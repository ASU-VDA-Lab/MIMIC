module fake_jpeg_8316_n_141 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_2),
.B(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

OR2x2_ASAP7_75t_SL g29 ( 
.A(n_0),
.B(n_4),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_15),
.B(n_1),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_15),
.B1(n_16),
.B2(n_27),
.Y(n_49)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_26),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_53),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_29),
.B(n_3),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_30),
.B(n_26),
.C(n_24),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_19),
.B1(n_24),
.B2(n_18),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_16),
.B1(n_27),
.B2(n_22),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_50),
.A2(n_37),
.B1(n_21),
.B2(n_22),
.Y(n_54)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_66),
.B1(n_71),
.B2(n_18),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_13),
.C(n_11),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_58),
.Y(n_72)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_57),
.Y(n_73)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_70),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_69),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_21),
.Y(n_65)
);

AO21x2_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_37),
.B(n_38),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_68),
.A2(n_52),
.B1(n_42),
.B2(n_38),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_36),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_33),
.B1(n_39),
.B2(n_19),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_39),
.C(n_46),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_75),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_46),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_79),
.B1(n_84),
.B2(n_68),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_33),
.B1(n_48),
.B2(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_68),
.B(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_85),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_38),
.B1(n_34),
.B2(n_25),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_2),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_34),
.C(n_14),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_64),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_89),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_66),
.B(n_59),
.Y(n_91)
);

FAx1_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_85),
.CI(n_72),
.CON(n_112),
.SN(n_112)
);

INVxp67_ASAP7_75t_SL g93 ( 
.A(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_100),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_98),
.B1(n_68),
.B2(n_57),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_87),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_64),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_99),
.Y(n_103)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_104),
.A2(n_110),
.B(n_63),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_75),
.C(n_74),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_88),
.C(n_96),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_76),
.B(n_68),
.C(n_77),
.D(n_82),
.Y(n_107)
);

MAJx2_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_94),
.C(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_76),
.Y(n_108)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_100),
.A2(n_86),
.B1(n_56),
.B2(n_63),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_90),
.B(n_98),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_118),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_106),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_119),
.C(n_109),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_105),
.B(n_14),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_107),
.B(n_103),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_110),
.B1(n_111),
.B2(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_123),
.Y(n_130)
);

OA21x2_ASAP7_75t_SL g129 ( 
.A1(n_124),
.A2(n_126),
.B(n_117),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_113),
.B1(n_116),
.B2(n_114),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_112),
.C(n_56),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_116),
.B1(n_115),
.B2(n_114),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_114),
.B1(n_126),
.B2(n_124),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_112),
.C(n_13),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_132),
.B(n_134),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_9),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_127),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_136),
.Y(n_139)
);

AOI322xp5_ASAP7_75t_L g136 ( 
.A1(n_133),
.A2(n_128),
.A3(n_25),
.B1(n_20),
.B2(n_6),
.C1(n_3),
.C2(n_5),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_25),
.B(n_20),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_139),
.Y(n_141)
);


endmodule