module fake_aes_2782_n_677 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_677);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_677;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g77 ( .A(n_73), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_14), .Y(n_78) );
INVxp67_ASAP7_75t_L g79 ( .A(n_50), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_9), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_23), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_6), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_17), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_32), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_62), .Y(n_85) );
BUFx3_ASAP7_75t_L g86 ( .A(n_58), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_8), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_20), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_59), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_70), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_1), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_57), .Y(n_92) );
OR2x2_ASAP7_75t_L g93 ( .A(n_29), .B(n_0), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_1), .Y(n_94) );
NOR2xp67_ASAP7_75t_L g95 ( .A(n_65), .B(n_30), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_72), .Y(n_96) );
INVxp33_ASAP7_75t_SL g97 ( .A(n_45), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_52), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_26), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_69), .Y(n_100) );
INVx2_ASAP7_75t_SL g101 ( .A(n_49), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_56), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_75), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_42), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_4), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_55), .Y(n_106) );
NOR2xp67_ASAP7_75t_L g107 ( .A(n_46), .B(n_6), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_34), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_40), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_12), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_10), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_66), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_18), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_8), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_44), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_31), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_9), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_67), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_47), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_0), .Y(n_120) );
CKINVDCx14_ASAP7_75t_R g121 ( .A(n_35), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_22), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_36), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_77), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_86), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_86), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_94), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_103), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_114), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_114), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_80), .B(n_2), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_82), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_108), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_101), .Y(n_134) );
NOR2xp33_ASAP7_75t_R g135 ( .A(n_121), .B(n_33), .Y(n_135) );
BUFx2_ASAP7_75t_L g136 ( .A(n_94), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_81), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_119), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_101), .B(n_2), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_80), .B(n_3), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_99), .B(n_3), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_87), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_87), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_90), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_119), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_78), .B(n_4), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_91), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_91), .Y(n_149) );
XOR2xp5_ASAP7_75t_L g150 ( .A(n_100), .B(n_5), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_84), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_84), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_85), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g154 ( .A1(n_93), .A2(n_5), .B1(n_7), .B2(n_10), .Y(n_154) );
OAI21x1_ASAP7_75t_L g155 ( .A1(n_85), .A2(n_39), .B(n_74), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_90), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_105), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_93), .Y(n_158) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_88), .A2(n_38), .B(n_71), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_111), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_88), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_89), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_89), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_112), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_102), .B(n_7), .Y(n_165) );
INVx4_ASAP7_75t_SL g166 ( .A(n_131), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_156), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_131), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_125), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_158), .B(n_92), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_158), .B(n_98), .Y(n_171) );
BUFx2_ASAP7_75t_L g172 ( .A(n_136), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_136), .B(n_92), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_134), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_125), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_128), .B(n_96), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_134), .B(n_96), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_145), .B(n_79), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_145), .B(n_97), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_131), .B(n_112), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_125), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_151), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_127), .Y(n_183) );
AO22x2_ASAP7_75t_L g184 ( .A1(n_154), .A2(n_115), .B1(n_113), .B2(n_118), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_141), .B(n_118), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_141), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_125), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_141), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_125), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_126), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_137), .A2(n_97), .B1(n_110), .B2(n_120), .Y(n_191) );
INVx4_ASAP7_75t_L g192 ( .A(n_126), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_126), .Y(n_193) );
AND2x6_ASAP7_75t_L g194 ( .A(n_137), .B(n_113), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_129), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_132), .B(n_98), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_130), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_124), .B(n_123), .Y(n_198) );
NOR2x1p5_ASAP7_75t_L g199 ( .A(n_124), .B(n_117), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_133), .B(n_122), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_151), .Y(n_201) );
INVx4_ASAP7_75t_L g202 ( .A(n_126), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_152), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_152), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_159), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_153), .Y(n_206) );
NAND3xp33_ASAP7_75t_SL g207 ( .A(n_156), .B(n_106), .C(n_109), .Y(n_207) );
AND2x2_ASAP7_75t_SL g208 ( .A(n_140), .B(n_115), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_143), .B(n_144), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_162), .B(n_104), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_159), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_138), .B(n_95), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_163), .B(n_116), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_148), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_138), .B(n_107), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_126), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_164), .B(n_110), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_139), .Y(n_218) );
OR2x2_ASAP7_75t_L g219 ( .A(n_133), .B(n_110), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_149), .B(n_110), .Y(n_220) );
AND2x6_ASAP7_75t_L g221 ( .A(n_164), .B(n_110), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_157), .B(n_83), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_166), .B(n_196), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_220), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_217), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_220), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_180), .B(n_161), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_170), .B(n_160), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_174), .Y(n_229) );
INVxp67_ASAP7_75t_L g230 ( .A(n_172), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_192), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_174), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_182), .Y(n_233) );
INVx2_ASAP7_75t_SL g234 ( .A(n_171), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_172), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_217), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_194), .Y(n_237) );
OR2x6_ASAP7_75t_L g238 ( .A(n_184), .B(n_147), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_217), .Y(n_239) );
INVx5_ASAP7_75t_L g240 ( .A(n_221), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_171), .B(n_165), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_209), .B(n_161), .Y(n_242) );
BUFx2_ASAP7_75t_L g243 ( .A(n_196), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_168), .A2(n_159), .B(n_155), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_166), .B(n_153), .Y(n_245) );
NAND2xp33_ASAP7_75t_SL g246 ( .A(n_199), .B(n_135), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_182), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_192), .Y(n_248) );
INVx2_ASAP7_75t_SL g249 ( .A(n_219), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_166), .B(n_142), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_183), .Y(n_251) );
NOR3xp33_ASAP7_75t_SL g252 ( .A(n_207), .B(n_150), .C(n_127), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_208), .A2(n_146), .B1(n_139), .B2(n_159), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_166), .B(n_155), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_203), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_208), .B(n_146), .Y(n_256) );
NOR2xp33_ASAP7_75t_SL g257 ( .A(n_194), .B(n_146), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_173), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_180), .B(n_146), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_194), .Y(n_260) );
NAND3xp33_ASAP7_75t_SL g261 ( .A(n_167), .B(n_183), .C(n_179), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_201), .Y(n_262) );
AND2x6_ASAP7_75t_L g263 ( .A(n_180), .B(n_139), .Y(n_263) );
INVxp67_ASAP7_75t_L g264 ( .A(n_176), .Y(n_264) );
INVx5_ASAP7_75t_L g265 ( .A(n_221), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_209), .B(n_146), .Y(n_266) );
OAI21xp33_ASAP7_75t_L g267 ( .A1(n_203), .A2(n_139), .B(n_150), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_185), .B(n_139), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_167), .Y(n_269) );
NAND2xp33_ASAP7_75t_L g270 ( .A(n_194), .B(n_37), .Y(n_270) );
CKINVDCx8_ASAP7_75t_R g271 ( .A(n_185), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_184), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_201), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_184), .A2(n_11), .B1(n_13), .B2(n_14), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_204), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_185), .B(n_15), .Y(n_276) );
NAND2xp33_ASAP7_75t_L g277 ( .A(n_194), .B(n_48), .Y(n_277) );
BUFx8_ASAP7_75t_L g278 ( .A(n_219), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_214), .B(n_43), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_213), .B(n_15), .Y(n_280) );
AND2x4_ASAP7_75t_SL g281 ( .A(n_186), .B(n_188), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_215), .B(n_222), .Y(n_282) );
INVxp67_ASAP7_75t_L g283 ( .A(n_177), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_178), .B(n_51), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_238), .A2(n_194), .B1(n_184), .B2(n_215), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_235), .B(n_230), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_242), .Y(n_287) );
BUFx2_ASAP7_75t_L g288 ( .A(n_278), .Y(n_288) );
INVx2_ASAP7_75t_SL g289 ( .A(n_278), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_225), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_269), .B(n_200), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_225), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_227), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_228), .B(n_191), .Y(n_294) );
OAI22xp33_ASAP7_75t_L g295 ( .A1(n_238), .A2(n_210), .B1(n_198), .B2(n_195), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_241), .B(n_197), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_249), .B(n_206), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_227), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_238), .A2(n_274), .B1(n_276), .B2(n_271), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_274), .A2(n_204), .B1(n_206), .B2(n_201), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_244), .A2(n_205), .B(n_211), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_237), .B(n_215), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_264), .B(n_211), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_236), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_224), .Y(n_305) );
OR2x6_ASAP7_75t_L g306 ( .A(n_223), .B(n_212), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_258), .B(n_205), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g308 ( .A1(n_234), .A2(n_205), .B1(n_211), .B2(n_192), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_236), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_266), .Y(n_310) );
OR2x6_ASAP7_75t_L g311 ( .A(n_223), .B(n_205), .Y(n_311) );
A2O1A1Ixp33_ASAP7_75t_L g312 ( .A1(n_233), .A2(n_205), .B(n_211), .C(n_216), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_226), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_243), .A2(n_211), .B1(n_202), .B2(n_221), .Y(n_314) );
INVx8_ASAP7_75t_L g315 ( .A(n_263), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_237), .B(n_202), .Y(n_316) );
AOI22xp33_ASAP7_75t_SL g317 ( .A1(n_272), .A2(n_221), .B1(n_202), .B2(n_16), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_282), .B(n_221), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_282), .B(n_221), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_283), .B(n_16), .Y(n_320) );
BUFx12f_ASAP7_75t_L g321 ( .A(n_251), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_247), .A2(n_218), .B1(n_216), .B2(n_193), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_239), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_237), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_261), .B(n_187), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_239), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_268), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_260), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_268), .Y(n_329) );
INVx4_ASAP7_75t_L g330 ( .A(n_260), .Y(n_330) );
BUFx3_ASAP7_75t_L g331 ( .A(n_262), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_246), .Y(n_332) );
NOR2x1_ASAP7_75t_L g333 ( .A(n_280), .B(n_218), .Y(n_333) );
NAND2x1p5_ASAP7_75t_L g334 ( .A(n_324), .B(n_260), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_324), .Y(n_335) );
INVx6_ASAP7_75t_L g336 ( .A(n_330), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_286), .Y(n_337) );
OA21x2_ASAP7_75t_L g338 ( .A1(n_312), .A2(n_253), .B(n_254), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_301), .A2(n_254), .B(n_256), .Y(n_339) );
OAI21x1_ASAP7_75t_L g340 ( .A1(n_333), .A2(n_279), .B(n_284), .Y(n_340) );
AO21x2_ASAP7_75t_L g341 ( .A1(n_295), .A2(n_279), .B(n_270), .Y(n_341) );
OAI21x1_ASAP7_75t_L g342 ( .A1(n_308), .A2(n_250), .B(n_255), .Y(n_342) );
INVx1_ASAP7_75t_SL g343 ( .A(n_297), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_299), .A2(n_267), .B1(n_272), .B2(n_281), .Y(n_344) );
OA21x2_ASAP7_75t_L g345 ( .A1(n_299), .A2(n_187), .B(n_175), .Y(n_345) );
OAI21x1_ASAP7_75t_L g346 ( .A1(n_322), .A2(n_275), .B(n_259), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_287), .Y(n_347) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_324), .B(n_245), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_297), .Y(n_349) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_300), .A2(n_181), .B(n_175), .Y(n_350) );
INVx2_ASAP7_75t_SL g351 ( .A(n_315), .Y(n_351) );
OAI21x1_ASAP7_75t_L g352 ( .A1(n_322), .A2(n_181), .B(n_189), .Y(n_352) );
OAI21xp5_ASAP7_75t_L g353 ( .A1(n_303), .A2(n_277), .B(n_229), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_293), .B(n_267), .Y(n_354) );
AO21x2_ASAP7_75t_L g355 ( .A1(n_300), .A2(n_169), .B(n_189), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_288), .Y(n_356) );
OAI21x1_ASAP7_75t_L g357 ( .A1(n_303), .A2(n_169), .B(n_190), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_328), .Y(n_358) );
NOR2xp67_ASAP7_75t_L g359 ( .A(n_330), .B(n_245), .Y(n_359) );
OAI21xp5_ASAP7_75t_L g360 ( .A1(n_307), .A2(n_232), .B(n_257), .Y(n_360) );
BUFx2_ASAP7_75t_L g361 ( .A(n_311), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_328), .Y(n_362) );
OAI221xp5_ASAP7_75t_L g363 ( .A1(n_285), .A2(n_252), .B1(n_273), .B2(n_257), .C(n_248), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_325), .A2(n_193), .B(n_190), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_344), .A2(n_291), .B1(n_289), .B2(n_320), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_363), .A2(n_321), .B1(n_317), .B2(n_298), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_363), .A2(n_294), .B1(n_313), .B2(n_305), .Y(n_367) );
AOI222xp33_ASAP7_75t_L g368 ( .A1(n_347), .A2(n_296), .B1(n_294), .B2(n_332), .C1(n_327), .C2(n_329), .Y(n_368) );
AOI222xp33_ASAP7_75t_L g369 ( .A1(n_347), .A2(n_307), .B1(n_326), .B2(n_323), .C1(n_302), .C2(n_310), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_341), .A2(n_311), .B(n_319), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_343), .A2(n_311), .B1(n_315), .B2(n_319), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_337), .A2(n_306), .B1(n_263), .B2(n_273), .Y(n_372) );
OAI211xp5_ASAP7_75t_L g373 ( .A1(n_356), .A2(n_318), .B(n_331), .C(n_314), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_343), .B(n_304), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_337), .A2(n_292), .B1(n_290), .B2(n_309), .C(n_318), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_336), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_349), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_357), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g379 ( .A1(n_349), .A2(n_306), .B1(n_231), .B2(n_316), .C(n_328), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_354), .A2(n_306), .B1(n_263), .B2(n_315), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_346), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_346), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_341), .A2(n_265), .B(n_240), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_341), .A2(n_265), .B(n_240), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_354), .A2(n_263), .B1(n_265), .B2(n_240), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_351), .B(n_19), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_361), .A2(n_21), .B1(n_24), .B2(n_25), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_350), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_361), .A2(n_27), .B1(n_28), .B2(n_41), .Y(n_389) );
OAI21xp5_ASAP7_75t_L g390 ( .A1(n_339), .A2(n_353), .B(n_342), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g391 ( .A1(n_353), .A2(n_53), .B1(n_54), .B2(n_60), .C(n_61), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_378), .Y(n_392) );
INVx4_ASAP7_75t_R g393 ( .A(n_376), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_377), .B(n_355), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_386), .B(n_335), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_386), .B(n_335), .Y(n_396) );
NAND2x1p5_ASAP7_75t_L g397 ( .A(n_386), .B(n_362), .Y(n_397) );
INVxp67_ASAP7_75t_SL g398 ( .A(n_377), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_381), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_381), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_378), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_374), .B(n_355), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_365), .B(n_351), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_382), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_374), .B(n_355), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_376), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_382), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_368), .B(n_355), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_388), .Y(n_409) );
INVxp67_ASAP7_75t_SL g410 ( .A(n_369), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_367), .B(n_345), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_388), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_366), .B(n_345), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_390), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_370), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_379), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_371), .B(n_345), .Y(n_417) );
OR2x6_ASAP7_75t_L g418 ( .A(n_383), .B(n_350), .Y(n_418) );
INVx2_ASAP7_75t_SL g419 ( .A(n_387), .Y(n_419) );
BUFx12f_ASAP7_75t_L g420 ( .A(n_373), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_391), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_375), .Y(n_422) );
OR2x6_ASAP7_75t_L g423 ( .A(n_384), .B(n_350), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_380), .B(n_345), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_372), .Y(n_425) );
OAI31xp33_ASAP7_75t_L g426 ( .A1(n_408), .A2(n_389), .A3(n_385), .B(n_348), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_392), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_392), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_409), .B(n_364), .Y(n_429) );
INVx3_ASAP7_75t_L g430 ( .A(n_392), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_409), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_401), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_412), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_408), .B(n_341), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_412), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_402), .B(n_338), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_406), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_399), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_402), .B(n_338), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_405), .B(n_338), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_405), .B(n_338), .Y(n_441) );
BUFx2_ASAP7_75t_L g442 ( .A(n_397), .Y(n_442) );
NOR3xp33_ASAP7_75t_L g443 ( .A(n_410), .B(n_359), .C(n_339), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_394), .B(n_364), .Y(n_444) );
BUFx2_ASAP7_75t_L g445 ( .A(n_397), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_399), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_400), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_400), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_401), .Y(n_449) );
AOI211xp5_ASAP7_75t_SL g450 ( .A1(n_422), .A2(n_359), .B(n_358), .C(n_335), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_394), .B(n_364), .Y(n_451) );
BUFx2_ASAP7_75t_L g452 ( .A(n_397), .Y(n_452) );
OAI221xp5_ASAP7_75t_L g453 ( .A1(n_403), .A2(n_360), .B1(n_336), .B2(n_348), .C(n_334), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_407), .Y(n_454) );
BUFx3_ASAP7_75t_L g455 ( .A(n_395), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_401), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_407), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_425), .A2(n_336), .B1(n_360), .B2(n_342), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_413), .B(n_414), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_404), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_413), .B(n_358), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_414), .B(n_358), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_404), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_404), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_398), .B(n_357), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_420), .Y(n_466) );
AOI221xp5_ASAP7_75t_L g467 ( .A1(n_416), .A2(n_348), .B1(n_362), .B2(n_334), .C(n_336), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_416), .B(n_352), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_415), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_415), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_419), .A2(n_362), .B1(n_334), .B2(n_336), .C(n_340), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_424), .B(n_352), .Y(n_472) );
INVxp67_ASAP7_75t_L g473 ( .A(n_424), .Y(n_473) );
NAND2x1_ASAP7_75t_L g474 ( .A(n_460), .B(n_393), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_455), .B(n_423), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_437), .B(n_419), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_431), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_466), .A2(n_420), .B1(n_421), .B2(n_396), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_431), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_433), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_459), .B(n_395), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_459), .B(n_417), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_436), .B(n_417), .Y(n_483) );
NOR2x1_ASAP7_75t_L g484 ( .A(n_442), .B(n_395), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_436), .B(n_423), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_440), .B(n_423), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_440), .B(n_423), .Y(n_487) );
INVxp67_ASAP7_75t_L g488 ( .A(n_442), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_433), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_455), .B(n_423), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_441), .B(n_418), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_435), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_439), .B(n_411), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_435), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_438), .Y(n_495) );
OAI222xp33_ASAP7_75t_L g496 ( .A1(n_453), .A2(n_418), .B1(n_421), .B2(n_396), .C1(n_395), .C2(n_393), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_441), .B(n_418), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_473), .B(n_418), .Y(n_498) );
INVx1_ASAP7_75t_SL g499 ( .A(n_445), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_473), .B(n_396), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_439), .B(n_418), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_438), .B(n_396), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_445), .Y(n_503) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_452), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_446), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_446), .B(n_340), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_447), .Y(n_507) );
NAND3xp33_ASAP7_75t_L g508 ( .A(n_443), .B(n_340), .C(n_64), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_463), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_444), .B(n_63), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_447), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_426), .A2(n_68), .B1(n_76), .B2(n_443), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_463), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_444), .B(n_451), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_451), .B(n_461), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_461), .B(n_472), .Y(n_516) );
INVx3_ASAP7_75t_L g517 ( .A(n_430), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_448), .B(n_457), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_455), .B(n_469), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_448), .Y(n_520) );
NAND2x1p5_ASAP7_75t_L g521 ( .A(n_452), .B(n_465), .Y(n_521) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_450), .A2(n_426), .B(n_467), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_472), .B(n_457), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_471), .B(n_467), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_469), .B(n_454), .Y(n_525) );
BUFx2_ASAP7_75t_SL g526 ( .A(n_463), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_454), .B(n_464), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_430), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_460), .B(n_464), .Y(n_529) );
INVx2_ASAP7_75t_SL g530 ( .A(n_430), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_514), .B(n_470), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_514), .B(n_470), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_515), .B(n_516), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_525), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_525), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_515), .B(n_429), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_516), .B(n_429), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_499), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_525), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_523), .B(n_434), .Y(n_540) );
OAI21xp33_ASAP7_75t_L g541 ( .A1(n_522), .A2(n_434), .B(n_450), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_523), .B(n_462), .Y(n_542) );
NOR3xp33_ASAP7_75t_SL g543 ( .A(n_524), .B(n_453), .C(n_471), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_503), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_477), .Y(n_545) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_524), .A2(n_468), .B(n_465), .Y(n_546) );
NAND2x1p5_ASAP7_75t_L g547 ( .A(n_474), .B(n_429), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_483), .B(n_429), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_483), .B(n_456), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_476), .B(n_462), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_482), .B(n_456), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g552 ( .A(n_512), .B(n_458), .C(n_468), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_479), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_482), .B(n_430), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_480), .Y(n_555) );
INVxp67_ASAP7_75t_SL g556 ( .A(n_521), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_485), .B(n_456), .Y(n_557) );
INVxp67_ASAP7_75t_SL g558 ( .A(n_521), .Y(n_558) );
A2O1A1O1Ixp25_ASAP7_75t_L g559 ( .A1(n_489), .A2(n_456), .B(n_428), .C(n_432), .D(n_449), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_485), .B(n_427), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_529), .Y(n_561) );
INVx2_ASAP7_75t_SL g562 ( .A(n_504), .Y(n_562) );
NOR2xp67_ASAP7_75t_SL g563 ( .A(n_526), .B(n_427), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_493), .B(n_427), .Y(n_564) );
NOR2xp67_ASAP7_75t_SL g565 ( .A(n_510), .B(n_428), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_492), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_486), .B(n_428), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_478), .B(n_432), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_486), .B(n_432), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_493), .B(n_449), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_475), .B(n_449), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_487), .B(n_491), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_487), .B(n_491), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_494), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_497), .B(n_498), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_497), .B(n_498), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_527), .B(n_511), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_495), .Y(n_578) );
NOR2x1_ASAP7_75t_L g579 ( .A(n_474), .B(n_496), .Y(n_579) );
NAND2x1_ASAP7_75t_L g580 ( .A(n_475), .B(n_490), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_501), .B(n_527), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_508), .A2(n_484), .B(n_506), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_533), .B(n_531), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_533), .B(n_531), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_532), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_561), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_577), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_532), .Y(n_588) );
OAI21xp5_ASAP7_75t_SL g589 ( .A1(n_579), .A2(n_488), .B(n_510), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_540), .B(n_529), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_581), .B(n_507), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_545), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g593 ( .A1(n_559), .A2(n_501), .B1(n_504), .B2(n_481), .Y(n_593) );
NOR3xp33_ASAP7_75t_L g594 ( .A(n_541), .B(n_518), .C(n_500), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_545), .Y(n_595) );
NOR2xp33_ASAP7_75t_SL g596 ( .A(n_563), .B(n_504), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_543), .B(n_504), .Y(n_597) );
INVxp67_ASAP7_75t_SL g598 ( .A(n_563), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_555), .Y(n_599) );
OAI22xp33_ASAP7_75t_L g600 ( .A1(n_580), .A2(n_528), .B1(n_530), .B2(n_517), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_538), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_547), .B(n_530), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_555), .Y(n_603) );
INVxp67_ASAP7_75t_SL g604 ( .A(n_565), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_568), .A2(n_519), .B1(n_490), .B2(n_475), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_572), .B(n_490), .Y(n_606) );
OAI22xp5_ASAP7_75t_SL g607 ( .A1(n_580), .A2(n_519), .B1(n_528), .B2(n_520), .Y(n_607) );
O2A1O1Ixp33_ASAP7_75t_L g608 ( .A1(n_544), .A2(n_505), .B(n_502), .C(n_517), .Y(n_608) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_552), .A2(n_519), .B(n_517), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_581), .B(n_509), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_553), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_564), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_550), .A2(n_509), .B1(n_513), .B2(n_534), .Y(n_613) );
AOI21xp33_ASAP7_75t_SL g614 ( .A1(n_547), .A2(n_513), .B(n_546), .Y(n_614) );
AOI21xp33_ASAP7_75t_L g615 ( .A1(n_556), .A2(n_558), .B(n_562), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_535), .A2(n_549), .B1(n_539), .B2(n_551), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_542), .B(n_574), .Y(n_617) );
AOI221xp5_ASAP7_75t_L g618 ( .A1(n_566), .A2(n_578), .B1(n_554), .B2(n_551), .C(n_539), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_549), .A2(n_565), .B1(n_548), .B2(n_569), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_586), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_592), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_595), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_589), .A2(n_547), .B(n_582), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_599), .Y(n_624) );
XOR2xp5_ASAP7_75t_L g625 ( .A(n_605), .B(n_564), .Y(n_625) );
XOR2x2_ASAP7_75t_L g626 ( .A(n_601), .B(n_573), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_603), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_610), .B(n_570), .Y(n_628) );
INVxp67_ASAP7_75t_L g629 ( .A(n_597), .Y(n_629) );
INVxp67_ASAP7_75t_L g630 ( .A(n_597), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_611), .Y(n_631) );
AOI21xp33_ASAP7_75t_SL g632 ( .A1(n_593), .A2(n_570), .B(n_562), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_612), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_591), .Y(n_634) );
OAI211xp5_ASAP7_75t_SL g635 ( .A1(n_593), .A2(n_573), .B(n_572), .C(n_575), .Y(n_635) );
OA22x2_ASAP7_75t_L g636 ( .A1(n_607), .A2(n_536), .B1(n_537), .B2(n_576), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_612), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_594), .B(n_548), .Y(n_638) );
AOI21xp33_ASAP7_75t_L g639 ( .A1(n_598), .A2(n_571), .B(n_557), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_585), .Y(n_640) );
XNOR2x1_ASAP7_75t_L g641 ( .A(n_587), .B(n_576), .Y(n_641) );
INVxp67_ASAP7_75t_SL g642 ( .A(n_608), .Y(n_642) );
AOI31xp33_ASAP7_75t_L g643 ( .A1(n_629), .A2(n_614), .A3(n_609), .B(n_615), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_623), .A2(n_602), .B(n_600), .Y(n_644) );
O2A1O1Ixp33_ASAP7_75t_L g645 ( .A1(n_642), .A2(n_604), .B(n_602), .C(n_600), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_621), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g647 ( .A1(n_629), .A2(n_619), .B(n_618), .Y(n_647) );
NOR2x1_ASAP7_75t_L g648 ( .A(n_635), .B(n_641), .Y(n_648) );
OAI22xp33_ASAP7_75t_L g649 ( .A1(n_636), .A2(n_596), .B1(n_584), .B2(n_583), .Y(n_649) );
OAI21xp33_ASAP7_75t_L g650 ( .A1(n_635), .A2(n_616), .B(n_619), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_636), .A2(n_616), .B1(n_613), .B2(n_617), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_622), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_624), .Y(n_653) );
AOI31xp33_ASAP7_75t_L g654 ( .A1(n_630), .A2(n_606), .A3(n_588), .B(n_536), .Y(n_654) );
NAND2x1_ASAP7_75t_SL g655 ( .A(n_620), .B(n_537), .Y(n_655) );
NAND3xp33_ASAP7_75t_SL g656 ( .A(n_644), .B(n_632), .C(n_630), .Y(n_656) );
A2O1A1Ixp33_ASAP7_75t_L g657 ( .A1(n_648), .A2(n_642), .B(n_638), .C(n_639), .Y(n_657) );
NAND2x1p5_ASAP7_75t_L g658 ( .A(n_644), .B(n_628), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_649), .A2(n_625), .B1(n_634), .B2(n_631), .C(n_633), .Y(n_659) );
AOI221x1_ASAP7_75t_L g660 ( .A1(n_650), .A2(n_627), .B1(n_637), .B2(n_633), .C(n_626), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_645), .A2(n_627), .B(n_637), .Y(n_661) );
OAI211xp5_ASAP7_75t_L g662 ( .A1(n_647), .A2(n_590), .B(n_640), .C(n_575), .Y(n_662) );
NOR3x1_ASAP7_75t_L g663 ( .A(n_643), .B(n_571), .C(n_557), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_657), .B(n_651), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_658), .B(n_654), .Y(n_665) );
NOR2x1_ASAP7_75t_L g666 ( .A(n_656), .B(n_646), .Y(n_666) );
AOI211xp5_ASAP7_75t_SL g667 ( .A1(n_659), .A2(n_652), .B(n_653), .C(n_655), .Y(n_667) );
NAND2x1p5_ASAP7_75t_L g668 ( .A(n_666), .B(n_663), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_665), .Y(n_669) );
AND3x4_ASAP7_75t_L g670 ( .A(n_667), .B(n_660), .C(n_662), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_669), .Y(n_671) );
OR3x1_ASAP7_75t_L g672 ( .A(n_670), .B(n_664), .C(n_661), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_671), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_673), .B(n_672), .Y(n_674) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_674), .Y(n_675) );
AOI222xp33_ASAP7_75t_L g676 ( .A1(n_675), .A2(n_668), .B1(n_571), .B2(n_569), .C1(n_567), .C2(n_560), .Y(n_676) );
AOI21xp33_ASAP7_75t_SL g677 ( .A1(n_676), .A2(n_560), .B(n_567), .Y(n_677) );
endmodule