module fake_netlist_5_2340_n_4387 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_451, n_408, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_452, n_397, n_111, n_155, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_470, n_325, n_449, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_457, n_297, n_156, n_5, n_225, n_377, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_430, n_313, n_88, n_479, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_213, n_129, n_342, n_482, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_309, n_30, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_85, n_463, n_239, n_466, n_420, n_55, n_49, n_310, n_54, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_441, n_450, n_312, n_476, n_429, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_480, n_237, n_425, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_409, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_391, n_434, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_52, n_278, n_110, n_4387);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_451;
input n_408;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_213;
input n_129;
input n_342;
input n_482;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_85;
input n_463;
input n_239;
input n_466;
input n_420;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_480;
input n_237;
input n_425;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_409;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_391;
input n_434;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_4387;

wire n_924;
wire n_1263;
wire n_3304;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_2756;
wire n_3912;
wire n_1423;
wire n_1126;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_3241;
wire n_785;
wire n_4129;
wire n_549;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_532;
wire n_1161;
wire n_3795;
wire n_3863;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_1780;
wire n_3256;
wire n_3732;
wire n_1488;
wire n_4250;
wire n_667;
wire n_2955;
wire n_2899;
wire n_790;
wire n_3619;
wire n_1055;
wire n_3541;
wire n_3622;
wire n_4112;
wire n_2386;
wire n_3596;
wire n_1501;
wire n_4337;
wire n_2395;
wire n_3906;
wire n_4138;
wire n_880;
wire n_4127;
wire n_3086;
wire n_3297;
wire n_544;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_552;
wire n_1528;
wire n_4217;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2821;
wire n_2520;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_4292;
wire n_2568;
wire n_3641;
wire n_956;
wire n_564;
wire n_4240;
wire n_1738;
wire n_2021;
wire n_3728;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_4236;
wire n_3088;
wire n_4202;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_551;
wire n_2143;
wire n_3713;
wire n_2853;
wire n_3615;
wire n_2059;
wire n_1323;
wire n_3663;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_3766;
wire n_1353;
wire n_800;
wire n_3595;
wire n_3246;
wire n_3202;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_3813;
wire n_1789;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_671;
wire n_4238;
wire n_819;
wire n_1451;
wire n_1022;
wire n_4038;
wire n_2302;
wire n_915;
wire n_4109;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_3341;
wire n_1947;
wire n_1264;
wire n_3587;
wire n_2114;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_1494;
wire n_3407;
wire n_3599;
wire n_3571;
wire n_3785;
wire n_625;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_854;
wire n_3621;
wire n_4211;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_3434;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1152;
wire n_3501;
wire n_3448;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_3019;
wire n_3039;
wire n_4013;
wire n_2011;
wire n_2096;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_877;
wire n_2105;
wire n_2538;
wire n_3776;
wire n_2024;
wire n_2530;
wire n_4242;
wire n_1696;
wire n_2483;
wire n_3163;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_3710;
wire n_4243;
wire n_3851;
wire n_1860;
wire n_2543;
wire n_4155;
wire n_1359;
wire n_530;
wire n_1728;
wire n_1107;
wire n_2031;
wire n_556;
wire n_2076;
wire n_3036;
wire n_2482;
wire n_3695;
wire n_3891;
wire n_4145;
wire n_2677;
wire n_1230;
wire n_4144;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_3010;
wire n_3180;
wire n_3379;
wire n_3832;
wire n_4374;
wire n_3532;
wire n_2770;
wire n_1124;
wire n_3987;
wire n_4061;
wire n_4131;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_902;
wire n_1705;
wire n_1294;
wire n_659;
wire n_1104;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_3531;
wire n_3403;
wire n_4021;
wire n_579;
wire n_1698;
wire n_3880;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2963;
wire n_3624;
wire n_3834;
wire n_2142;
wire n_3186;
wire n_3461;
wire n_3082;
wire n_1154;
wire n_2189;
wire n_3796;
wire n_3332;
wire n_1242;
wire n_3283;
wire n_1135;
wire n_3048;
wire n_3258;
wire n_3937;
wire n_3696;
wire n_519;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1243;
wire n_1016;
wire n_4315;
wire n_546;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_1280;
wire n_3277;
wire n_3782;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_2478;
wire n_3650;
wire n_3786;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_3638;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_2537;
wire n_2983;
wire n_3763;
wire n_569;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_920;
wire n_2515;
wire n_3022;
wire n_3810;
wire n_2466;
wire n_1517;
wire n_2091;
wire n_2652;
wire n_2635;
wire n_4311;
wire n_1289;
wire n_4264;
wire n_3631;
wire n_2715;
wire n_3806;
wire n_3087;
wire n_4197;
wire n_2085;
wire n_3489;
wire n_1669;
wire n_2566;
wire n_1949;
wire n_976;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_3060;
wire n_4276;
wire n_2651;
wire n_3947;
wire n_4358;
wire n_3490;
wire n_3656;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_3437;
wire n_3868;
wire n_4369;
wire n_2099;
wire n_2408;
wire n_4168;
wire n_3446;
wire n_3353;
wire n_1877;
wire n_4203;
wire n_3687;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_1723;
wire n_955;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_4350;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_3156;
wire n_550;
wire n_696;
wire n_3101;
wire n_3669;
wire n_897;
wire n_798;
wire n_3376;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_3653;
wire n_1414;
wire n_1216;
wire n_580;
wire n_2693;
wire n_3798;
wire n_3702;
wire n_1040;
wire n_4065;
wire n_3836;
wire n_2202;
wire n_2648;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1852;
wire n_2159;
wire n_578;
wire n_2976;
wire n_3876;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_4135;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_4187;
wire n_1547;
wire n_1070;
wire n_777;
wire n_4166;
wire n_2089;
wire n_3420;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1071;
wire n_485;
wire n_1561;
wire n_1267;
wire n_1165;
wire n_496;
wire n_1801;
wire n_3985;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_3361;
wire n_1600;
wire n_521;
wire n_3744;
wire n_663;
wire n_845;
wire n_2235;
wire n_4263;
wire n_1862;
wire n_673;
wire n_837;
wire n_3980;
wire n_1239;
wire n_2915;
wire n_528;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_3291;
wire n_4255;
wire n_680;
wire n_1587;
wire n_1473;
wire n_2682;
wire n_3755;
wire n_553;
wire n_901;
wire n_2432;
wire n_3668;
wire n_813;
wire n_4258;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_3440;
wire n_3405;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_3563;
wire n_2934;
wire n_1672;
wire n_4237;
wire n_2699;
wire n_675;
wire n_2506;
wire n_4064;
wire n_888;
wire n_1880;
wire n_2769;
wire n_3550;
wire n_2337;
wire n_3542;
wire n_1167;
wire n_1626;
wire n_3436;
wire n_637;
wire n_2615;
wire n_3940;
wire n_1384;
wire n_1556;
wire n_3907;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_3841;
wire n_2238;
wire n_2118;
wire n_923;
wire n_2985;
wire n_691;
wire n_1151;
wire n_2944;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_3418;
wire n_2932;
wire n_2753;
wire n_2980;
wire n_1582;
wire n_3637;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_3262;
wire n_3136;
wire n_1836;
wire n_2868;
wire n_3395;
wire n_1450;
wire n_4080;
wire n_4006;
wire n_3141;
wire n_4226;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_3570;
wire n_3690;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_3986;
wire n_4376;
wire n_3716;
wire n_4025;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_3191;
wire n_571;
wire n_1585;
wire n_2712;
wire n_2684;
wire n_3837;
wire n_3593;
wire n_3193;
wire n_3885;
wire n_3936;
wire n_1971;
wire n_1599;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3507;
wire n_3273;
wire n_3821;
wire n_2713;
wire n_3544;
wire n_2700;
wire n_2644;
wire n_4310;
wire n_1211;
wire n_1197;
wire n_3367;
wire n_4020;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_3709;
wire n_1447;
wire n_907;
wire n_2251;
wire n_3096;
wire n_1377;
wire n_3915;
wire n_2370;
wire n_3496;
wire n_3954;
wire n_4114;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_3339;
wire n_2055;
wire n_3427;
wire n_3025;
wire n_3349;
wire n_1403;
wire n_3735;
wire n_4067;
wire n_2248;
wire n_4042;
wire n_4176;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_4385;
wire n_3320;
wire n_3007;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_3899;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_4159;
wire n_3714;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_3071;
wire n_3739;
wire n_4089;
wire n_3651;
wire n_3310;
wire n_3487;
wire n_593;
wire n_4333;
wire n_2258;
wire n_4069;
wire n_748;
wire n_1058;
wire n_1667;
wire n_586;
wire n_3359;
wire n_838;
wire n_2784;
wire n_3718;
wire n_3983;
wire n_2919;
wire n_3092;
wire n_1053;
wire n_3470;
wire n_1224;
wire n_2865;
wire n_4327;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_4195;
wire n_953;
wire n_1014;
wire n_4218;
wire n_1241;
wire n_3676;
wire n_2150;
wire n_3146;
wire n_4375;
wire n_2241;
wire n_2757;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_3781;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_3580;
wire n_4246;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_4353;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_534;
wire n_3106;
wire n_1882;
wire n_4164;
wire n_884;
wire n_3328;
wire n_944;
wire n_4130;
wire n_4234;
wire n_1754;
wire n_3889;
wire n_3611;
wire n_1623;
wire n_2862;
wire n_4256;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2674;
wire n_2606;
wire n_3187;
wire n_1565;
wire n_4088;
wire n_4224;
wire n_3508;
wire n_2828;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_4161;
wire n_647;
wire n_3433;
wire n_4024;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_3392;
wire n_3430;
wire n_3975;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_1319;
wire n_561;
wire n_2379;
wire n_3331;
wire n_3447;
wire n_2616;
wire n_2911;
wire n_3992;
wire n_3305;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_4148;
wire n_4151;
wire n_1883;
wire n_1906;
wire n_4103;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_3528;
wire n_3649;
wire n_2262;
wire n_4302;
wire n_2462;
wire n_2514;
wire n_4373;
wire n_1532;
wire n_4252;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_3625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_4331;
wire n_4160;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2293;
wire n_686;
wire n_3989;
wire n_2837;
wire n_847;
wire n_3804;
wire n_4051;
wire n_4344;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_3481;
wire n_2762;
wire n_4097;
wire n_558;
wire n_3655;
wire n_2808;
wire n_1276;
wire n_702;
wire n_3009;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_3981;
wire n_2108;
wire n_3640;
wire n_728;
wire n_1162;
wire n_1538;
wire n_2930;
wire n_4206;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3514;
wire n_3116;
wire n_1884;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_3602;
wire n_1038;
wire n_2967;
wire n_1369;
wire n_520;
wire n_3909;
wire n_2611;
wire n_4261;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_3207;
wire n_2581;
wire n_3944;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_3752;
wire n_4090;
wire n_809;
wire n_3923;
wire n_931;
wire n_1711;
wire n_599;
wire n_1891;
wire n_1662;
wire n_870;
wire n_1481;
wire n_2626;
wire n_3441;
wire n_3042;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_4001;
wire n_3047;
wire n_2510;
wire n_3526;
wire n_4219;
wire n_868;
wire n_2454;
wire n_4371;
wire n_639;
wire n_2804;
wire n_914;
wire n_3659;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_3120;
wire n_965;
wire n_1876;
wire n_1743;
wire n_4007;
wire n_3790;
wire n_4011;
wire n_4268;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2825;
wire n_2813;
wire n_2009;
wire n_1888;
wire n_759;
wire n_3643;
wire n_3895;
wire n_4194;
wire n_2222;
wire n_1892;
wire n_4120;
wire n_3510;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_4278;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_4142;
wire n_1189;
wire n_2690;
wire n_4082;
wire n_4028;
wire n_3370;
wire n_2215;
wire n_3479;
wire n_4085;
wire n_1259;
wire n_4073;
wire n_1690;
wire n_4260;
wire n_3819;
wire n_706;
wire n_746;
wire n_1649;
wire n_3150;
wire n_4163;
wire n_747;
wire n_2064;
wire n_784;
wire n_3978;
wire n_4325;
wire n_2449;
wire n_3867;
wire n_1733;
wire n_4372;
wire n_1244;
wire n_3500;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_3660;
wire n_2297;
wire n_4186;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_615;
wire n_851;
wire n_1759;
wire n_1788;
wire n_2177;
wire n_843;
wire n_2491;
wire n_3747;
wire n_523;
wire n_1537;
wire n_913;
wire n_705;
wire n_3833;
wire n_865;
wire n_2227;
wire n_3775;
wire n_4133;
wire n_678;
wire n_2671;
wire n_697;
wire n_4262;
wire n_4184;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_1798;
wire n_2022;
wire n_776;
wire n_3814;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_4099;
wire n_2592;
wire n_3416;
wire n_4379;
wire n_525;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_4340;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_3513;
wire n_4295;
wire n_649;
wire n_547;
wire n_2563;
wire n_1444;
wire n_4030;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_4334;
wire n_1674;
wire n_3725;
wire n_1833;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_3128;
wire n_1734;
wire n_3038;
wire n_744;
wire n_629;
wire n_590;
wire n_3770;
wire n_4014;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_3144;
wire n_4244;
wire n_2943;
wire n_2913;
wire n_4254;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_1233;
wire n_4179;
wire n_3469;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_1615;
wire n_4175;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_3317;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_3355;
wire n_604;
wire n_2007;
wire n_3220;
wire n_949;
wire n_2539;
wire n_3917;
wire n_3942;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_3855;
wire n_946;
wire n_1539;
wire n_2736;
wire n_4157;
wire n_4283;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_3765;
wire n_498;
wire n_1468;
wire n_1559;
wire n_3823;
wire n_1765;
wire n_3455;
wire n_1866;
wire n_4173;
wire n_689;
wire n_3158;
wire n_738;
wire n_1624;
wire n_3000;
wire n_640;
wire n_3452;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_3816;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_3113;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_2577;
wire n_3760;
wire n_4108;
wire n_4078;
wire n_1760;
wire n_2875;
wire n_936;
wire n_1500;
wire n_568;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_757;
wire n_3844;
wire n_3280;
wire n_2342;
wire n_633;
wire n_2856;
wire n_4054;
wire n_3471;
wire n_1832;
wire n_4156;
wire n_1851;
wire n_758;
wire n_999;
wire n_3205;
wire n_2046;
wire n_4146;
wire n_2848;
wire n_2741;
wire n_4360;
wire n_2937;
wire n_3666;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_3828;
wire n_2290;
wire n_1656;
wire n_3564;
wire n_3288;
wire n_1158;
wire n_3095;
wire n_3866;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_3988;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_3667;
wire n_1145;
wire n_878;
wire n_524;
wire n_3843;
wire n_3457;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_3856;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_3703;
wire n_4324;
wire n_1068;
wire n_3030;
wire n_3558;
wire n_1871;
wire n_2580;
wire n_3630;
wire n_2545;
wire n_2787;
wire n_3685;
wire n_4249;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_906;
wire n_3271;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_4086;
wire n_2412;
wire n_4356;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_724;
wire n_3753;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_3648;
wire n_2035;
wire n_658;
wire n_2061;
wire n_3773;
wire n_3555;
wire n_3579;
wire n_3918;
wire n_3075;
wire n_3173;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_4317;
wire n_3969;
wire n_2857;
wire n_3932;
wire n_1586;
wire n_4291;
wire n_959;
wire n_2459;
wire n_3031;
wire n_4154;
wire n_535;
wire n_3396;
wire n_3701;
wire n_940;
wire n_4386;
wire n_1445;
wire n_3516;
wire n_4023;
wire n_4149;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1923;
wire n_1773;
wire n_592;
wire n_3243;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_2666;
wire n_2982;
wire n_3385;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_3545;
wire n_2171;
wire n_978;
wire n_2768;
wire n_4299;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_4019;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_3343;
wire n_3515;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_514;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2473;
wire n_3287;
wire n_2137;
wire n_3378;
wire n_603;
wire n_1431;
wire n_2583;
wire n_484;
wire n_1593;
wire n_1033;
wire n_3767;
wire n_4279;
wire n_3426;
wire n_3454;
wire n_2299;
wire n_2873;
wire n_2540;
wire n_3820;
wire n_636;
wire n_4367;
wire n_3741;
wire n_660;
wire n_3410;
wire n_2087;
wire n_1640;
wire n_4294;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_750;
wire n_2029;
wire n_742;
wire n_995;
wire n_3221;
wire n_4125;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_4232;
wire n_3629;
wire n_3021;
wire n_1989;
wire n_3818;
wire n_2359;
wire n_2941;
wire n_3674;
wire n_1887;
wire n_3502;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_3990;
wire n_962;
wire n_3475;
wire n_1215;
wire n_3015;
wire n_4170;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_3719;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_3681;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_3672;
wire n_2399;
wire n_3058;
wire n_4147;
wire n_4308;
wire n_2812;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_3607;
wire n_2355;
wire n_2133;
wire n_4365;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_3830;
wire n_1043;
wire n_2585;
wire n_3505;
wire n_486;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_3730;
wire n_3883;
wire n_1177;
wire n_3276;
wire n_1355;
wire n_2565;
wire n_974;
wire n_4152;
wire n_727;
wire n_3897;
wire n_1159;
wire n_3845;
wire n_957;
wire n_3787;
wire n_773;
wire n_2124;
wire n_743;
wire n_3001;
wire n_2081;
wire n_3945;
wire n_3149;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_3268;
wire n_3597;
wire n_4296;
wire n_2418;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_4281;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_4200;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_3614;
wire n_4198;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_3301;
wire n_4285;
wire n_3466;
wire n_3458;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_3185;
wire n_1132;
wire n_3330;
wire n_1366;
wire n_1300;
wire n_3960;
wire n_2595;
wire n_1127;
wire n_3248;
wire n_2277;
wire n_761;
wire n_2477;
wire n_3523;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_4329;
wire n_1006;
wire n_3411;
wire n_3887;
wire n_4087;
wire n_2110;
wire n_3811;
wire n_4093;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_4271;
wire n_1486;
wire n_582;
wire n_3586;
wire n_1332;
wire n_3519;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_4174;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_1870;
wire n_512;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_4071;
wire n_4330;
wire n_4341;
wire n_4257;
wire n_3453;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_3399;
wire n_4312;
wire n_2896;
wire n_652;
wire n_1111;
wire n_3213;
wire n_1365;
wire n_4074;
wire n_1927;
wire n_3065;
wire n_4361;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_3645;
wire n_609;
wire n_1041;
wire n_1265;
wire n_3223;
wire n_1909;
wire n_3838;
wire n_3929;
wire n_3077;
wire n_4277;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_834;
wire n_3474;
wire n_765;
wire n_4140;
wire n_3675;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_3984;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_3938;
wire n_1913;
wire n_2878;
wire n_504;
wire n_1823;
wire n_511;
wire n_3679;
wire n_3779;
wire n_874;
wire n_2464;
wire n_3422;
wire n_3888;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_4326;
wire n_1456;
wire n_3557;
wire n_2230;
wire n_3498;
wire n_4189;
wire n_2015;
wire n_2365;
wire n_1982;
wire n_1875;
wire n_4110;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_3707;
wire n_987;
wire n_4207;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_4305;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_3429;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_3849;
wire n_3946;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_545;
wire n_860;
wire n_3229;
wire n_4213;
wire n_2849;
wire n_1805;
wire n_3925;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_3692;
wire n_948;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4059;
wire n_2455;
wire n_4349;
wire n_628;
wire n_1849;
wire n_3788;
wire n_4084;
wire n_2410;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_4313;
wire n_970;
wire n_4037;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2467;
wire n_513;
wire n_3366;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_560;
wire n_2288;
wire n_3421;
wire n_4139;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_4063;
wire n_1205;
wire n_1044;
wire n_2436;
wire n_1209;
wire n_3029;
wire n_1552;
wire n_2508;
wire n_3242;
wire n_3592;
wire n_3618;
wire n_4031;
wire n_495;
wire n_602;
wire n_3525;
wire n_574;
wire n_2593;
wire n_3486;
wire n_1435;
wire n_879;
wire n_3394;
wire n_3793;
wire n_3683;
wire n_2416;
wire n_2405;
wire n_3642;
wire n_623;
wire n_3995;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_3808;
wire n_824;
wire n_4339;
wire n_4036;
wire n_1645;
wire n_3881;
wire n_4041;
wire n_2461;
wire n_490;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_4060;
wire n_996;
wire n_1684;
wire n_921;
wire n_2658;
wire n_3590;
wire n_1717;
wire n_572;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_4210;
wire n_2578;
wire n_3097;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_2929;
wire n_3424;
wire n_3478;
wire n_1381;
wire n_2555;
wire n_3751;
wire n_2662;
wire n_2740;
wire n_3824;
wire n_3890;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_3388;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_3583;
wire n_2890;
wire n_3560;
wire n_3059;
wire n_3524;
wire n_4076;
wire n_2554;
wire n_3465;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_3215;
wire n_1438;
wire n_3698;
wire n_3927;
wire n_1082;
wire n_1840;
wire n_589;
wire n_3961;
wire n_1630;
wire n_2122;
wire n_716;
wire n_2512;
wire n_3589;
wire n_4102;
wire n_562;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_3658;
wire n_3449;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_3559;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_3993;
wire n_2216;
wire n_531;
wire n_3020;
wire n_3677;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1424;
wire n_1056;
wire n_960;
wire n_3462;
wire n_3588;
wire n_2933;
wire n_4230;
wire n_2308;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_3419;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_3860;
wire n_1382;
wire n_1029;
wire n_925;
wire n_3546;
wire n_1206;
wire n_4248;
wire n_2647;
wire n_3784;
wire n_3160;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_2969;
wire n_3941;
wire n_3195;
wire n_1519;
wire n_950;
wire n_3190;
wire n_2428;
wire n_1553;
wire n_3678;
wire n_3847;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_3456;
wire n_1346;
wire n_3053;
wire n_1299;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3893;
wire n_3290;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_3298;
wire n_3548;
wire n_968;
wire n_912;
wire n_3569;
wire n_4348;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_3334;
wire n_967;
wire n_1442;
wire n_2923;
wire n_4162;
wire n_3665;
wire n_4355;
wire n_3494;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_2731;
wire n_3264;
wire n_515;
wire n_2333;
wire n_3953;
wire n_885;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_3875;
wire n_3976;
wire n_4122;
wire n_1357;
wire n_483;
wire n_2125;
wire n_3771;
wire n_3979;
wire n_4297;
wire n_683;
wire n_1632;
wire n_3110;
wire n_2998;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_4003;
wire n_3800;
wire n_721;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_4301;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_4048;
wire n_4026;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_983;
wire n_1844;
wire n_4104;
wire n_2760;
wire n_2792;
wire n_3554;
wire n_3377;
wire n_2870;
wire n_3777;
wire n_4377;
wire n_1305;
wire n_3749;
wire n_3178;
wire n_873;
wire n_1826;
wire n_3962;
wire n_3991;
wire n_1112;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_762;
wire n_1283;
wire n_1644;
wire n_4172;
wire n_2334;
wire n_2637;
wire n_4384;
wire n_690;
wire n_4046;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_3537;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_4096;
wire n_4199;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_3750;
wire n_3282;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_3231;
wire n_3105;
wire n_1966;
wire n_3632;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_753;
wire n_621;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_2993;
wire n_4286;
wire n_3864;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_507;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3274;
wire n_3041;
wire n_3299;
wire n_2646;
wire n_1560;
wire n_3715;
wire n_1605;
wire n_4362;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_972;
wire n_3504;
wire n_692;
wire n_2037;
wire n_2685;
wire n_3920;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3568;
wire n_3664;
wire n_2589;
wire n_3203;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_3737;
wire n_3913;
wire n_1185;
wire n_991;
wire n_2903;
wire n_3417;
wire n_3482;
wire n_3921;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_3717;
wire n_4106;
wire n_4034;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_945;
wire n_2997;
wire n_492;
wire n_3743;
wire n_3327;
wire n_1504;
wire n_943;
wire n_3326;
wire n_3956;
wire n_3572;
wire n_992;
wire n_3067;
wire n_4215;
wire n_1932;
wire n_4280;
wire n_3375;
wire n_2755;
wire n_4047;
wire n_543;
wire n_842;
wire n_3734;
wire n_650;
wire n_984;
wire n_694;
wire n_3237;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_3167;
wire n_4239;
wire n_4029;
wire n_3400;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_3423;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_3870;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3574;
wire n_4352;
wire n_918;
wire n_3529;
wire n_3854;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_4201;
wire n_1610;
wire n_4347;
wire n_1077;
wire n_1422;
wire n_3196;
wire n_4095;
wire n_3078;
wire n_2364;
wire n_2533;
wire n_4338;
wire n_540;
wire n_3492;
wire n_618;
wire n_3094;
wire n_896;
wire n_2310;
wire n_2780;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_3099;
wire n_4043;
wire n_3704;
wire n_2596;
wire n_1636;
wire n_894;
wire n_2056;
wire n_3253;
wire n_1730;
wire n_3601;
wire n_3603;
wire n_4027;
wire n_831;
wire n_2280;
wire n_4123;
wire n_2192;
wire n_964;
wire n_3633;
wire n_3363;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_2973;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2318;
wire n_2393;
wire n_3689;
wire n_2020;
wire n_3831;
wire n_1646;
wire n_2502;
wire n_3801;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_2974;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2751;
wire n_2707;
wire n_2793;
wire n_3372;
wire n_3451;
wire n_2971;
wire n_3442;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_3950;
wire n_4000;
wire n_655;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_4121;
wire n_3998;
wire n_1446;
wire n_2285;
wire n_3147;
wire n_2758;
wire n_4141;
wire n_1458;
wire n_669;
wire n_1176;
wire n_1472;
wire n_2471;
wire n_2298;
wire n_1807;
wire n_3869;
wire n_4307;
wire n_1149;
wire n_2618;
wire n_4359;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_3230;
wire n_1020;
wire n_1062;
wire n_3342;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_3386;
wire n_3931;
wire n_3708;
wire n_1204;
wire n_4010;
wire n_4107;
wire n_2840;
wire n_3729;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_3488;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_3861;
wire n_3780;
wire n_1848;
wire n_1928;
wire n_555;
wire n_783;
wire n_2126;
wire n_4117;
wire n_2893;
wire n_3636;
wire n_1188;
wire n_2962;
wire n_2588;
wire n_4004;
wire n_4118;
wire n_1722;
wire n_3957;
wire n_661;
wire n_2441;
wire n_3848;
wire n_1802;
wire n_3083;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_4079;
wire n_3898;
wire n_849;
wire n_2795;
wire n_4091;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2002;
wire n_2282;
wire n_3608;
wire n_510;
wire n_2800;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_3233;
wire n_3829;
wire n_3380;
wire n_3177;
wire n_4053;
wire n_830;
wire n_4274;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_3409;
wire n_3460;
wire n_2352;
wire n_3538;
wire n_1413;
wire n_801;
wire n_4040;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_3552;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_3198;
wire n_749;
wire n_1895;
wire n_3123;
wire n_3684;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_4316;
wire n_939;
wire n_3697;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_3393;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_4247;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_4018;
wire n_4044;
wire n_3900;
wire n_4062;
wire n_4113;
wire n_3520;
wire n_3971;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_3759;
wire n_1338;
wire n_577;
wire n_4005;
wire n_2016;
wire n_1522;
wire n_4321;
wire n_4342;
wire n_3872;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_4336;
wire n_3933;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_3206;
wire n_2653;
wire n_3578;
wire n_3966;
wire n_990;
wire n_836;
wire n_2867;
wire n_3812;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_567;
wire n_1465;
wire n_3145;
wire n_4183;
wire n_3124;
wire n_778;
wire n_1122;
wire n_4068;
wire n_4253;
wire n_4290;
wire n_4233;
wire n_3192;
wire n_2608;
wire n_3877;
wire n_3764;
wire n_2657;
wire n_770;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_3547;
wire n_2649;
wire n_3977;
wire n_1102;
wire n_3727;
wire n_2852;
wire n_3774;
wire n_4052;
wire n_2392;
wire n_3459;
wire n_3093;
wire n_1843;
wire n_1499;
wire n_711;
wire n_3061;
wire n_3155;
wire n_1187;
wire n_3517;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1929;
wire n_1597;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_489;
wire n_1174;
wire n_2431;
wire n_3356;
wire n_3324;
wire n_3758;
wire n_2835;
wire n_3914;
wire n_4304;
wire n_3911;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_3803;
wire n_3182;
wire n_1572;
wire n_1968;
wire n_4192;
wire n_3742;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_1516;
wire n_876;
wire n_3736;
wire n_1190;
wire n_3506;
wire n_3896;
wire n_1736;
wire n_3605;
wire n_1685;
wire n_3958;
wire n_2409;
wire n_601;
wire n_917;
wire n_3450;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_3402;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3565;
wire n_4115;
wire n_726;
wire n_3174;
wire n_982;
wire n_2575;
wire n_2988;
wire n_3390;
wire n_1573;
wire n_1731;
wire n_1453;
wire n_2217;
wire n_3746;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_2766;
wire n_3817;
wire n_1658;
wire n_899;
wire n_1253;
wire n_2722;
wire n_1737;
wire n_2201;
wire n_2745;
wire n_2117;
wire n_3408;
wire n_1904;
wire n_4167;
wire n_2640;
wire n_1993;
wire n_774;
wire n_3835;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_3432;
wire n_1514;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_3967;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_3401;
wire n_1899;
wire n_3226;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_3090;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_3762;
wire n_3902;
wire n_3533;
wire n_2877;
wire n_3318;
wire n_4070;
wire n_2148;
wire n_4282;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_3485;
wire n_4180;
wire n_487;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_665;
wire n_3035;
wire n_3654;
wire n_1440;
wire n_3839;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_910;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_4143;
wire n_4323;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_3972;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_3639;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4105;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_3791;
wire n_4204;
wire n_3308;
wire n_2665;
wire n_3905;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_3368;
wire n_2924;
wire n_3467;
wire n_808;
wire n_2484;
wire n_4111;
wire n_797;
wire n_3530;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_3731;
wire n_2765;
wire n_3329;
wire n_4322;
wire n_500;
wire n_2994;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_3135;
wire n_4354;
wire n_3657;
wire n_2003;
wire n_1457;
wire n_766;
wire n_3928;
wire n_541;
wire n_2692;
wire n_3573;
wire n_3148;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_3534;
wire n_715;
wire n_3901;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3757;
wire n_536;
wire n_3438;
wire n_4098;
wire n_872;
wire n_2012;
wire n_594;
wire n_3792;
wire n_4272;
wire n_1291;
wire n_3974;
wire n_3381;
wire n_3871;
wire n_4094;
wire n_3503;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_1782;
wire n_2245;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_4269;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_2965;
wire n_3536;
wire n_3661;
wire n_3635;
wire n_4150;
wire n_827;
wire n_3217;
wire n_3425;
wire n_3404;
wire n_1703;
wire n_3312;
wire n_4055;
wire n_1352;
wire n_2926;
wire n_626;
wire n_2197;
wire n_2199;
wire n_3540;
wire n_1650;
wire n_3670;
wire n_3973;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3046;
wire n_3882;
wire n_3934;
wire n_2213;
wire n_1170;
wire n_2023;
wire n_3826;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_3922;
wire n_3846;
wire n_676;
wire n_2103;
wire n_653;
wire n_3968;
wire n_2160;
wire n_642;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_3074;
wire n_3204;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_1999;
wire n_664;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_3673;
wire n_2480;
wire n_4017;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_3943;
wire n_1822;
wire n_3397;
wire n_3740;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_4072;
wire n_916;
wire n_1081;
wire n_2549;
wire n_493;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_4380;
wire n_703;
wire n_980;
wire n_1115;
wire n_698;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2977;
wire n_3606;
wire n_2601;
wire n_3043;
wire n_4022;
wire n_998;
wire n_3802;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_3600;
wire n_501;
wire n_823;
wire n_2686;
wire n_2528;
wire n_4134;
wire n_725;
wire n_2344;
wire n_3892;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_4035;
wire n_2316;
wire n_672;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3711;
wire n_3315;
wire n_581;
wire n_2906;
wire n_554;
wire n_1625;
wire n_2130;
wire n_3415;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_3239;
wire n_3139;
wire n_2773;
wire n_3292;
wire n_3172;
wire n_2598;
wire n_3878;
wire n_1762;
wire n_1013;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_1452;
wire n_718;
wire n_2687;
wire n_3023;
wire n_3553;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_4220;
wire n_4251;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_4075;
wire n_4193;
wire n_3982;
wire n_2654;
wire n_997;
wire n_3431;
wire n_3104;
wire n_932;
wire n_3169;
wire n_3151;
wire n_612;
wire n_3822;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_3850;
wire n_788;
wire n_1326;
wire n_3070;
wire n_3284;
wire n_4066;
wire n_3647;
wire n_3176;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_559;
wire n_825;
wire n_4351;
wire n_2819;
wire n_3126;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_4368;
wire n_737;
wire n_1718;
wire n_4050;
wire n_3700;
wire n_3609;
wire n_4136;
wire n_986;
wire n_2315;
wire n_509;
wire n_3228;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_1952;
wire n_4223;
wire n_1281;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1063;
wire n_3720;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_733;
wire n_1922;
wire n_2966;
wire n_4049;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_3862;
wire n_1569;
wire n_2188;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_867;
wire n_2422;
wire n_3959;
wire n_2239;
wire n_587;
wire n_2950;
wire n_792;
wire n_1429;
wire n_756;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_4346;
wire n_3852;
wire n_548;
wire n_3170;
wire n_3724;
wire n_812;
wire n_2104;
wire n_2748;
wire n_3311;
wire n_518;
wire n_505;
wire n_2057;
wire n_3272;
wire n_4008;
wire n_3011;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_4196;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_3345;
wire n_862;
wire n_3584;
wire n_1425;
wire n_760;
wire n_3858;
wire n_1901;
wire n_3069;
wire n_3756;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_3691;
wire n_3628;
wire n_2889;
wire n_4235;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_4382;
wire n_2939;
wire n_1745;
wire n_3924;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_3412;
wire n_3999;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_3807;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2447;
wire n_1813;
wire n_2343;
wire n_3761;
wire n_886;
wire n_3439;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_654;
wire n_1172;
wire n_2535;
wire n_4205;
wire n_1341;
wire n_2774;
wire n_570;
wire n_2726;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_2382;
wire n_1707;
wire n_853;
wire n_4178;
wire n_3062;
wire n_3161;
wire n_2317;
wire n_751;
wire n_3289;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_4229;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_3477;
wire n_3017;
wire n_3626;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_4100;
wire n_4228;
wire n_2456;
wire n_3904;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_522;
wire n_3364;
wire n_1287;
wire n_4363;
wire n_1262;
wire n_2691;
wire n_930;
wire n_4092;
wire n_3908;
wire n_1873;
wire n_1411;
wire n_3926;
wire n_3201;
wire n_3054;
wire n_4335;
wire n_1962;
wire n_622;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2423;
wire n_3671;
wire n_1087;
wire n_3472;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_4181;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_3302;
wire n_3235;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_4225;
wire n_3391;
wire n_682;
wire n_1567;
wire n_4259;
wire n_2567;
wire n_3949;
wire n_3543;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_922;
wire n_3122;
wire n_816;
wire n_1648;
wire n_4015;
wire n_591;
wire n_3842;
wire n_1536;
wire n_3050;
wire n_3265;
wire n_1857;
wire n_4056;
wire n_4153;
wire n_1344;
wire n_2041;
wire n_631;
wire n_3627;
wire n_1246;
wire n_3840;
wire n_4300;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_2957;
wire n_839;
wire n_3551;
wire n_3903;
wire n_1210;
wire n_3518;
wire n_2964;
wire n_3769;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_3733;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_4267;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_3865;
wire n_3722;
wire n_3859;
wire n_4171;
wire n_1842;
wire n_871;
wire n_2442;
wire n_3309;
wire n_3738;
wire n_4045;
wire n_685;
wire n_598;
wire n_928;
wire n_1367;
wire n_608;
wire n_1943;
wire n_3634;
wire n_1460;
wire n_772;
wire n_2018;
wire n_3464;
wire n_3260;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_3245;
wire n_3357;
wire n_499;
wire n_2531;
wire n_1589;
wire n_4116;
wire n_517;
wire n_3428;
wire n_2961;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_3351;
wire n_1619;
wire n_3527;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_3754;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1752;
wire n_1525;
wire n_2397;
wire n_740;
wire n_2883;
wire n_3115;
wire n_4287;
wire n_3509;
wire n_3352;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_4182;
wire n_3063;
wire n_3617;
wire n_2912;
wire n_1794;
wire n_3535;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_3251;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_3955;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4270;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_3118;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_2321;
wire n_3511;
wire n_1226;
wire n_1277;
wire n_722;
wire n_3680;
wire n_2591;
wire n_3443;
wire n_2146;
wire n_844;
wire n_3384;
wire n_852;
wire n_3497;
wire n_1487;
wire n_1864;
wire n_3644;
wire n_1601;
wire n_1028;
wire n_4016;
wire n_3336;
wire n_3935;
wire n_781;
wire n_2940;
wire n_542;
wire n_3435;
wire n_3521;
wire n_3575;
wire n_1546;
wire n_595;
wire n_502;
wire n_3562;
wire n_3948;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_4231;
wire n_979;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3322;
wire n_3232;
wire n_3652;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_3250;
wire n_1937;
wire n_585;
wire n_2112;
wire n_4083;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_616;
wire n_2278;
wire n_2594;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3234;
wire n_1914;
wire n_3612;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_3493;
wire n_745;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_4328;
wire n_3004;
wire n_3323;
wire n_3916;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_4081;
wire n_3132;
wire n_3556;
wire n_648;
wire n_1379;
wire n_2734;
wire n_3874;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3951;
wire n_3024;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_3512;
wire n_494;
wire n_1761;
wire n_641;
wire n_3238;
wire n_3210;
wire n_3930;
wire n_730;
wire n_3175;
wire n_3522;
wire n_2036;
wire n_1325;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_575;
wire n_795;
wire n_2404;
wire n_4345;
wire n_2083;
wire n_695;
wire n_3281;
wire n_656;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_3964;
wire n_3266;
wire n_2485;
wire n_4318;
wire n_3772;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_3884;
wire n_4185;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_3726;
wire n_2210;
wire n_4169;
wire n_805;
wire n_3247;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_2525;
wire n_2513;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_3480;
wire n_2892;
wire n_4032;
wire n_3057;
wire n_3194;
wire n_3582;
wire n_3066;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_3577;
wire n_3539;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_3662;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_4319;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_657;
wire n_4320;
wire n_644;
wire n_1741;
wire n_2229;
wire n_4124;
wire n_1160;
wire n_1397;
wire n_4057;
wire n_4332;
wire n_491;
wire n_1258;
wire n_4314;
wire n_1074;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_1621;
wire n_2708;
wire n_3809;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_3694;
wire n_1448;
wire n_4245;
wire n_4288;
wire n_4364;
wire n_2225;
wire n_3613;
wire n_3567;
wire n_1507;
wire n_4378;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3444;
wire n_3853;
wire n_1181;
wire n_1505;
wire n_4216;
wire n_4222;
wire n_1634;
wire n_3939;
wire n_1196;
wire n_4012;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_811;
wire n_1558;
wire n_3225;
wire n_4241;
wire n_807;
wire n_3321;
wire n_2166;
wire n_3910;
wire n_2938;
wire n_3212;
wire n_835;
wire n_666;
wire n_3319;
wire n_3594;
wire n_1433;
wire n_4309;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_3721;
wire n_3335;
wire n_1254;
wire n_3799;
wire n_4119;
wire n_4298;
wire n_1026;
wire n_3413;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_2044;
wire n_2013;
wire n_1089;
wire n_1990;
wire n_927;
wire n_2920;
wire n_2689;
wire n_3259;
wire n_4265;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_4191;
wire n_2511;
wire n_4293;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_3688;
wire n_3383;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_3585;
wire n_2975;
wire n_3473;
wire n_4188;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_4214;
wire n_1622;
wire n_2237;
wire n_3414;
wire n_3463;
wire n_3699;
wire n_1180;
wire n_1827;
wire n_3360;
wire n_4209;
wire n_2524;
wire n_3873;
wire n_1271;
wire n_3705;
wire n_2802;
wire n_533;
wire n_1542;
wire n_1251;
wire n_3693;
wire n_4366;
wire n_4009;
wire n_3159;
wire n_2728;
wire n_3857;
wire n_2268;
wire n_3778;

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_256),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_13),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_390),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_41),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_439),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_278),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_135),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_407),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_61),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_289),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_309),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_166),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_326),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_27),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_43),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_110),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_93),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_225),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_38),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_167),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_14),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_481),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_257),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_356),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_4),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_233),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_30),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_421),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_283),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_213),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_51),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_139),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_336),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_102),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_94),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_20),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_469),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_267),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g521 ( 
.A(n_88),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_363),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_75),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_126),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_114),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_339),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_51),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_91),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_171),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_329),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_134),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_328),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_225),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_206),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_185),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_291),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_449),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_3),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_482),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_31),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_340),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_73),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_35),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_145),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_81),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_313),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_59),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_48),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_65),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_142),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_114),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_330),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_268),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_59),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_8),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_256),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_89),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_130),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_288),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_6),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_164),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_400),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_306),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_416),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_315),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_180),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_23),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_165),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_110),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_362),
.Y(n_570)
);

BUFx10_ASAP7_75t_L g571 ( 
.A(n_170),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_317),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_75),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_151),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_172),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_109),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_465),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_234),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_217),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g580 ( 
.A(n_472),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_480),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_358),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_291),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_106),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_289),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_109),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_467),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_207),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_160),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_113),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_447),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_397),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_377),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_134),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_153),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_16),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_389),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_24),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_77),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_258),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_107),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_165),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_267),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_413),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_364),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_212),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_329),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_268),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_387),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_434),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_331),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_399),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_314),
.Y(n_613)
);

BUFx2_ASAP7_75t_SL g614 ( 
.A(n_196),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_60),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_215),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_361),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_235),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_348),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_45),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_426),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_100),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_324),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_411),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_325),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_257),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_9),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_143),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_23),
.Y(n_629)
);

BUFx10_ASAP7_75t_L g630 ( 
.A(n_50),
.Y(n_630)
);

BUFx10_ASAP7_75t_L g631 ( 
.A(n_318),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_104),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_452),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_83),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_409),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_272),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_133),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_433),
.Y(n_638)
);

CKINVDCx16_ASAP7_75t_R g639 ( 
.A(n_220),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_405),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_315),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_238),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_349),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_342),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_94),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_476),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_64),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_130),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_290),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_148),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_88),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_125),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_121),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_332),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_450),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_420),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_286),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_34),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_77),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_319),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_406),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_331),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_378),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_16),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_248),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_334),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_320),
.Y(n_667)
);

CKINVDCx14_ASAP7_75t_R g668 ( 
.A(n_344),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_349),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_292),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_95),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_95),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_276),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_150),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_375),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_356),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_140),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_228),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_401),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_415),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_260),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_334),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_212),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_38),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_137),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_326),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_264),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_343),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_136),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_115),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_432),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_173),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_281),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_197),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_72),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_200),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_359),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_86),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_166),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_91),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_380),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_269),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_242),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_321),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_479),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_442),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_231),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_383),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_194),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_215),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_316),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_86),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_163),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_299),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_7),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_40),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_443),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_170),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_211),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_466),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_330),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_198),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_101),
.Y(n_723)
);

BUFx10_ASAP7_75t_L g724 ( 
.A(n_337),
.Y(n_724)
);

BUFx2_ASAP7_75t_SL g725 ( 
.A(n_66),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_151),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_50),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_31),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_8),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_79),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_200),
.Y(n_731)
);

CKINVDCx16_ASAP7_75t_R g732 ( 
.A(n_226),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_155),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_393),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_408),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_156),
.Y(n_736)
);

CKINVDCx16_ASAP7_75t_R g737 ( 
.A(n_169),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_463),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_197),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_214),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_29),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_328),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_459),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_159),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_111),
.Y(n_745)
);

CKINVDCx14_ASAP7_75t_R g746 ( 
.A(n_398),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_237),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_318),
.Y(n_748)
);

BUFx10_ASAP7_75t_L g749 ( 
.A(n_4),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_20),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_97),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_402),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_457),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_446),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_19),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_24),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_232),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_430),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_58),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_27),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_173),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_388),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_273),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_392),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_117),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_63),
.Y(n_766)
);

CKINVDCx16_ASAP7_75t_R g767 ( 
.A(n_213),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_347),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_144),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_322),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_141),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_303),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_266),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_0),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_385),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_346),
.Y(n_776)
);

BUFx10_ASAP7_75t_L g777 ( 
.A(n_32),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_270),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_160),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_49),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_423),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_108),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_118),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_353),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_185),
.Y(n_785)
);

CKINVDCx16_ASAP7_75t_R g786 ( 
.A(n_182),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_111),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_128),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_499),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_564),
.Y(n_790)
);

INVxp33_ASAP7_75t_L g791 ( 
.A(n_629),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_499),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_519),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_499),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_624),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_499),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_485),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_499),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_541),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_499),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_668),
.B(n_640),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_487),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_541),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_497),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_497),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_580),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_524),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_497),
.Y(n_808)
);

CKINVDCx16_ASAP7_75t_R g809 ( 
.A(n_639),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_538),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_538),
.Y(n_811)
);

CKINVDCx20_ASAP7_75t_R g812 ( 
.A(n_580),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_538),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_746),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_546),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_519),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_682),
.Y(n_817)
);

INVxp67_ASAP7_75t_SL g818 ( 
.A(n_524),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_546),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_490),
.Y(n_820)
);

CKINVDCx14_ASAP7_75t_R g821 ( 
.A(n_682),
.Y(n_821)
);

INVxp33_ASAP7_75t_SL g822 ( 
.A(n_703),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_546),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_585),
.Y(n_824)
);

INVxp67_ASAP7_75t_SL g825 ( 
.A(n_524),
.Y(n_825)
);

INVxp67_ASAP7_75t_SL g826 ( 
.A(n_542),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_585),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_585),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_588),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_504),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_588),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_588),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_510),
.Y(n_833)
);

CKINVDCx16_ASAP7_75t_R g834 ( 
.A(n_639),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_607),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_607),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_607),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_522),
.Y(n_838)
);

INVxp67_ASAP7_75t_SL g839 ( 
.A(n_542),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_636),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_537),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_636),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_636),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_570),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_642),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_642),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_581),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_642),
.Y(n_848)
);

INVxp33_ASAP7_75t_SL g849 ( 
.A(n_703),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_591),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_688),
.Y(n_851)
);

INVx1_ASAP7_75t_SL g852 ( 
.A(n_778),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_593),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_688),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_597),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_522),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_778),
.Y(n_857)
);

INVxp67_ASAP7_75t_SL g858 ( 
.A(n_542),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_539),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_539),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_562),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_562),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_577),
.Y(n_863)
);

INVxp67_ASAP7_75t_SL g864 ( 
.A(n_577),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_688),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_609),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_740),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_740),
.Y(n_868)
);

CKINVDCx14_ASAP7_75t_R g869 ( 
.A(n_571),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_740),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_780),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_780),
.Y(n_872)
);

CKINVDCx14_ASAP7_75t_R g873 ( 
.A(n_571),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_610),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_571),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_614),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_780),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_732),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_732),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_484),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_646),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_484),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_587),
.Y(n_883)
);

INVxp67_ASAP7_75t_SL g884 ( 
.A(n_587),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_663),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_489),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_489),
.Y(n_887)
);

INVxp67_ASAP7_75t_SL g888 ( 
.A(n_592),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_737),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_493),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_655),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_493),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_496),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_496),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_656),
.Y(n_895)
);

INVxp67_ASAP7_75t_SL g896 ( 
.A(n_592),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_675),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_691),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_498),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_498),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_501),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_501),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_604),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_701),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_604),
.Y(n_905)
);

NAND2xp33_ASAP7_75t_R g906 ( 
.A(n_708),
.B(n_0),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_506),
.Y(n_907)
);

INVx1_ASAP7_75t_SL g908 ( 
.A(n_509),
.Y(n_908)
);

INVxp67_ASAP7_75t_L g909 ( 
.A(n_614),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_506),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_511),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_511),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_514),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_514),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_527),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_605),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_527),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_640),
.B(n_605),
.Y(n_918)
);

BUFx5_ASAP7_75t_L g919 ( 
.A(n_612),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_529),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_529),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_612),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_533),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_533),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_535),
.Y(n_925)
);

INVxp33_ASAP7_75t_SL g926 ( 
.A(n_483),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_535),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_717),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_551),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_551),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_735),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_558),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_753),
.Y(n_933)
);

INVxp67_ASAP7_75t_SL g934 ( 
.A(n_617),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_558),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_663),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_754),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_559),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_818),
.B(n_670),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_822),
.A2(n_767),
.B1(n_786),
.B2(n_737),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_789),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_821),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_789),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_797),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_792),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_825),
.B(n_670),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_796),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_796),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_936),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_936),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_809),
.B(n_767),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_849),
.A2(n_786),
.B1(n_526),
.B2(n_528),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_792),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_936),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_794),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_936),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_826),
.B(n_712),
.Y(n_957)
);

BUFx12f_ASAP7_75t_L g958 ( 
.A(n_802),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_926),
.B(n_582),
.Y(n_959)
);

NOR2x1_ASAP7_75t_L g960 ( 
.A(n_885),
.B(n_663),
.Y(n_960)
);

CKINVDCx20_ASAP7_75t_R g961 ( 
.A(n_790),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_839),
.B(n_712),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_936),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_794),
.Y(n_964)
);

BUFx12f_ASAP7_75t_L g965 ( 
.A(n_820),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_798),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_798),
.Y(n_967)
);

BUFx8_ASAP7_75t_L g968 ( 
.A(n_889),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_800),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_800),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_811),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_811),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_819),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_819),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_829),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_829),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_842),
.Y(n_977)
);

BUFx8_ASAP7_75t_L g978 ( 
.A(n_889),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_864),
.B(n_752),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_806),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_842),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_884),
.B(n_888),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_896),
.B(n_752),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_878),
.Y(n_984)
);

CKINVDCx6p67_ASAP7_75t_R g985 ( 
.A(n_814),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_830),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_845),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_845),
.Y(n_988)
);

OA21x2_ASAP7_75t_L g989 ( 
.A1(n_804),
.A2(n_621),
.B(n_617),
.Y(n_989)
);

INVx4_ASAP7_75t_L g990 ( 
.A(n_885),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_804),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_805),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_885),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_879),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_805),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_808),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_852),
.A2(n_601),
.B1(n_556),
.B2(n_488),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_919),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_812),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_834),
.A2(n_531),
.B1(n_573),
.B2(n_517),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_880),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_833),
.B(n_758),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_919),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_799),
.A2(n_653),
.B1(n_657),
.B2(n_615),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_880),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_817),
.A2(n_491),
.B1(n_492),
.B2(n_486),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_841),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_919),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_808),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_908),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_807),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_844),
.Y(n_1012)
);

BUFx8_ASAP7_75t_L g1013 ( 
.A(n_803),
.Y(n_1013)
);

AND2x6_ASAP7_75t_L g1014 ( 
.A(n_918),
.B(n_752),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_810),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_810),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_813),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_813),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_803),
.A2(n_692),
.B1(n_696),
.B2(n_658),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_SL g1020 ( 
.A(n_875),
.B(n_582),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_SL g1021 ( 
.A1(n_795),
.A2(n_750),
.B1(n_760),
.B2(n_726),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_882),
.Y(n_1022)
);

OA21x2_ASAP7_75t_L g1023 ( 
.A1(n_815),
.A2(n_633),
.B(n_621),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_815),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_823),
.Y(n_1025)
);

INVx5_ASAP7_75t_L g1026 ( 
.A(n_793),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_791),
.A2(n_495),
.B1(n_500),
.B2(n_494),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_823),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_824),
.Y(n_1029)
);

INVx5_ASAP7_75t_L g1030 ( 
.A(n_793),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_824),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_875),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_858),
.B(n_771),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_827),
.Y(n_1034)
);

INVx6_ASAP7_75t_L g1035 ( 
.A(n_816),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_847),
.B(n_781),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_934),
.B(n_633),
.Y(n_1037)
);

INVx5_ASAP7_75t_L g1038 ( 
.A(n_816),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_827),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_828),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_882),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_807),
.B(n_771),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_850),
.B(n_635),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_919),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_828),
.Y(n_1045)
);

AND2x6_ASAP7_75t_L g1046 ( 
.A(n_801),
.B(n_775),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_886),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_SL g1048 ( 
.A1(n_869),
.A2(n_768),
.B1(n_623),
.B2(n_654),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_838),
.B(n_559),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_886),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_838),
.B(n_563),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_855),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_881),
.B(n_635),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_831),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_891),
.B(n_638),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_831),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_887),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_887),
.Y(n_1058)
);

BUFx12f_ASAP7_75t_L g1059 ( 
.A(n_895),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_883),
.B(n_638),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_857),
.A2(n_534),
.B1(n_654),
.B2(n_623),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_873),
.Y(n_1062)
);

BUFx8_ASAP7_75t_L g1063 ( 
.A(n_856),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_972),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_947),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_950),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_947),
.Y(n_1067)
);

NAND2x1_ASAP7_75t_L g1068 ( 
.A(n_990),
.B(n_1014),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_950),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_972),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_972),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_982),
.B(n_904),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_947),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_982),
.B(n_928),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_972),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_941),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_941),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_SL g1078 ( 
.A1(n_1021),
.A2(n_684),
.B1(n_685),
.B2(n_534),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_972),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_950),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_972),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_943),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_943),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_945),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_945),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_953),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_982),
.B(n_931),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_953),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_950),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_950),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_955),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_975),
.Y(n_1092)
);

XOR2xp5_ASAP7_75t_L g1093 ( 
.A(n_1021),
.B(n_853),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_982),
.B(n_937),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_1010),
.Y(n_1095)
);

NAND2xp33_ASAP7_75t_SL g1096 ( 
.A(n_1032),
.B(n_866),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1046),
.B(n_919),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1046),
.B(n_919),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_955),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1042),
.B(n_883),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_966),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_975),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_1020),
.B(n_959),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_975),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_966),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_1032),
.B(n_874),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_969),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_969),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_975),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_970),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_950),
.Y(n_1111)
);

INVx4_ASAP7_75t_L g1112 ( 
.A(n_993),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_970),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_975),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1042),
.B(n_916),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1037),
.B(n_916),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_975),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1001),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1046),
.B(n_919),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1043),
.B(n_897),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_956),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1001),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1005),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_994),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1005),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_977),
.Y(n_1126)
);

BUFx8_ASAP7_75t_L g1127 ( 
.A(n_1062),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_942),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_977),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_956),
.Y(n_1130)
);

NAND2x1p5_ASAP7_75t_L g1131 ( 
.A(n_989),
.B(n_705),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1022),
.Y(n_1132)
);

NOR2x1_ASAP7_75t_L g1133 ( 
.A(n_1002),
.B(n_661),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_956),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1022),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1062),
.B(n_898),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1041),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1041),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1047),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_SL g1140 ( 
.A(n_958),
.B(n_933),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1047),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1050),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_977),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_956),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_977),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1050),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1057),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_977),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_977),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1046),
.B(n_919),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1057),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1058),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_987),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_987),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_961),
.Y(n_1155)
);

INVxp67_ASAP7_75t_L g1156 ( 
.A(n_1027),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_984),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_987),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1046),
.B(n_919),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_1011),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_956),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1058),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_944),
.B(n_986),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_948),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_987),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1013),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_948),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_980),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_987),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_987),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_964),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1053),
.A2(n_860),
.B(n_859),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_964),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1046),
.B(n_861),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1037),
.B(n_939),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_967),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_956),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1007),
.B(n_876),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1046),
.B(n_862),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1037),
.B(n_922),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1037),
.B(n_922),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_967),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1055),
.B(n_863),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_990),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_993),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_990),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_990),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_949),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_949),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1060),
.B(n_661),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_993),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_940),
.A2(n_906),
.B1(n_684),
.B2(n_707),
.Y(n_1192)
);

INVx6_ASAP7_75t_L g1193 ( 
.A(n_1026),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_993),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_954),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_993),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_954),
.Y(n_1197)
);

INVxp67_ASAP7_75t_L g1198 ( 
.A(n_951),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_963),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_993),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_995),
.Y(n_1201)
);

INVx5_ASAP7_75t_L g1202 ( 
.A(n_1014),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_979),
.B(n_903),
.Y(n_1203)
);

INVx4_ASAP7_75t_L g1204 ( 
.A(n_995),
.Y(n_1204)
);

OA21x2_ASAP7_75t_L g1205 ( 
.A1(n_963),
.A2(n_905),
.B(n_835),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_995),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_995),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_979),
.B(n_705),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_989),
.Y(n_1209)
);

INVxp67_ASAP7_75t_L g1210 ( 
.A(n_1006),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_989),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1060),
.B(n_679),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_989),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1023),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_979),
.B(n_706),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_995),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1023),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_995),
.Y(n_1218)
);

INVx1_ASAP7_75t_SL g1219 ( 
.A(n_980),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1023),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1023),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_996),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_974),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_998),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_996),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_974),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_996),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_981),
.Y(n_1228)
);

CKINVDCx8_ASAP7_75t_R g1229 ( 
.A(n_999),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_1035),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_996),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_981),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_996),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1049),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_996),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1009),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1052),
.B(n_1063),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1009),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1009),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1009),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1009),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1060),
.B(n_979),
.Y(n_1242)
);

AND2x2_ASAP7_75t_SL g1243 ( 
.A(n_983),
.B(n_679),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_939),
.B(n_832),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_998),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1009),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1015),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1035),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1015),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_998),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1015),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1015),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1015),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1015),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1024),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1024),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1024),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1024),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_946),
.B(n_832),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1024),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1011),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1024),
.Y(n_1262)
);

BUFx8_ASAP7_75t_L g1263 ( 
.A(n_999),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1025),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1060),
.B(n_680),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1025),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1025),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1003),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1049),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_1051),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_983),
.B(n_680),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1025),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1025),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1025),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1039),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1039),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_983),
.B(n_706),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1039),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1039),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_946),
.B(n_835),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1039),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_983),
.B(n_764),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1039),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1014),
.B(n_1036),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1040),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_971),
.A2(n_837),
.B(n_836),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1040),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1040),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1040),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1242),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1243),
.B(n_1175),
.Y(n_1291)
);

BUFx10_ASAP7_75t_L g1292 ( 
.A(n_1120),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1103),
.B(n_1072),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1074),
.B(n_1063),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1156),
.A2(n_957),
.B1(n_1033),
.B2(n_962),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1205),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1205),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1230),
.Y(n_1298)
);

OR2x6_ASAP7_75t_L g1299 ( 
.A(n_1166),
.B(n_958),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1243),
.A2(n_1014),
.B1(n_962),
.B2(n_957),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1243),
.B(n_1014),
.Y(n_1301)
);

NAND3x1_ASAP7_75t_L g1302 ( 
.A(n_1192),
.B(n_952),
.C(n_1019),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1205),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1087),
.B(n_1012),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1242),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1175),
.B(n_1014),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1095),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1242),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1094),
.B(n_1198),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1242),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1133),
.B(n_1014),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1210),
.B(n_965),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1133),
.B(n_1033),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1095),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1116),
.B(n_1180),
.Y(n_1315)
);

INVx6_ASAP7_75t_L g1316 ( 
.A(n_1112),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_1234),
.B(n_952),
.C(n_1063),
.Y(n_1317)
);

INVx4_ASAP7_75t_L g1318 ( 
.A(n_1207),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1205),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1065),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1286),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1230),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1100),
.B(n_1115),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1208),
.B(n_1063),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1248),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1271),
.A2(n_697),
.B1(n_734),
.B2(n_720),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1286),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1215),
.A2(n_764),
.B1(n_697),
.B2(n_734),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1271),
.A2(n_1212),
.B1(n_1265),
.B2(n_1190),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1065),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1068),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1067),
.Y(n_1332)
);

INVx5_ASAP7_75t_L g1333 ( 
.A(n_1193),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1271),
.A2(n_1212),
.B1(n_1265),
.B2(n_1190),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1277),
.B(n_965),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1286),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1282),
.B(n_1059),
.Y(n_1337)
);

BUFx10_ASAP7_75t_L g1338 ( 
.A(n_1271),
.Y(n_1338)
);

OAI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1192),
.A2(n_1004),
.B1(n_1061),
.B2(n_1019),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1286),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1157),
.B(n_1059),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1116),
.B(n_1035),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1067),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1073),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1180),
.B(n_1013),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1181),
.B(n_1035),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1076),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_1068),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1076),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1073),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1248),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1077),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1077),
.Y(n_1353)
);

AND2x6_ASAP7_75t_L g1354 ( 
.A(n_1209),
.B(n_720),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1181),
.B(n_1003),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1224),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1082),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1155),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1100),
.B(n_1051),
.Y(n_1359)
);

INVx4_ASAP7_75t_L g1360 ( 
.A(n_1207),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1224),
.Y(n_1361)
);

NAND2xp33_ASAP7_75t_L g1362 ( 
.A(n_1202),
.B(n_1131),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1118),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1118),
.Y(n_1364)
);

INVx5_ASAP7_75t_L g1365 ( 
.A(n_1193),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1115),
.B(n_909),
.Y(n_1366)
);

AND2x6_ASAP7_75t_L g1367 ( 
.A(n_1209),
.B(n_738),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1168),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1082),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1127),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1124),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1083),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_1219),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1083),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1080),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1084),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1184),
.B(n_1003),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_SL g1378 ( 
.A(n_1160),
.B(n_1013),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1084),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1244),
.B(n_1061),
.Y(n_1380)
);

NAND2xp33_ASAP7_75t_L g1381 ( 
.A(n_1202),
.B(n_738),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1261),
.B(n_1013),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1224),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1085),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1184),
.B(n_1008),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1183),
.B(n_1048),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1085),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1086),
.Y(n_1388)
);

BUFx4f_ASAP7_75t_L g1389 ( 
.A(n_1190),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1269),
.B(n_1004),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1122),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1127),
.Y(n_1392)
);

AND2x6_ASAP7_75t_L g1393 ( 
.A(n_1211),
.B(n_743),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1270),
.A2(n_743),
.B1(n_775),
.B2(n_762),
.Y(n_1394)
);

NAND2xp33_ASAP7_75t_L g1395 ( 
.A(n_1202),
.B(n_762),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1080),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1244),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1202),
.B(n_1026),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1086),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1088),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1088),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1186),
.B(n_1008),
.Y(n_1402)
);

INVx4_ASAP7_75t_SL g1403 ( 
.A(n_1211),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1186),
.B(n_1008),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1187),
.B(n_1044),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_SL g1406 ( 
.A(n_1166),
.B(n_985),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1091),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1224),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1096),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1091),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1099),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1178),
.B(n_1048),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1099),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1106),
.B(n_1000),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1203),
.B(n_997),
.C(n_1000),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1190),
.B(n_890),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1187),
.B(n_1044),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1101),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1101),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1259),
.Y(n_1420)
);

AND2x6_ASAP7_75t_L g1421 ( 
.A(n_1213),
.B(n_563),
.Y(n_1421)
);

NAND2x1p5_ASAP7_75t_L g1422 ( 
.A(n_1202),
.B(n_960),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1259),
.B(n_1017),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1202),
.B(n_1030),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1105),
.Y(n_1425)
);

AO22x2_ASAP7_75t_L g1426 ( 
.A1(n_1093),
.A2(n_725),
.B1(n_707),
.B2(n_710),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1127),
.Y(n_1427)
);

NOR3xp33_ASAP7_75t_L g1428 ( 
.A(n_1078),
.B(n_521),
.C(n_685),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1080),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1105),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1280),
.B(n_1044),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1280),
.B(n_1026),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1107),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1107),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1212),
.B(n_890),
.Y(n_1435)
);

BUFx10_ASAP7_75t_L g1436 ( 
.A(n_1212),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_SL g1437 ( 
.A(n_1140),
.B(n_985),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1207),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1108),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1108),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_SL g1441 ( 
.A(n_1265),
.B(n_1026),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1245),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1122),
.B(n_1017),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1123),
.B(n_1026),
.Y(n_1444)
);

BUFx10_ASAP7_75t_L g1445 ( 
.A(n_1265),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1110),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1284),
.B(n_1026),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1128),
.B(n_968),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1123),
.B(n_1125),
.Y(n_1449)
);

INVx4_ASAP7_75t_L g1450 ( 
.A(n_1207),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1125),
.B(n_968),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1110),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1132),
.B(n_1030),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1132),
.B(n_1030),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_SL g1455 ( 
.A(n_1135),
.B(n_1030),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1113),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1263),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1113),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1223),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1136),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1135),
.B(n_1137),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1223),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1226),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1093),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1137),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1138),
.Y(n_1466)
);

NAND2xp33_ASAP7_75t_L g1467 ( 
.A(n_1131),
.B(n_960),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1226),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1138),
.Y(n_1469)
);

NAND2xp33_ASAP7_75t_L g1470 ( 
.A(n_1131),
.B(n_1030),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1229),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1139),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1228),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1213),
.A2(n_725),
.B1(n_1045),
.B2(n_1040),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1228),
.Y(n_1475)
);

INVx4_ASAP7_75t_L g1476 ( 
.A(n_1207),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1245),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1232),
.Y(n_1478)
);

INVx4_ASAP7_75t_L g1479 ( 
.A(n_1216),
.Y(n_1479)
);

INVxp67_ASAP7_75t_SL g1480 ( 
.A(n_1245),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1139),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1127),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1141),
.B(n_1017),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1080),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1141),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1232),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1142),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1142),
.B(n_1030),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1245),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1146),
.Y(n_1490)
);

INVx4_ASAP7_75t_SL g1491 ( 
.A(n_1214),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1146),
.B(n_1038),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1171),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1147),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1147),
.B(n_1038),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1151),
.B(n_968),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1080),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1151),
.B(n_1038),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1121),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1152),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1152),
.B(n_1038),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1162),
.Y(n_1502)
);

INVx4_ASAP7_75t_L g1503 ( 
.A(n_1216),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1162),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1164),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_SL g1506 ( 
.A(n_1174),
.B(n_1038),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_1179),
.B(n_1038),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1164),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1250),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1250),
.B(n_1017),
.Y(n_1510)
);

CKINVDCx20_ASAP7_75t_R g1511 ( 
.A(n_1229),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_R g1512 ( 
.A(n_1263),
.B(n_968),
.Y(n_1512)
);

BUFx10_ASAP7_75t_L g1513 ( 
.A(n_1214),
.Y(n_1513)
);

NAND3xp33_ASAP7_75t_L g1514 ( 
.A(n_1163),
.B(n_978),
.C(n_503),
.Y(n_1514)
);

NAND3xp33_ASAP7_75t_L g1515 ( 
.A(n_1237),
.B(n_978),
.C(n_505),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1167),
.Y(n_1516)
);

INVx4_ASAP7_75t_L g1517 ( 
.A(n_1216),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1078),
.B(n_710),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1167),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1172),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1171),
.Y(n_1521)
);

INVx4_ASAP7_75t_SL g1522 ( 
.A(n_1217),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1188),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1172),
.Y(n_1524)
);

INVx4_ASAP7_75t_L g1525 ( 
.A(n_1216),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1217),
.B(n_1220),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1220),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1097),
.B(n_978),
.Y(n_1528)
);

AND2x2_ASAP7_75t_SL g1529 ( 
.A(n_1221),
.B(n_567),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1182),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1182),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1250),
.B(n_1018),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1173),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1173),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1293),
.B(n_1250),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1313),
.B(n_1268),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1315),
.B(n_1268),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1347),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1320),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1320),
.Y(n_1540)
);

INVx4_ASAP7_75t_L g1541 ( 
.A(n_1290),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1423),
.B(n_1268),
.Y(n_1542)
);

INVxp67_ASAP7_75t_L g1543 ( 
.A(n_1307),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1291),
.B(n_1331),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1309),
.B(n_1304),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1366),
.B(n_718),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1386),
.A2(n_1221),
.B1(n_1176),
.B2(n_1268),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1366),
.B(n_718),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1423),
.B(n_1194),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1347),
.Y(n_1550)
);

NAND2xp33_ASAP7_75t_SL g1551 ( 
.A(n_1331),
.B(n_1098),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1330),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1331),
.B(n_1119),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1397),
.B(n_1200),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1331),
.B(n_1150),
.Y(n_1555)
);

AND2x6_ASAP7_75t_SL g1556 ( 
.A(n_1412),
.B(n_567),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1330),
.Y(n_1557)
);

AND2x4_ASAP7_75t_SL g1558 ( 
.A(n_1338),
.B(n_571),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1323),
.B(n_774),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1368),
.B(n_1373),
.Y(n_1560)
);

NAND2x1p5_ASAP7_75t_L g1561 ( 
.A(n_1290),
.B(n_1194),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1349),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1292),
.B(n_978),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1397),
.B(n_1194),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1349),
.Y(n_1565)
);

NAND2x1p5_ASAP7_75t_L g1566 ( 
.A(n_1290),
.B(n_1194),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1420),
.B(n_1196),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1332),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1420),
.B(n_1196),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_SL g1570 ( 
.A(n_1370),
.Y(n_1570)
);

AND2x6_ASAP7_75t_SL g1571 ( 
.A(n_1341),
.B(n_1312),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1529),
.A2(n_1421),
.B1(n_1300),
.B2(n_1306),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1323),
.B(n_1196),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1526),
.B(n_1352),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1332),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1331),
.B(n_1159),
.Y(n_1576)
);

NAND3xp33_ASAP7_75t_L g1577 ( 
.A(n_1415),
.B(n_1263),
.C(n_507),
.Y(n_1577)
);

NAND2xp33_ASAP7_75t_L g1578 ( 
.A(n_1301),
.B(n_1185),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1305),
.A2(n_1235),
.B1(n_1241),
.B2(n_1236),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1369),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1529),
.A2(n_1176),
.B1(n_1189),
.B2(n_1188),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1369),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1526),
.B(n_1196),
.Y(n_1583)
);

BUFx6f_ASAP7_75t_L g1584 ( 
.A(n_1375),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1352),
.B(n_1200),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1372),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1380),
.B(n_774),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1353),
.B(n_1200),
.Y(n_1588)
);

BUFx5_ASAP7_75t_L g1589 ( 
.A(n_1297),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1389),
.B(n_1348),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1380),
.B(n_630),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1343),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1353),
.B(n_1200),
.Y(n_1593)
);

A2O1A1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1295),
.A2(n_579),
.B(n_594),
.C(n_576),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1357),
.B(n_1189),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1389),
.B(n_1201),
.Y(n_1596)
);

O2A1O1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1328),
.A2(n_1197),
.B(n_1199),
.C(n_1195),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1372),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1292),
.B(n_1263),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1292),
.B(n_1112),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1348),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1314),
.B(n_1112),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1308),
.A2(n_1279),
.B1(n_1283),
.B2(n_1276),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1389),
.B(n_1201),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1470),
.A2(n_1204),
.B(n_1112),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1359),
.B(n_630),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1371),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1329),
.A2(n_1197),
.B1(n_1199),
.B2(n_1195),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1357),
.B(n_1066),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1371),
.B(n_502),
.Y(n_1610)
);

INVx8_ASAP7_75t_L g1611 ( 
.A(n_1421),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1374),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1374),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1348),
.Y(n_1614)
);

O2A1O1Ixp33_ASAP7_75t_L g1615 ( 
.A1(n_1394),
.A2(n_579),
.B(n_594),
.C(n_576),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1403),
.B(n_1206),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1376),
.Y(n_1617)
);

INVxp67_ASAP7_75t_SL g1618 ( 
.A(n_1375),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1376),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1400),
.B(n_1066),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1400),
.B(n_1066),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1401),
.B(n_1410),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1513),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1343),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1403),
.B(n_1491),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1401),
.B(n_1066),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1403),
.B(n_1206),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1344),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1403),
.B(n_1222),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1379),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1410),
.B(n_1111),
.Y(n_1631)
);

NOR2xp67_ASAP7_75t_L g1632 ( 
.A(n_1515),
.B(n_1222),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1344),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1434),
.B(n_1111),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1434),
.B(n_1111),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1460),
.B(n_1390),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1491),
.B(n_1225),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1439),
.B(n_1111),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1491),
.B(n_1225),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1439),
.B(n_1440),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1491),
.B(n_1227),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1440),
.B(n_1130),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1350),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1379),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1310),
.B(n_1064),
.Y(n_1645)
);

AOI22x1_ASAP7_75t_L g1646 ( 
.A1(n_1350),
.A2(n_1070),
.B1(n_1071),
.B2(n_1064),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1446),
.B(n_1130),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1513),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1421),
.A2(n_1236),
.B1(n_1241),
.B2(n_1235),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1384),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1384),
.Y(n_1651)
);

A2O1A1Ixp33_ASAP7_75t_L g1652 ( 
.A1(n_1446),
.A2(n_603),
.B(n_611),
.C(n_600),
.Y(n_1652)
);

AOI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1334),
.A2(n_1342),
.B1(n_1346),
.B2(n_1359),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1527),
.A2(n_1070),
.B1(n_1075),
.B2(n_1071),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1387),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1390),
.B(n_630),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1456),
.B(n_1130),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1387),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1471),
.B(n_630),
.Y(n_1659)
);

AOI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1416),
.A2(n_1288),
.B1(n_1285),
.B2(n_1246),
.Y(n_1660)
);

NOR3xp33_ASAP7_75t_L g1661 ( 
.A(n_1339),
.B(n_512),
.C(n_508),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1522),
.B(n_1227),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1456),
.B(n_1130),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1458),
.B(n_1161),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1388),
.Y(n_1665)
);

NAND2xp33_ASAP7_75t_L g1666 ( 
.A(n_1354),
.B(n_1185),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1388),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1399),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1414),
.B(n_513),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1409),
.B(n_631),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1522),
.B(n_1231),
.Y(n_1671)
);

BUFx8_ASAP7_75t_L g1672 ( 
.A(n_1457),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1399),
.Y(n_1673)
);

XOR2xp5_ASAP7_75t_L g1674 ( 
.A(n_1358),
.B(n_360),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1416),
.A2(n_1272),
.B1(n_1276),
.B2(n_1267),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1421),
.A2(n_1247),
.B1(n_1249),
.B2(n_1246),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1458),
.B(n_1161),
.Y(n_1677)
);

NOR3xp33_ASAP7_75t_L g1678 ( 
.A(n_1317),
.B(n_516),
.C(n_515),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1416),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1465),
.B(n_1161),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1522),
.B(n_1231),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1435),
.A2(n_1283),
.B1(n_1285),
.B2(n_1279),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1522),
.B(n_1233),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1414),
.B(n_518),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1465),
.B(n_1161),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1512),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1311),
.B(n_1233),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1494),
.B(n_1177),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1494),
.B(n_1177),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1298),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1431),
.B(n_1338),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1338),
.B(n_1238),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1407),
.Y(n_1693)
);

NOR2xp67_ASAP7_75t_SL g1694 ( 
.A(n_1316),
.B(n_600),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1407),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1500),
.B(n_1177),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1411),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1464),
.B(n_892),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1527),
.B(n_1238),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1411),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1500),
.B(n_1177),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1413),
.Y(n_1702)
);

NAND2xp33_ASAP7_75t_L g1703 ( 
.A(n_1354),
.B(n_1185),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1413),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1418),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1418),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1518),
.B(n_892),
.Y(n_1707)
);

AND2x4_ASAP7_75t_SL g1708 ( 
.A(n_1436),
.B(n_631),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1421),
.A2(n_1249),
.B1(n_1252),
.B2(n_1247),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1502),
.B(n_1255),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1419),
.Y(n_1711)
);

NOR2xp67_ASAP7_75t_L g1712 ( 
.A(n_1514),
.B(n_1240),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1419),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1425),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1425),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1375),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1430),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1502),
.B(n_1255),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1504),
.B(n_1363),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1451),
.B(n_631),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1335),
.B(n_520),
.Y(n_1721)
);

INVx2_ASAP7_75t_SL g1722 ( 
.A(n_1513),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1430),
.Y(n_1723)
);

OR2x6_ASAP7_75t_L g1724 ( 
.A(n_1370),
.B(n_1240),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1433),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1504),
.B(n_1255),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1433),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1452),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1452),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_SL g1730 ( 
.A1(n_1511),
.A2(n_1518),
.B1(n_1358),
.B2(n_1457),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1296),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1296),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1496),
.B(n_631),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1364),
.B(n_1256),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1319),
.Y(n_1735)
);

AND2x2_ASAP7_75t_SL g1736 ( 
.A(n_1362),
.B(n_603),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1319),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1435),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1505),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1459),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1391),
.B(n_1256),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_SL g1742 ( 
.A(n_1355),
.B(n_1251),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1436),
.B(n_1251),
.Y(n_1743)
);

NOR3xp33_ASAP7_75t_L g1744 ( 
.A(n_1337),
.B(n_525),
.C(n_523),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1435),
.A2(n_1288),
.B1(n_1252),
.B2(n_1254),
.Y(n_1745)
);

NAND2xp33_ASAP7_75t_L g1746 ( 
.A(n_1354),
.B(n_1185),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1448),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_L g1748 ( 
.A(n_1375),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1505),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1294),
.B(n_1324),
.Y(n_1750)
);

BUFx3_ASAP7_75t_L g1751 ( 
.A(n_1298),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1508),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1466),
.B(n_530),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1508),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1469),
.B(n_532),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1472),
.B(n_1256),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1511),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1481),
.B(n_536),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1485),
.B(n_1253),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1375),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1356),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1516),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1436),
.B(n_1266),
.Y(n_1763)
);

BUFx3_ASAP7_75t_L g1764 ( 
.A(n_1322),
.Y(n_1764)
);

INVx3_ASAP7_75t_L g1765 ( 
.A(n_1356),
.Y(n_1765)
);

INVx4_ASAP7_75t_L g1766 ( 
.A(n_1316),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1428),
.B(n_724),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1487),
.B(n_1253),
.Y(n_1768)
);

A2O1A1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1449),
.A2(n_613),
.B(n_627),
.C(n_611),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1490),
.B(n_1254),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1299),
.Y(n_1771)
);

BUFx6f_ASAP7_75t_SL g1772 ( 
.A(n_1392),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1445),
.B(n_1266),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1443),
.B(n_1483),
.Y(n_1774)
);

OR2x6_ASAP7_75t_L g1775 ( 
.A(n_1392),
.B(n_1275),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1445),
.Y(n_1776)
);

NOR2x1p5_ASAP7_75t_L g1777 ( 
.A(n_1427),
.B(n_540),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1443),
.B(n_1257),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1483),
.B(n_1257),
.Y(n_1779)
);

OAI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1474),
.A2(n_1075),
.B1(n_1081),
.B2(n_1079),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1459),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1470),
.A2(n_1204),
.B(n_1134),
.Y(n_1782)
);

BUFx2_ASAP7_75t_L g1783 ( 
.A(n_1607),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1545),
.B(n_1461),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1559),
.B(n_1421),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_R g1786 ( 
.A(n_1686),
.B(n_1437),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1731),
.Y(n_1787)
);

INVx4_ASAP7_75t_L g1788 ( 
.A(n_1584),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1538),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1766),
.A2(n_1362),
.B(n_1605),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1538),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1774),
.B(n_1533),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1541),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1560),
.Y(n_1794)
);

NAND2x1p5_ASAP7_75t_L g1795 ( 
.A(n_1766),
.B(n_1351),
.Y(n_1795)
);

O2A1O1Ixp5_ASAP7_75t_L g1796 ( 
.A1(n_1750),
.A2(n_1528),
.B(n_1447),
.C(n_1345),
.Y(n_1796)
);

BUFx2_ASAP7_75t_L g1797 ( 
.A(n_1543),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1550),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1550),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1669),
.B(n_1533),
.Y(n_1800)
);

OR2x6_ASAP7_75t_L g1801 ( 
.A(n_1757),
.B(n_1427),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1636),
.A2(n_1302),
.B1(n_1382),
.B2(n_1378),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1736),
.A2(n_1426),
.B1(n_1354),
.B2(n_1393),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1731),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1562),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1736),
.A2(n_1426),
.B1(n_1661),
.B2(n_1574),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1684),
.A2(n_1426),
.B1(n_1354),
.B2(n_1393),
.Y(n_1807)
);

AND2x6_ASAP7_75t_SL g1808 ( 
.A(n_1599),
.B(n_1299),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1541),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1738),
.A2(n_1302),
.B1(n_1467),
.B2(n_1325),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1562),
.Y(n_1811)
);

BUFx12f_ASAP7_75t_L g1812 ( 
.A(n_1672),
.Y(n_1812)
);

NOR2x2_ASAP7_75t_L g1813 ( 
.A(n_1724),
.B(n_1299),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1690),
.B(n_1322),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1565),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1546),
.B(n_1548),
.Y(n_1816)
);

INVx4_ASAP7_75t_L g1817 ( 
.A(n_1584),
.Y(n_1817)
);

BUFx2_ASAP7_75t_L g1818 ( 
.A(n_1690),
.Y(n_1818)
);

INVx2_ASAP7_75t_SL g1819 ( 
.A(n_1698),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1732),
.Y(n_1820)
);

BUFx4f_ASAP7_75t_L g1821 ( 
.A(n_1724),
.Y(n_1821)
);

BUFx3_ASAP7_75t_L g1822 ( 
.A(n_1751),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1732),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1686),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1565),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1587),
.B(n_1516),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1766),
.B(n_1445),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1580),
.Y(n_1828)
);

INVx2_ASAP7_75t_SL g1829 ( 
.A(n_1670),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1751),
.B(n_1325),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1735),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1719),
.B(n_1519),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1591),
.B(n_1519),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1539),
.B(n_1540),
.Y(n_1834)
);

BUFx6f_ASAP7_75t_L g1835 ( 
.A(n_1584),
.Y(n_1835)
);

BUFx6f_ASAP7_75t_L g1836 ( 
.A(n_1584),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1572),
.B(n_1509),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1552),
.B(n_1557),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1679),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1568),
.B(n_1534),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1580),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_1570),
.Y(n_1842)
);

NOR3xp33_ASAP7_75t_SL g1843 ( 
.A(n_1577),
.B(n_544),
.C(n_543),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1575),
.A2(n_1426),
.B1(n_1354),
.B2(n_1393),
.Y(n_1844)
);

INVx3_ASAP7_75t_L g1845 ( 
.A(n_1541),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1589),
.B(n_1356),
.Y(n_1846)
);

BUFx6f_ASAP7_75t_L g1847 ( 
.A(n_1716),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_R g1848 ( 
.A(n_1571),
.B(n_1406),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1707),
.B(n_1747),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1592),
.B(n_1534),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1624),
.A2(n_1367),
.B1(n_1393),
.B2(n_1326),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1589),
.B(n_1361),
.Y(n_1852)
);

OR2x6_ASAP7_75t_L g1853 ( 
.A(n_1738),
.B(n_1482),
.Y(n_1853)
);

BUFx12f_ASAP7_75t_L g1854 ( 
.A(n_1672),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1582),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1582),
.Y(n_1856)
);

AO22x1_ASAP7_75t_L g1857 ( 
.A1(n_1721),
.A2(n_1482),
.B1(n_1393),
.B2(n_1367),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1628),
.B(n_1367),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1735),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1633),
.B(n_1367),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1643),
.A2(n_1393),
.B1(n_1367),
.B2(n_1462),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_SL g1862 ( 
.A1(n_1730),
.A2(n_1674),
.B1(n_1771),
.B2(n_1299),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1586),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_L g1864 ( 
.A(n_1716),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1573),
.B(n_1367),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1573),
.B(n_1377),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1656),
.B(n_1523),
.Y(n_1867)
);

BUFx3_ASAP7_75t_L g1868 ( 
.A(n_1764),
.Y(n_1868)
);

INVx2_ASAP7_75t_SL g1869 ( 
.A(n_1659),
.Y(n_1869)
);

INVx2_ASAP7_75t_SL g1870 ( 
.A(n_1764),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1586),
.Y(n_1871)
);

AOI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1573),
.A2(n_1467),
.B1(n_1432),
.B2(n_1441),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1589),
.B(n_1509),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1678),
.A2(n_1653),
.B1(n_1733),
.B2(n_1720),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1570),
.Y(n_1875)
);

BUFx3_ASAP7_75t_L g1876 ( 
.A(n_1672),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1737),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1598),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1622),
.B(n_1385),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1776),
.B(n_1351),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_SL g1881 ( 
.A(n_1563),
.B(n_724),
.Y(n_1881)
);

NAND2xp33_ASAP7_75t_L g1882 ( 
.A(n_1589),
.B(n_1351),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1610),
.B(n_1462),
.Y(n_1883)
);

BUFx3_ASAP7_75t_L g1884 ( 
.A(n_1724),
.Y(n_1884)
);

BUFx2_ASAP7_75t_L g1885 ( 
.A(n_1724),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1640),
.A2(n_1316),
.B1(n_1480),
.B2(n_1509),
.Y(n_1886)
);

NAND2x1p5_ASAP7_75t_L g1887 ( 
.A(n_1625),
.B(n_1351),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1589),
.B(n_1361),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1589),
.B(n_1402),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1589),
.B(n_1361),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1598),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1776),
.B(n_1351),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1612),
.A2(n_1468),
.B1(n_1473),
.B2(n_1463),
.Y(n_1893)
);

AOI211xp5_ASAP7_75t_L g1894 ( 
.A1(n_1767),
.A2(n_627),
.B(n_637),
.C(n_613),
.Y(n_1894)
);

BUFx3_ASAP7_75t_L g1895 ( 
.A(n_1775),
.Y(n_1895)
);

NOR3xp33_ASAP7_75t_SL g1896 ( 
.A(n_1594),
.B(n_547),
.C(n_545),
.Y(n_1896)
);

NAND2x1p5_ASAP7_75t_L g1897 ( 
.A(n_1625),
.B(n_1318),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1570),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1716),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1602),
.B(n_1463),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1612),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1613),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1613),
.Y(n_1903)
);

INVxp67_ASAP7_75t_L g1904 ( 
.A(n_1606),
.Y(n_1904)
);

A2O1A1Ixp33_ASAP7_75t_L g1905 ( 
.A1(n_1594),
.A2(n_1615),
.B(n_1749),
.C(n_1739),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_1601),
.B(n_1383),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1617),
.Y(n_1907)
);

AOI211xp5_ASAP7_75t_L g1908 ( 
.A1(n_1744),
.A2(n_641),
.B(n_644),
.C(n_637),
.Y(n_1908)
);

BUFx4f_ASAP7_75t_L g1909 ( 
.A(n_1775),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1601),
.B(n_1383),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1617),
.Y(n_1911)
);

A2O1A1Ixp33_ASAP7_75t_L g1912 ( 
.A1(n_1752),
.A2(n_1524),
.B(n_1520),
.C(n_1303),
.Y(n_1912)
);

OR2x6_ASAP7_75t_L g1913 ( 
.A(n_1611),
.B(n_1316),
.Y(n_1913)
);

HB1xp67_ASAP7_75t_L g1914 ( 
.A(n_1716),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1754),
.B(n_1404),
.Y(n_1915)
);

BUFx12f_ASAP7_75t_L g1916 ( 
.A(n_1771),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1753),
.B(n_724),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1755),
.B(n_1758),
.Y(n_1918)
);

BUFx4f_ASAP7_75t_L g1919 ( 
.A(n_1775),
.Y(n_1919)
);

HB1xp67_ASAP7_75t_L g1920 ( 
.A(n_1748),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1619),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1737),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1762),
.B(n_1405),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1619),
.Y(n_1924)
);

AND2x6_ASAP7_75t_L g1925 ( 
.A(n_1601),
.B(n_1614),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1535),
.B(n_1417),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1630),
.B(n_1468),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1630),
.B(n_1473),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_1772),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1644),
.B(n_1475),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1775),
.B(n_1475),
.Y(n_1931)
);

INVx5_ASAP7_75t_L g1932 ( 
.A(n_1748),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1644),
.B(n_1658),
.Y(n_1933)
);

BUFx6f_ASAP7_75t_L g1934 ( 
.A(n_1748),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1658),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1668),
.B(n_1478),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1668),
.B(n_1478),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1693),
.B(n_1486),
.Y(n_1938)
);

AOI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1544),
.A2(n_1495),
.B1(n_1498),
.B2(n_1455),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1693),
.Y(n_1940)
);

AOI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1544),
.A2(n_1486),
.B1(n_1531),
.B2(n_1530),
.Y(n_1941)
);

INVx3_ASAP7_75t_L g1942 ( 
.A(n_1748),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1702),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1702),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1705),
.Y(n_1945)
);

OR2x6_ASAP7_75t_L g1946 ( 
.A(n_1611),
.B(n_1524),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1705),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1706),
.B(n_1530),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1706),
.Y(n_1949)
);

AND2x6_ASAP7_75t_SL g1950 ( 
.A(n_1556),
.B(n_641),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1713),
.Y(n_1951)
);

OAI22xp5_ASAP7_75t_SL g1952 ( 
.A1(n_1722),
.A2(n_566),
.B1(n_584),
.B2(n_552),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1713),
.B(n_1531),
.Y(n_1953)
);

AND2x2_ASAP7_75t_SL g1954 ( 
.A(n_1666),
.B(n_1381),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_1772),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1717),
.Y(n_1956)
);

INVxp67_ASAP7_75t_SL g1957 ( 
.A(n_1760),
.Y(n_1957)
);

AOI21xp33_ASAP7_75t_L g1958 ( 
.A1(n_1722),
.A2(n_1520),
.B(n_1493),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1717),
.B(n_1493),
.Y(n_1959)
);

NAND2x1p5_ASAP7_75t_L g1960 ( 
.A(n_1623),
.B(n_1503),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1614),
.B(n_1383),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1727),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1727),
.Y(n_1963)
);

INVx3_ASAP7_75t_L g1964 ( 
.A(n_1760),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1614),
.B(n_1761),
.Y(n_1965)
);

BUFx6f_ASAP7_75t_L g1966 ( 
.A(n_1760),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1761),
.B(n_1408),
.Y(n_1967)
);

OR2x6_ASAP7_75t_L g1968 ( 
.A(n_1611),
.B(n_1777),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1650),
.Y(n_1969)
);

O2A1O1Ixp5_ASAP7_75t_L g1970 ( 
.A1(n_1694),
.A2(n_1507),
.B(n_1506),
.C(n_1453),
.Y(n_1970)
);

AOI211xp5_ASAP7_75t_L g1971 ( 
.A1(n_1769),
.A2(n_648),
.B(n_649),
.C(n_644),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1651),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1632),
.B(n_1521),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1655),
.Y(n_1974)
);

BUFx3_ASAP7_75t_L g1975 ( 
.A(n_1760),
.Y(n_1975)
);

NOR2x1_ASAP7_75t_R g1976 ( 
.A(n_1772),
.B(n_548),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1665),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1558),
.Y(n_1978)
);

OR2x6_ASAP7_75t_L g1979 ( 
.A(n_1611),
.B(n_1297),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1740),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_L g1981 ( 
.A(n_1667),
.B(n_1408),
.Y(n_1981)
);

AOI22xp33_ASAP7_75t_SL g1982 ( 
.A1(n_1558),
.A2(n_749),
.B1(n_777),
.B2(n_724),
.Y(n_1982)
);

OR2x6_ASAP7_75t_L g1983 ( 
.A(n_1590),
.B(n_1303),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1708),
.B(n_1521),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1761),
.B(n_1408),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1673),
.B(n_1442),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1740),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1695),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1781),
.Y(n_1989)
);

INVx5_ASAP7_75t_L g1990 ( 
.A(n_1623),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1708),
.B(n_749),
.Y(n_1991)
);

AO22x1_ASAP7_75t_L g1992 ( 
.A1(n_1623),
.A2(n_550),
.B1(n_553),
.B2(n_549),
.Y(n_1992)
);

INVx3_ASAP7_75t_L g1993 ( 
.A(n_1765),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1697),
.B(n_1700),
.Y(n_1994)
);

OAI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1547),
.A2(n_1489),
.B1(n_1477),
.B2(n_1442),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1704),
.B(n_1442),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1781),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1711),
.B(n_1477),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1918),
.B(n_1648),
.Y(n_1999)
);

NAND2xp33_ASAP7_75t_SL g2000 ( 
.A(n_1786),
.B(n_1648),
.Y(n_2000)
);

NAND2xp33_ASAP7_75t_SL g2001 ( 
.A(n_1786),
.B(n_1648),
.Y(n_2001)
);

NAND2xp33_ASAP7_75t_SL g2002 ( 
.A(n_1848),
.B(n_1590),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1816),
.B(n_1714),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_SL g2004 ( 
.A(n_1918),
.B(n_1600),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1829),
.B(n_1715),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1784),
.B(n_1883),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1800),
.B(n_1723),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_SL g2008 ( 
.A(n_1883),
.B(n_1725),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1826),
.B(n_1536),
.Y(n_2009)
);

NAND2xp33_ASAP7_75t_SL g2010 ( 
.A(n_1848),
.B(n_1649),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1849),
.B(n_1728),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1849),
.B(n_1729),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_SL g2013 ( 
.A(n_1802),
.B(n_1765),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1867),
.B(n_1833),
.Y(n_2014)
);

AND2x4_ASAP7_75t_L g2015 ( 
.A(n_1884),
.B(n_1645),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1869),
.B(n_1765),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1867),
.B(n_1537),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1819),
.B(n_1645),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_1874),
.B(n_1645),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1794),
.B(n_1712),
.Y(n_2020)
);

NAND2xp33_ASAP7_75t_SL g2021 ( 
.A(n_1824),
.B(n_1978),
.Y(n_2021)
);

NAND2xp33_ASAP7_75t_SL g2022 ( 
.A(n_1896),
.B(n_1676),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1794),
.B(n_1691),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1783),
.B(n_1691),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_1881),
.B(n_1709),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1904),
.B(n_1660),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_SL g2027 ( 
.A(n_1814),
.B(n_1675),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_1814),
.B(n_1682),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1830),
.B(n_1745),
.Y(n_2029)
);

NAND2xp33_ASAP7_75t_SL g2030 ( 
.A(n_1896),
.B(n_1616),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1830),
.B(n_1542),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1806),
.B(n_1769),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_1797),
.B(n_1778),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1917),
.B(n_1779),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_SL g2035 ( 
.A(n_1810),
.B(n_1554),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1982),
.B(n_1564),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1818),
.B(n_1822),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1900),
.B(n_1549),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1806),
.B(n_1583),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1900),
.B(n_1595),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1798),
.B(n_1652),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1822),
.B(n_1868),
.Y(n_2042)
);

NAND2xp33_ASAP7_75t_SL g2043 ( 
.A(n_1843),
.B(n_1616),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1868),
.B(n_1567),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1832),
.B(n_1759),
.Y(n_2045)
);

NAND2xp33_ASAP7_75t_SL g2046 ( 
.A(n_1843),
.B(n_1627),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1785),
.B(n_1569),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1894),
.B(n_1991),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1792),
.B(n_1879),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_1870),
.B(n_1768),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_SL g2051 ( 
.A(n_1839),
.B(n_1770),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_SL g2052 ( 
.A(n_1839),
.B(n_1579),
.Y(n_2052)
);

AND2x2_ASAP7_75t_SL g2053 ( 
.A(n_1954),
.B(n_1666),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1908),
.B(n_1603),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1984),
.B(n_1551),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1901),
.B(n_1903),
.Y(n_2056)
);

NAND2xp33_ASAP7_75t_SL g2057 ( 
.A(n_1842),
.B(n_1627),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_SL g2058 ( 
.A(n_1931),
.B(n_1551),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1931),
.B(n_1834),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1838),
.B(n_1734),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_SL g2061 ( 
.A(n_1821),
.B(n_1741),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_1821),
.B(n_1756),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_1909),
.B(n_1710),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1909),
.B(n_1718),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1915),
.B(n_1652),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_SL g2066 ( 
.A(n_1919),
.B(n_1807),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_SL g2067 ( 
.A(n_1919),
.B(n_1726),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1807),
.B(n_1561),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1990),
.B(n_1561),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1923),
.B(n_1926),
.Y(n_2070)
);

NAND2xp33_ASAP7_75t_SL g2071 ( 
.A(n_1875),
.B(n_1629),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_SL g2072 ( 
.A(n_1990),
.B(n_1566),
.Y(n_2072)
);

NAND2xp33_ASAP7_75t_SL g2073 ( 
.A(n_1898),
.B(n_1629),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_1990),
.B(n_1566),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1866),
.B(n_1585),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_SL g2076 ( 
.A(n_1990),
.B(n_1803),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1803),
.B(n_1692),
.Y(n_2077)
);

NAND2xp33_ASAP7_75t_SL g2078 ( 
.A(n_1929),
.B(n_1637),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_SL g2079 ( 
.A(n_1955),
.B(n_1692),
.Y(n_2079)
);

NAND2xp33_ASAP7_75t_SL g2080 ( 
.A(n_1862),
.B(n_1637),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_SL g2081 ( 
.A(n_1952),
.B(n_1844),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1844),
.B(n_1743),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1924),
.B(n_1588),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_SL g2084 ( 
.A(n_1932),
.B(n_1743),
.Y(n_2084)
);

NAND2xp33_ASAP7_75t_SL g2085 ( 
.A(n_1885),
.B(n_1639),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_SL g2086 ( 
.A(n_1932),
.B(n_1865),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_SL g2087 ( 
.A(n_1932),
.B(n_1763),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_SL g2088 ( 
.A(n_1932),
.B(n_1763),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_1880),
.B(n_1773),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_SL g2090 ( 
.A(n_1880),
.B(n_1773),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_SL g2091 ( 
.A(n_1892),
.B(n_1581),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_SL g2092 ( 
.A(n_1892),
.B(n_1593),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_1796),
.B(n_1596),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1840),
.B(n_1742),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_SL g2095 ( 
.A(n_1969),
.B(n_1596),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_SL g2096 ( 
.A(n_1972),
.B(n_1604),
.Y(n_2096)
);

NAND2xp33_ASAP7_75t_SL g2097 ( 
.A(n_1835),
.B(n_1639),
.Y(n_2097)
);

NAND2xp33_ASAP7_75t_SL g2098 ( 
.A(n_1835),
.B(n_1641),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_SL g2099 ( 
.A(n_1974),
.B(n_1604),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1850),
.B(n_1742),
.Y(n_2100)
);

AND2x2_ASAP7_75t_SL g2101 ( 
.A(n_1954),
.B(n_1703),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_1977),
.B(n_1396),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_SL g2103 ( 
.A(n_1988),
.B(n_1396),
.Y(n_2103)
);

NAND2xp33_ASAP7_75t_SL g2104 ( 
.A(n_1835),
.B(n_1836),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_SL g2105 ( 
.A(n_1973),
.B(n_1396),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_SL g2106 ( 
.A(n_1973),
.B(n_1396),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_SL g2107 ( 
.A(n_1876),
.B(n_1396),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_1876),
.B(n_1429),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1905),
.B(n_1609),
.Y(n_2109)
);

NAND2xp33_ASAP7_75t_SL g2110 ( 
.A(n_1835),
.B(n_1641),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_1993),
.B(n_1429),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1905),
.B(n_1620),
.Y(n_2112)
);

NAND2xp33_ASAP7_75t_SL g2113 ( 
.A(n_1836),
.B(n_1662),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_1993),
.B(n_1429),
.Y(n_2114)
);

NAND2xp33_ASAP7_75t_SL g2115 ( 
.A(n_1836),
.B(n_1662),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_SL g2116 ( 
.A(n_1884),
.B(n_1429),
.Y(n_2116)
);

OR2x2_ASAP7_75t_L g2117 ( 
.A(n_1994),
.B(n_1680),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1943),
.B(n_1321),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_SL g2119 ( 
.A(n_1895),
.B(n_1429),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1895),
.B(n_1484),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_1947),
.B(n_1321),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_1793),
.B(n_1484),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1787),
.B(n_1621),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_1793),
.B(n_1484),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_1809),
.B(n_1484),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_SL g2126 ( 
.A(n_1809),
.B(n_1845),
.Y(n_2126)
);

NAND2x1_ASAP7_75t_L g2127 ( 
.A(n_1913),
.B(n_1318),
.Y(n_2127)
);

NAND2xp33_ASAP7_75t_SL g2128 ( 
.A(n_1836),
.B(n_1671),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_1845),
.B(n_1858),
.Y(n_2129)
);

NAND2xp33_ASAP7_75t_SL g2130 ( 
.A(n_1847),
.B(n_1864),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_1949),
.B(n_1980),
.Y(n_2131)
);

NAND2xp33_ASAP7_75t_SL g2132 ( 
.A(n_1847),
.B(n_1671),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_SL g2133 ( 
.A(n_1860),
.B(n_1851),
.Y(n_2133)
);

AND2x4_ASAP7_75t_L g2134 ( 
.A(n_1968),
.B(n_1681),
.Y(n_2134)
);

AND2x4_ASAP7_75t_L g2135 ( 
.A(n_1968),
.B(n_1681),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_1851),
.B(n_1484),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1787),
.B(n_1327),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_SL g2138 ( 
.A(n_1847),
.B(n_1497),
.Y(n_2138)
);

NAND2xp33_ASAP7_75t_SL g2139 ( 
.A(n_1847),
.B(n_1683),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_SL g2140 ( 
.A(n_1864),
.B(n_1497),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_SL g2141 ( 
.A(n_1864),
.B(n_1497),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_SL g2142 ( 
.A(n_1864),
.B(n_1934),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_SL g2143 ( 
.A(n_1934),
.B(n_1497),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_SL g2144 ( 
.A(n_1934),
.B(n_1497),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_SL g2145 ( 
.A(n_1934),
.B(n_1499),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_SL g2146 ( 
.A(n_1966),
.B(n_1916),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_SL g2147 ( 
.A(n_1966),
.B(n_1499),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_SL g2148 ( 
.A(n_1966),
.B(n_1499),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_SL g2149 ( 
.A(n_1966),
.B(n_1499),
.Y(n_2149)
);

NAND2xp33_ASAP7_75t_SL g2150 ( 
.A(n_1788),
.B(n_1817),
.Y(n_2150)
);

AND2x4_ASAP7_75t_L g2151 ( 
.A(n_1968),
.B(n_1683),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1804),
.B(n_1327),
.Y(n_2152)
);

NAND2xp33_ASAP7_75t_SL g2153 ( 
.A(n_1788),
.B(n_1626),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_SL g2154 ( 
.A(n_1872),
.B(n_1499),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1804),
.B(n_1336),
.Y(n_2155)
);

NAND2xp33_ASAP7_75t_SL g2156 ( 
.A(n_1817),
.B(n_1631),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_SL g2157 ( 
.A(n_1889),
.B(n_1634),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_SL g2158 ( 
.A(n_1861),
.B(n_1893),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_SL g2159 ( 
.A(n_1861),
.B(n_1635),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1820),
.B(n_1336),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1820),
.B(n_1340),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_SL g2162 ( 
.A(n_1893),
.B(n_1663),
.Y(n_2162)
);

NAND2xp33_ASAP7_75t_SL g2163 ( 
.A(n_1914),
.B(n_1638),
.Y(n_2163)
);

NAND2xp33_ASAP7_75t_SL g2164 ( 
.A(n_1914),
.B(n_1642),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1823),
.B(n_1340),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_SL g2166 ( 
.A(n_1975),
.B(n_1688),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_SL g2167 ( 
.A(n_1975),
.B(n_1689),
.Y(n_2167)
);

NAND2xp33_ASAP7_75t_SL g2168 ( 
.A(n_1920),
.B(n_1647),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_1812),
.B(n_1696),
.Y(n_2169)
);

NAND2xp33_ASAP7_75t_SL g2170 ( 
.A(n_1920),
.B(n_1657),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1823),
.B(n_1618),
.Y(n_2171)
);

NAND2xp33_ASAP7_75t_SL g2172 ( 
.A(n_1837),
.B(n_1664),
.Y(n_2172)
);

AND2x4_ASAP7_75t_L g2173 ( 
.A(n_1913),
.B(n_1553),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_SL g2174 ( 
.A(n_1854),
.B(n_1677),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_SL g2175 ( 
.A(n_1886),
.B(n_1685),
.Y(n_2175)
);

NAND2xp33_ASAP7_75t_SL g2176 ( 
.A(n_1837),
.B(n_1701),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_1940),
.B(n_1687),
.Y(n_2177)
);

NAND2xp33_ASAP7_75t_SL g2178 ( 
.A(n_1827),
.B(n_1553),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_1940),
.B(n_1477),
.Y(n_2179)
);

NAND2xp33_ASAP7_75t_SL g2180 ( 
.A(n_1827),
.B(n_1555),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_1944),
.B(n_1489),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1831),
.B(n_1555),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_1944),
.B(n_1489),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1831),
.B(n_1576),
.Y(n_2184)
);

NAND2xp33_ASAP7_75t_SL g2185 ( 
.A(n_1899),
.B(n_1576),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1962),
.B(n_1608),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_SL g2187 ( 
.A(n_1962),
.B(n_1318),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_1963),
.B(n_1360),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_SL g2189 ( 
.A(n_1963),
.B(n_1360),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_SL g2190 ( 
.A(n_1987),
.B(n_1989),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_SL g2191 ( 
.A(n_1987),
.B(n_1360),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_SL g2192 ( 
.A(n_1989),
.B(n_1438),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1859),
.B(n_1687),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1859),
.B(n_1877),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_1997),
.B(n_1438),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_SL g2196 ( 
.A(n_1997),
.B(n_1438),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_SL g2197 ( 
.A(n_1789),
.B(n_1450),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_SL g2198 ( 
.A(n_1791),
.B(n_1799),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_SL g2199 ( 
.A(n_1805),
.B(n_1811),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_SL g2200 ( 
.A(n_1815),
.B(n_1450),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_1825),
.B(n_1450),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_SL g2202 ( 
.A(n_1828),
.B(n_1476),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_1841),
.B(n_1476),
.Y(n_2203)
);

NAND2xp33_ASAP7_75t_SL g2204 ( 
.A(n_1899),
.B(n_1476),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_SL g2205 ( 
.A(n_1855),
.B(n_1479),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_SL g2206 ( 
.A(n_1856),
.B(n_1479),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_SL g2207 ( 
.A(n_1863),
.B(n_1479),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_1871),
.B(n_1503),
.Y(n_2208)
);

NAND2xp33_ASAP7_75t_SL g2209 ( 
.A(n_1942),
.B(n_1503),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_SL g2210 ( 
.A(n_1878),
.B(n_1517),
.Y(n_2210)
);

NAND2xp33_ASAP7_75t_SL g2211 ( 
.A(n_1942),
.B(n_1517),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1877),
.B(n_1699),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_SL g2213 ( 
.A(n_1891),
.B(n_1517),
.Y(n_2213)
);

NAND2xp33_ASAP7_75t_SL g2214 ( 
.A(n_1964),
.B(n_1525),
.Y(n_2214)
);

NAND2xp33_ASAP7_75t_R g2215 ( 
.A(n_1801),
.B(n_1444),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_1902),
.B(n_1699),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1922),
.B(n_1510),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_1907),
.B(n_1525),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_SL g2219 ( 
.A(n_1911),
.B(n_1525),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_SL g2220 ( 
.A(n_1921),
.B(n_1422),
.Y(n_2220)
);

NAND2xp33_ASAP7_75t_SL g2221 ( 
.A(n_1964),
.B(n_1703),
.Y(n_2221)
);

AND2x4_ASAP7_75t_L g2222 ( 
.A(n_1913),
.B(n_1782),
.Y(n_2222)
);

AND2x4_ASAP7_75t_L g2223 ( 
.A(n_1979),
.B(n_1532),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_SL g2224 ( 
.A(n_1935),
.B(n_1945),
.Y(n_2224)
);

NAND2xp33_ASAP7_75t_SL g2225 ( 
.A(n_1951),
.B(n_1746),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_1956),
.B(n_1422),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1922),
.B(n_1780),
.Y(n_2227)
);

NAND2xp33_ASAP7_75t_SL g2228 ( 
.A(n_1846),
.B(n_1746),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1933),
.B(n_1578),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_SL g2230 ( 
.A(n_1981),
.B(n_1422),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_SL g2231 ( 
.A(n_1981),
.B(n_1597),
.Y(n_2231)
);

NAND2xp33_ASAP7_75t_SL g2232 ( 
.A(n_1846),
.B(n_1654),
.Y(n_2232)
);

NAND2xp33_ASAP7_75t_SL g2233 ( 
.A(n_1852),
.B(n_1454),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_SL g2234 ( 
.A(n_1941),
.B(n_1488),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2003),
.B(n_1801),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2056),
.Y(n_2236)
);

OAI21x1_ASAP7_75t_L g2237 ( 
.A1(n_2093),
.A2(n_1790),
.B(n_1646),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_2021),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_2002),
.Y(n_2239)
);

CKINVDCx5p33_ASAP7_75t_R g2240 ( 
.A(n_2146),
.Y(n_2240)
);

OR2x2_ASAP7_75t_L g2241 ( 
.A(n_2014),
.B(n_1801),
.Y(n_2241)
);

INVx4_ASAP7_75t_L g2242 ( 
.A(n_2015),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_2003),
.B(n_1992),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2006),
.B(n_1971),
.Y(n_2244)
);

NOR2xp33_ASAP7_75t_R g2245 ( 
.A(n_2000),
.B(n_1808),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2070),
.B(n_1950),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2056),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2118),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_2042),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_2118),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2131),
.Y(n_2251)
);

INVxp67_ASAP7_75t_L g2252 ( 
.A(n_2037),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2131),
.Y(n_2253)
);

CKINVDCx16_ASAP7_75t_R g2254 ( 
.A(n_2215),
.Y(n_2254)
);

INVx3_ASAP7_75t_L g2255 ( 
.A(n_2015),
.Y(n_2255)
);

AO21x1_ASAP7_75t_L g2256 ( 
.A1(n_2004),
.A2(n_1882),
.B(n_1578),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2194),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2194),
.Y(n_2258)
);

INVx1_ASAP7_75t_SL g2259 ( 
.A(n_2001),
.Y(n_2259)
);

AOI22xp33_ASAP7_75t_SL g2260 ( 
.A1(n_2053),
.A2(n_1853),
.B1(n_777),
.B2(n_749),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2049),
.B(n_1853),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2121),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2121),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2177),
.Y(n_2264)
);

AOI22xp33_ASAP7_75t_L g2265 ( 
.A1(n_2081),
.A2(n_777),
.B1(n_749),
.B2(n_649),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2177),
.Y(n_2266)
);

CKINVDCx5p33_ASAP7_75t_R g2267 ( 
.A(n_2010),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2137),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2017),
.B(n_1853),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2009),
.B(n_1927),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_2137),
.Y(n_2271)
);

BUFx2_ASAP7_75t_L g2272 ( 
.A(n_2015),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2184),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2040),
.B(n_1928),
.Y(n_2274)
);

BUFx4f_ASAP7_75t_L g2275 ( 
.A(n_2134),
.Y(n_2275)
);

INVx1_ASAP7_75t_SL g2276 ( 
.A(n_2020),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2034),
.B(n_2033),
.Y(n_2277)
);

AOI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_2048),
.A2(n_1857),
.B1(n_1983),
.B2(n_1939),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2045),
.B(n_1930),
.Y(n_2279)
);

NOR2xp33_ASAP7_75t_L g2280 ( 
.A(n_2054),
.B(n_1983),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2184),
.Y(n_2281)
);

OAI22xp5_ASAP7_75t_SL g2282 ( 
.A1(n_2053),
.A2(n_555),
.B1(n_557),
.B2(n_554),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2015),
.B(n_893),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2152),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2038),
.B(n_1936),
.Y(n_2285)
);

BUFx4f_ASAP7_75t_L g2286 ( 
.A(n_2134),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_2080),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2041),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_2057),
.Y(n_2289)
);

NOR2xp33_ASAP7_75t_R g2290 ( 
.A(n_2071),
.B(n_1925),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2152),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2041),
.Y(n_2292)
);

HB1xp67_ASAP7_75t_L g2293 ( 
.A(n_2018),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2182),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1999),
.B(n_2007),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2212),
.Y(n_2296)
);

AND2x4_ASAP7_75t_L g2297 ( 
.A(n_2134),
.B(n_1979),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2059),
.B(n_1937),
.Y(n_2298)
);

NOR2xp67_ASAP7_75t_L g2299 ( 
.A(n_2169),
.B(n_1965),
.Y(n_2299)
);

NAND2xp33_ASAP7_75t_L g2300 ( 
.A(n_2228),
.B(n_1925),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2051),
.B(n_893),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_2155),
.Y(n_2302)
);

INVxp67_ASAP7_75t_L g2303 ( 
.A(n_2011),
.Y(n_2303)
);

OAI22xp5_ASAP7_75t_L g2304 ( 
.A1(n_2053),
.A2(n_1983),
.B1(n_1979),
.B2(n_1946),
.Y(n_2304)
);

AOI22xp33_ASAP7_75t_L g2305 ( 
.A1(n_2032),
.A2(n_777),
.B1(n_650),
.B2(n_652),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_2023),
.B(n_894),
.Y(n_2306)
);

AND2x2_ASAP7_75t_SL g2307 ( 
.A(n_2101),
.B(n_1813),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2012),
.B(n_1938),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2024),
.B(n_894),
.Y(n_2309)
);

INVxp67_ASAP7_75t_SL g2310 ( 
.A(n_2171),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2031),
.B(n_1957),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2008),
.B(n_1957),
.Y(n_2312)
);

AOI22xp33_ASAP7_75t_SL g2313 ( 
.A1(n_2101),
.A2(n_1925),
.B1(n_650),
.B2(n_652),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2032),
.B(n_899),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_2026),
.B(n_2079),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2065),
.B(n_1948),
.Y(n_2316)
);

AOI22xp33_ASAP7_75t_L g2317 ( 
.A1(n_2025),
.A2(n_660),
.B1(n_664),
.B2(n_648),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2212),
.Y(n_2318)
);

AND3x1_ASAP7_75t_SL g2319 ( 
.A(n_2022),
.B(n_664),
.C(n_660),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_2101),
.B(n_1958),
.Y(n_2320)
);

A2O1A1Ixp33_ASAP7_75t_L g2321 ( 
.A1(n_2158),
.A2(n_2136),
.B(n_2077),
.C(n_2066),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2075),
.B(n_2083),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2083),
.B(n_2039),
.Y(n_2323)
);

A2O1A1Ixp33_ASAP7_75t_L g2324 ( 
.A1(n_2076),
.A2(n_1912),
.B(n_1995),
.C(n_1970),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2039),
.B(n_1953),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2216),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2216),
.Y(n_2327)
);

BUFx4f_ASAP7_75t_L g2328 ( 
.A(n_2134),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_L g2329 ( 
.A(n_2019),
.B(n_1965),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2117),
.B(n_2050),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2117),
.B(n_1976),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2036),
.B(n_1959),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2052),
.B(n_1986),
.Y(n_2333)
);

CKINVDCx5p33_ASAP7_75t_R g2334 ( 
.A(n_2073),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2198),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2094),
.B(n_1996),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2005),
.B(n_899),
.Y(n_2337)
);

CKINVDCx5p33_ASAP7_75t_R g2338 ( 
.A(n_2078),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2155),
.Y(n_2339)
);

CKINVDCx5p33_ASAP7_75t_R g2340 ( 
.A(n_2174),
.Y(n_2340)
);

OAI22xp5_ASAP7_75t_SL g2341 ( 
.A1(n_2135),
.A2(n_561),
.B1(n_565),
.B2(n_560),
.Y(n_2341)
);

BUFx8_ASAP7_75t_L g2342 ( 
.A(n_2135),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2199),
.Y(n_2343)
);

OAI22xp5_ASAP7_75t_L g2344 ( 
.A1(n_2027),
.A2(n_1946),
.B1(n_1795),
.B2(n_1960),
.Y(n_2344)
);

CKINVDCx20_ASAP7_75t_R g2345 ( 
.A(n_2043),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2224),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2100),
.B(n_2028),
.Y(n_2347)
);

OAI21x1_ASAP7_75t_L g2348 ( 
.A1(n_2154),
.A2(n_1873),
.B(n_1852),
.Y(n_2348)
);

BUFx8_ASAP7_75t_L g2349 ( 
.A(n_2135),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2193),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_2109),
.B(n_1960),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2029),
.B(n_1998),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2016),
.B(n_2044),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2160),
.Y(n_2354)
);

AOI22xp33_ASAP7_75t_SL g2355 ( 
.A1(n_2173),
.A2(n_1925),
.B1(n_667),
.B2(n_672),
.Y(n_2355)
);

BUFx8_ASAP7_75t_L g2356 ( 
.A(n_2135),
.Y(n_2356)
);

OAI22xp5_ASAP7_75t_L g2357 ( 
.A1(n_2091),
.A2(n_2068),
.B1(n_2058),
.B2(n_2112),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2160),
.Y(n_2358)
);

NOR3xp33_ASAP7_75t_L g2359 ( 
.A(n_2046),
.B(n_2030),
.C(n_2061),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2161),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2151),
.B(n_2107),
.Y(n_2361)
);

INVx6_ASAP7_75t_L g2362 ( 
.A(n_2151),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2161),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_2013),
.B(n_1873),
.Y(n_2364)
);

OAI22xp5_ASAP7_75t_SL g2365 ( 
.A1(n_2151),
.A2(n_569),
.B1(n_572),
.B2(n_568),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2060),
.B(n_574),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2165),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2151),
.B(n_900),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2035),
.B(n_575),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_2063),
.B(n_1888),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2055),
.B(n_578),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2165),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2064),
.B(n_583),
.Y(n_2373)
);

A2O1A1Ixp33_ASAP7_75t_L g2374 ( 
.A1(n_2082),
.A2(n_1912),
.B(n_1890),
.C(n_1888),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_2108),
.Y(n_2375)
);

AOI22xp33_ASAP7_75t_L g2376 ( 
.A1(n_2231),
.A2(n_667),
.B1(n_672),
.B2(n_666),
.Y(n_2376)
);

CKINVDCx20_ASAP7_75t_R g2377 ( 
.A(n_2150),
.Y(n_2377)
);

AOI22xp5_ASAP7_75t_L g2378 ( 
.A1(n_2085),
.A2(n_1925),
.B1(n_589),
.B2(n_590),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_2173),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2089),
.B(n_900),
.Y(n_2380)
);

AND3x1_ASAP7_75t_SL g2381 ( 
.A(n_2163),
.B(n_673),
.C(n_666),
.Y(n_2381)
);

NOR2xp33_ASAP7_75t_L g2382 ( 
.A(n_2133),
.B(n_1967),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2067),
.B(n_586),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2190),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2171),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2227),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_2090),
.B(n_901),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2227),
.Y(n_2388)
);

AOI22xp33_ASAP7_75t_L g2389 ( 
.A1(n_2172),
.A2(n_2176),
.B1(n_674),
.B2(n_677),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2062),
.B(n_595),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2092),
.B(n_2095),
.Y(n_2391)
);

AOI22xp33_ASAP7_75t_L g2392 ( 
.A1(n_2186),
.A2(n_674),
.B1(n_677),
.B2(n_673),
.Y(n_2392)
);

INVx6_ASAP7_75t_L g2393 ( 
.A(n_2173),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2123),
.Y(n_2394)
);

AND2x2_ASAP7_75t_SL g2395 ( 
.A(n_2222),
.B(n_1381),
.Y(n_2395)
);

AOI22x1_ASAP7_75t_L g2396 ( 
.A1(n_2173),
.A2(n_1887),
.B1(n_1897),
.B2(n_1795),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2217),
.Y(n_2397)
);

AO22x1_ASAP7_75t_L g2398 ( 
.A1(n_2223),
.A2(n_598),
.B1(n_599),
.B2(n_596),
.Y(n_2398)
);

INVx3_ASAP7_75t_L g2399 ( 
.A(n_2127),
.Y(n_2399)
);

OAI221xp5_ASAP7_75t_L g2400 ( 
.A1(n_2178),
.A2(n_902),
.B1(n_910),
.B2(n_907),
.C(n_901),
.Y(n_2400)
);

INVx3_ASAP7_75t_L g2401 ( 
.A(n_2127),
.Y(n_2401)
);

CKINVDCx20_ASAP7_75t_R g2402 ( 
.A(n_2104),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2116),
.B(n_902),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2096),
.B(n_602),
.Y(n_2404)
);

BUFx3_ASAP7_75t_L g2405 ( 
.A(n_2223),
.Y(n_2405)
);

AOI22xp5_ASAP7_75t_L g2406 ( 
.A1(n_2180),
.A2(n_2164),
.B1(n_2170),
.B2(n_2168),
.Y(n_2406)
);

INVx2_ASAP7_75t_SL g2407 ( 
.A(n_2142),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2119),
.B(n_2120),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2099),
.B(n_606),
.Y(n_2409)
);

NAND2xp33_ASAP7_75t_L g2410 ( 
.A(n_2225),
.B(n_1897),
.Y(n_2410)
);

BUFx3_ASAP7_75t_L g2411 ( 
.A(n_2223),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2179),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2181),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2223),
.B(n_907),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2183),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2086),
.B(n_910),
.Y(n_2416)
);

AOI22xp5_ASAP7_75t_L g2417 ( 
.A1(n_2222),
.A2(n_616),
.B1(n_618),
.B2(n_608),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2102),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2103),
.Y(n_2419)
);

OAI22xp5_ASAP7_75t_L g2420 ( 
.A1(n_2230),
.A2(n_1946),
.B1(n_1887),
.B2(n_1890),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2157),
.B(n_2229),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2166),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2167),
.Y(n_2423)
);

CKINVDCx20_ASAP7_75t_R g2424 ( 
.A(n_2130),
.Y(n_2424)
);

CKINVDCx11_ASAP7_75t_R g2425 ( 
.A(n_2222),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2105),
.B(n_619),
.Y(n_2426)
);

NAND2xp33_ASAP7_75t_L g2427 ( 
.A(n_2221),
.B(n_1906),
.Y(n_2427)
);

INVx3_ASAP7_75t_L g2428 ( 
.A(n_2222),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2111),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2106),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2114),
.Y(n_2431)
);

OR2x2_ASAP7_75t_L g2432 ( 
.A(n_2047),
.B(n_1967),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_2097),
.Y(n_2433)
);

AND2x2_ASAP7_75t_L g2434 ( 
.A(n_2084),
.B(n_911),
.Y(n_2434)
);

NOR2xp67_ASAP7_75t_SL g2435 ( 
.A(n_2069),
.B(n_1906),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2087),
.B(n_911),
.Y(n_2436)
);

CKINVDCx5p33_ASAP7_75t_R g2437 ( 
.A(n_2098),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_2088),
.B(n_912),
.Y(n_2438)
);

AOI22xp5_ASAP7_75t_L g2439 ( 
.A1(n_2185),
.A2(n_622),
.B1(n_625),
.B2(n_620),
.Y(n_2439)
);

OR2x2_ASAP7_75t_L g2440 ( 
.A(n_2129),
.B(n_1985),
.Y(n_2440)
);

AND3x1_ASAP7_75t_SL g2441 ( 
.A(n_2110),
.B(n_681),
.C(n_678),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2126),
.B(n_912),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2162),
.B(n_626),
.Y(n_2443)
);

BUFx6f_ASAP7_75t_L g2444 ( 
.A(n_2072),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2138),
.Y(n_2445)
);

OR2x2_ASAP7_75t_L g2446 ( 
.A(n_2220),
.B(n_1985),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_2153),
.B(n_2156),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2122),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2226),
.B(n_913),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2124),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2074),
.B(n_628),
.Y(n_2451)
);

AOI22xp5_ASAP7_75t_L g2452 ( 
.A1(n_2113),
.A2(n_634),
.B1(n_643),
.B2(n_632),
.Y(n_2452)
);

INVx4_ASAP7_75t_L g2453 ( 
.A(n_2115),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2140),
.B(n_913),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2125),
.Y(n_2455)
);

CKINVDCx5p33_ASAP7_75t_R g2456 ( 
.A(n_2128),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2159),
.B(n_645),
.Y(n_2457)
);

INVx4_ASAP7_75t_L g2458 ( 
.A(n_2132),
.Y(n_2458)
);

AOI22xp33_ASAP7_75t_SL g2459 ( 
.A1(n_2232),
.A2(n_681),
.B1(n_693),
.B2(n_678),
.Y(n_2459)
);

INVx3_ASAP7_75t_L g2460 ( 
.A(n_2139),
.Y(n_2460)
);

OAI22xp5_ASAP7_75t_L g2461 ( 
.A1(n_2197),
.A2(n_1961),
.B1(n_1910),
.B2(n_651),
.Y(n_2461)
);

INVx3_ASAP7_75t_L g2462 ( 
.A(n_2204),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2141),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2143),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_2175),
.B(n_647),
.Y(n_2465)
);

OR2x2_ASAP7_75t_L g2466 ( 
.A(n_2144),
.B(n_1910),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2145),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2147),
.B(n_659),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2148),
.B(n_914),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2149),
.Y(n_2470)
);

AND2x4_ASAP7_75t_L g2471 ( 
.A(n_2200),
.B(n_1961),
.Y(n_2471)
);

BUFx6f_ASAP7_75t_L g2472 ( 
.A(n_2201),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2202),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2203),
.B(n_914),
.Y(n_2474)
);

BUFx3_ASAP7_75t_L g2475 ( 
.A(n_2209),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2187),
.Y(n_2476)
);

AOI22xp33_ASAP7_75t_L g2477 ( 
.A1(n_2234),
.A2(n_698),
.B1(n_714),
.B2(n_693),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2188),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2205),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2206),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2207),
.B(n_915),
.Y(n_2481)
);

A2O1A1Ixp33_ASAP7_75t_L g2482 ( 
.A1(n_2233),
.A2(n_1395),
.B(n_756),
.C(n_770),
.Y(n_2482)
);

INVx3_ASAP7_75t_L g2483 ( 
.A(n_2211),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2208),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2189),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2210),
.B(n_662),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2213),
.B(n_665),
.Y(n_2487)
);

AOI22xp5_ASAP7_75t_L g2488 ( 
.A1(n_2214),
.A2(n_2219),
.B1(n_2218),
.B2(n_2192),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2196),
.B(n_669),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_SL g2490 ( 
.A(n_2191),
.B(n_1492),
.Y(n_2490)
);

INVx5_ASAP7_75t_L g2491 ( 
.A(n_2195),
.Y(n_2491)
);

OAI22xp5_ASAP7_75t_SL g2492 ( 
.A1(n_2006),
.A2(n_676),
.B1(n_683),
.B2(n_671),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2006),
.B(n_686),
.Y(n_2493)
);

AND2x2_ASAP7_75t_L g2494 ( 
.A(n_2003),
.B(n_915),
.Y(n_2494)
);

NAND3xp33_ASAP7_75t_SL g2495 ( 
.A(n_2048),
.B(n_689),
.C(n_687),
.Y(n_2495)
);

AND2x4_ASAP7_75t_L g2496 ( 
.A(n_2015),
.B(n_1275),
.Y(n_2496)
);

AOI22xp33_ASAP7_75t_L g2497 ( 
.A1(n_2081),
.A2(n_714),
.B1(n_722),
.B2(n_698),
.Y(n_2497)
);

NAND2x1p5_ASAP7_75t_L g2498 ( 
.A(n_2127),
.B(n_1258),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2118),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2006),
.B(n_690),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2056),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2006),
.B(n_694),
.Y(n_2502)
);

OAI221xp5_ASAP7_75t_L g2503 ( 
.A1(n_2048),
.A2(n_921),
.B1(n_923),
.B2(n_920),
.C(n_917),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_2021),
.Y(n_2504)
);

AOI22x1_ASAP7_75t_L g2505 ( 
.A1(n_2287),
.A2(n_727),
.B1(n_728),
.B2(n_722),
.Y(n_2505)
);

AO21x2_ASAP7_75t_L g2506 ( 
.A1(n_2447),
.A2(n_1395),
.B(n_1501),
.Y(n_2506)
);

BUFx2_ASAP7_75t_SL g2507 ( 
.A(n_2377),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2322),
.B(n_695),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2264),
.Y(n_2509)
);

INVx3_ASAP7_75t_L g2510 ( 
.A(n_2428),
.Y(n_2510)
);

INVxp67_ASAP7_75t_L g2511 ( 
.A(n_2246),
.Y(n_2511)
);

OAI21x1_ASAP7_75t_L g2512 ( 
.A1(n_2237),
.A2(n_1081),
.B(n_1079),
.Y(n_2512)
);

NAND2x1p5_ASAP7_75t_L g2513 ( 
.A(n_2447),
.B(n_2453),
.Y(n_2513)
);

AND2x4_ASAP7_75t_L g2514 ( 
.A(n_2405),
.B(n_1092),
.Y(n_2514)
);

AO21x2_ASAP7_75t_L g2515 ( 
.A1(n_2237),
.A2(n_837),
.B(n_836),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2264),
.Y(n_2516)
);

BUFx8_ASAP7_75t_SL g2517 ( 
.A(n_2238),
.Y(n_2517)
);

AOI22x1_ASAP7_75t_L g2518 ( 
.A1(n_2287),
.A2(n_728),
.B1(n_731),
.B2(n_727),
.Y(n_2518)
);

NOR2x1_ASAP7_75t_R g2519 ( 
.A(n_2239),
.B(n_699),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2266),
.Y(n_2520)
);

OAI21x1_ASAP7_75t_L g2521 ( 
.A1(n_2348),
.A2(n_2396),
.B(n_2399),
.Y(n_2521)
);

AO21x2_ASAP7_75t_L g2522 ( 
.A1(n_2406),
.A2(n_843),
.B(n_840),
.Y(n_2522)
);

INVx1_ASAP7_75t_SL g2523 ( 
.A(n_2249),
.Y(n_2523)
);

BUFx3_ASAP7_75t_L g2524 ( 
.A(n_2342),
.Y(n_2524)
);

AO21x2_ASAP7_75t_L g2525 ( 
.A1(n_2320),
.A2(n_2324),
.B(n_2359),
.Y(n_2525)
);

OAI21x1_ASAP7_75t_L g2526 ( 
.A1(n_2399),
.A2(n_1102),
.B(n_1092),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2266),
.Y(n_2527)
);

INVx8_ASAP7_75t_L g2528 ( 
.A(n_2496),
.Y(n_2528)
);

CKINVDCx14_ASAP7_75t_R g2529 ( 
.A(n_2238),
.Y(n_2529)
);

CKINVDCx11_ASAP7_75t_R g2530 ( 
.A(n_2254),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2330),
.B(n_700),
.Y(n_2531)
);

OAI21x1_ASAP7_75t_SL g2532 ( 
.A1(n_2256),
.A2(n_1278),
.B(n_1104),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2386),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2326),
.Y(n_2534)
);

OAI21x1_ASAP7_75t_SL g2535 ( 
.A1(n_2357),
.A2(n_1278),
.B(n_1104),
.Y(n_2535)
);

AO21x2_ASAP7_75t_L g2536 ( 
.A1(n_2320),
.A2(n_843),
.B(n_840),
.Y(n_2536)
);

NOR2x1_ASAP7_75t_L g2537 ( 
.A(n_2453),
.B(n_917),
.Y(n_2537)
);

OA21x2_ASAP7_75t_L g2538 ( 
.A1(n_2324),
.A2(n_848),
.B(n_846),
.Y(n_2538)
);

OA21x2_ASAP7_75t_L g2539 ( 
.A1(n_2374),
.A2(n_848),
.B(n_846),
.Y(n_2539)
);

BUFx6f_ASAP7_75t_L g2540 ( 
.A(n_2425),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2347),
.B(n_702),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2327),
.B(n_731),
.Y(n_2542)
);

AOI22x1_ASAP7_75t_L g2543 ( 
.A1(n_2267),
.A2(n_742),
.B1(n_748),
.B2(n_733),
.Y(n_2543)
);

CKINVDCx5p33_ASAP7_75t_R g2544 ( 
.A(n_2504),
.Y(n_2544)
);

BUFx4f_ASAP7_75t_L g2545 ( 
.A(n_2395),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2288),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2292),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2273),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2386),
.Y(n_2549)
);

INVx3_ASAP7_75t_L g2550 ( 
.A(n_2428),
.Y(n_2550)
);

AOI22xp33_ASAP7_75t_L g2551 ( 
.A1(n_2495),
.A2(n_742),
.B1(n_748),
.B2(n_733),
.Y(n_2551)
);

INVx3_ASAP7_75t_L g2552 ( 
.A(n_2401),
.Y(n_2552)
);

OAI21x1_ASAP7_75t_L g2553 ( 
.A1(n_2401),
.A2(n_1109),
.B(n_1102),
.Y(n_2553)
);

OAI21x1_ASAP7_75t_L g2554 ( 
.A1(n_2490),
.A2(n_1114),
.B(n_1109),
.Y(n_2554)
);

OA21x2_ASAP7_75t_L g2555 ( 
.A1(n_2374),
.A2(n_854),
.B(n_851),
.Y(n_2555)
);

AOI21xp5_ASAP7_75t_L g2556 ( 
.A1(n_2410),
.A2(n_1424),
.B(n_1398),
.Y(n_2556)
);

AO21x2_ASAP7_75t_L g2557 ( 
.A1(n_2410),
.A2(n_854),
.B(n_851),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2388),
.Y(n_2558)
);

INVx4_ASAP7_75t_L g2559 ( 
.A(n_2453),
.Y(n_2559)
);

INVxp67_ASAP7_75t_SL g2560 ( 
.A(n_2310),
.Y(n_2560)
);

NAND2x1p5_ASAP7_75t_L g2561 ( 
.A(n_2458),
.B(n_1258),
.Y(n_2561)
);

OAI21x1_ASAP7_75t_L g2562 ( 
.A1(n_2490),
.A2(n_1117),
.B(n_1114),
.Y(n_2562)
);

OR2x6_ASAP7_75t_L g2563 ( 
.A(n_2304),
.B(n_2458),
.Y(n_2563)
);

BUFx4f_ASAP7_75t_L g2564 ( 
.A(n_2395),
.Y(n_2564)
);

INVxp67_ASAP7_75t_L g2565 ( 
.A(n_2241),
.Y(n_2565)
);

INVx2_ASAP7_75t_SL g2566 ( 
.A(n_2362),
.Y(n_2566)
);

OAI21x1_ASAP7_75t_L g2567 ( 
.A1(n_2351),
.A2(n_1126),
.B(n_1117),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2388),
.Y(n_2568)
);

BUFx12f_ASAP7_75t_L g2569 ( 
.A(n_2504),
.Y(n_2569)
);

OAI21x1_ASAP7_75t_L g2570 ( 
.A1(n_2351),
.A2(n_1129),
.B(n_1126),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2281),
.Y(n_2571)
);

OAI21x1_ASAP7_75t_L g2572 ( 
.A1(n_2420),
.A2(n_1143),
.B(n_1129),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2296),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2323),
.B(n_751),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2318),
.Y(n_2575)
);

OAI21x1_ASAP7_75t_L g2576 ( 
.A1(n_2498),
.A2(n_1145),
.B(n_1143),
.Y(n_2576)
);

INVxp67_ASAP7_75t_L g2577 ( 
.A(n_2331),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2294),
.Y(n_2578)
);

AOI21xp5_ASAP7_75t_L g2579 ( 
.A1(n_2300),
.A2(n_1365),
.B(n_1333),
.Y(n_2579)
);

BUFx4f_ASAP7_75t_SL g2580 ( 
.A(n_2377),
.Y(n_2580)
);

INVx3_ASAP7_75t_L g2581 ( 
.A(n_2379),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2350),
.Y(n_2582)
);

AND2x4_ASAP7_75t_L g2583 ( 
.A(n_2405),
.B(n_1145),
.Y(n_2583)
);

INVx2_ASAP7_75t_SL g2584 ( 
.A(n_2362),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2421),
.Y(n_2585)
);

AND2x4_ASAP7_75t_L g2586 ( 
.A(n_2411),
.B(n_1148),
.Y(n_2586)
);

BUFx8_ASAP7_75t_SL g2587 ( 
.A(n_2340),
.Y(n_2587)
);

INVx2_ASAP7_75t_SL g2588 ( 
.A(n_2362),
.Y(n_2588)
);

OAI21x1_ASAP7_75t_L g2589 ( 
.A1(n_2498),
.A2(n_1149),
.B(n_1148),
.Y(n_2589)
);

OAI21x1_ASAP7_75t_L g2590 ( 
.A1(n_2462),
.A2(n_1153),
.B(n_1149),
.Y(n_2590)
);

INVx1_ASAP7_75t_SL g2591 ( 
.A(n_2249),
.Y(n_2591)
);

OAI21x1_ASAP7_75t_L g2592 ( 
.A1(n_2462),
.A2(n_1154),
.B(n_1153),
.Y(n_2592)
);

BUFx12f_ASAP7_75t_L g2593 ( 
.A(n_2340),
.Y(n_2593)
);

OAI21x1_ASAP7_75t_L g2594 ( 
.A1(n_2483),
.A2(n_1158),
.B(n_1154),
.Y(n_2594)
);

OAI21xp5_ASAP7_75t_L g2595 ( 
.A1(n_2369),
.A2(n_756),
.B(n_751),
.Y(n_2595)
);

AO21x2_ASAP7_75t_L g2596 ( 
.A1(n_2278),
.A2(n_2364),
.B(n_2482),
.Y(n_2596)
);

BUFx3_ASAP7_75t_L g2597 ( 
.A(n_2342),
.Y(n_2597)
);

AO21x2_ASAP7_75t_L g2598 ( 
.A1(n_2364),
.A2(n_867),
.B(n_865),
.Y(n_2598)
);

OAI21x1_ASAP7_75t_L g2599 ( 
.A1(n_2483),
.A2(n_1165),
.B(n_1158),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2379),
.B(n_770),
.Y(n_2600)
);

AND2x4_ASAP7_75t_L g2601 ( 
.A(n_2411),
.B(n_2379),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2257),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2268),
.Y(n_2603)
);

INVx2_ASAP7_75t_SL g2604 ( 
.A(n_2393),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_2267),
.B(n_704),
.Y(n_2605)
);

OAI21x1_ASAP7_75t_L g2606 ( 
.A1(n_2344),
.A2(n_1169),
.B(n_1165),
.Y(n_2606)
);

OAI22xp5_ASAP7_75t_L g2607 ( 
.A1(n_2239),
.A2(n_711),
.B1(n_713),
.B2(n_709),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2258),
.Y(n_2608)
);

INVx3_ASAP7_75t_L g2609 ( 
.A(n_2379),
.Y(n_2609)
);

AO21x2_ASAP7_75t_L g2610 ( 
.A1(n_2482),
.A2(n_867),
.B(n_865),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2385),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2268),
.Y(n_2612)
);

INVx3_ASAP7_75t_L g2613 ( 
.A(n_2297),
.Y(n_2613)
);

AO21x2_ASAP7_75t_L g2614 ( 
.A1(n_2427),
.A2(n_870),
.B(n_868),
.Y(n_2614)
);

BUFx12f_ASAP7_75t_L g2615 ( 
.A(n_2240),
.Y(n_2615)
);

INVx3_ASAP7_75t_L g2616 ( 
.A(n_2297),
.Y(n_2616)
);

AOI21xp5_ASAP7_75t_L g2617 ( 
.A1(n_2300),
.A2(n_2316),
.B(n_2427),
.Y(n_2617)
);

INVx3_ASAP7_75t_L g2618 ( 
.A(n_2297),
.Y(n_2618)
);

OAI21x1_ASAP7_75t_L g2619 ( 
.A1(n_2370),
.A2(n_1169),
.B(n_1170),
.Y(n_2619)
);

CKINVDCx14_ASAP7_75t_R g2620 ( 
.A(n_2245),
.Y(n_2620)
);

NOR2xp33_ASAP7_75t_SL g2621 ( 
.A(n_2259),
.B(n_715),
.Y(n_2621)
);

OAI21x1_ASAP7_75t_L g2622 ( 
.A1(n_2370),
.A2(n_1170),
.B(n_1260),
.Y(n_2622)
);

AOI22x1_ASAP7_75t_L g2623 ( 
.A1(n_2458),
.A2(n_788),
.B1(n_776),
.B2(n_719),
.Y(n_2623)
);

INVx3_ASAP7_75t_L g2624 ( 
.A(n_2393),
.Y(n_2624)
);

BUFx2_ASAP7_75t_L g2625 ( 
.A(n_2361),
.Y(n_2625)
);

BUFx6f_ASAP7_75t_L g2626 ( 
.A(n_2425),
.Y(n_2626)
);

OAI21x1_ASAP7_75t_L g2627 ( 
.A1(n_2389),
.A2(n_1264),
.B(n_1260),
.Y(n_2627)
);

AOI21xp5_ASAP7_75t_L g2628 ( 
.A1(n_2279),
.A2(n_1365),
.B(n_1333),
.Y(n_2628)
);

OAI21x1_ASAP7_75t_L g2629 ( 
.A1(n_2389),
.A2(n_1267),
.B(n_1264),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2271),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2307),
.B(n_776),
.Y(n_2631)
);

OAI21x1_ASAP7_75t_L g2632 ( 
.A1(n_2460),
.A2(n_1272),
.B(n_1089),
.Y(n_2632)
);

OAI21x1_ASAP7_75t_L g2633 ( 
.A1(n_2460),
.A2(n_1089),
.B(n_1069),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2394),
.B(n_716),
.Y(n_2634)
);

BUFx2_ASAP7_75t_SL g2635 ( 
.A(n_2402),
.Y(n_2635)
);

BUFx3_ASAP7_75t_L g2636 ( 
.A(n_2342),
.Y(n_2636)
);

AOI22x1_ASAP7_75t_L g2637 ( 
.A1(n_2433),
.A2(n_788),
.B1(n_723),
.B2(n_729),
.Y(n_2637)
);

BUFx12f_ASAP7_75t_L g2638 ( 
.A(n_2240),
.Y(n_2638)
);

AOI22x1_ASAP7_75t_L g2639 ( 
.A1(n_2433),
.A2(n_730),
.B1(n_736),
.B2(n_721),
.Y(n_2639)
);

OAI21x1_ASAP7_75t_L g2640 ( 
.A1(n_2271),
.A2(n_1089),
.B(n_1069),
.Y(n_2640)
);

CKINVDCx20_ASAP7_75t_R g2641 ( 
.A(n_2345),
.Y(n_2641)
);

INVx4_ASAP7_75t_L g2642 ( 
.A(n_2475),
.Y(n_2642)
);

NAND2x1p5_ASAP7_75t_L g2643 ( 
.A(n_2475),
.B(n_1204),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2284),
.Y(n_2644)
);

INVx1_ASAP7_75t_SL g2645 ( 
.A(n_2235),
.Y(n_2645)
);

BUFx12f_ASAP7_75t_L g2646 ( 
.A(n_2289),
.Y(n_2646)
);

OAI21x1_ASAP7_75t_L g2647 ( 
.A1(n_2284),
.A2(n_1090),
.B(n_1069),
.Y(n_2647)
);

BUFx2_ASAP7_75t_SL g2648 ( 
.A(n_2402),
.Y(n_2648)
);

AO21x2_ASAP7_75t_L g2649 ( 
.A1(n_2321),
.A2(n_2488),
.B(n_2332),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2291),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_2245),
.Y(n_2651)
);

AO21x2_ASAP7_75t_L g2652 ( 
.A1(n_2321),
.A2(n_870),
.B(n_868),
.Y(n_2652)
);

INVx5_ASAP7_75t_L g2653 ( 
.A(n_2393),
.Y(n_2653)
);

BUFx2_ASAP7_75t_L g2654 ( 
.A(n_2349),
.Y(n_2654)
);

INVx2_ASAP7_75t_SL g2655 ( 
.A(n_2275),
.Y(n_2655)
);

OAI21x1_ASAP7_75t_L g2656 ( 
.A1(n_2291),
.A2(n_1090),
.B(n_872),
.Y(n_2656)
);

OAI21x1_ASAP7_75t_L g2657 ( 
.A1(n_2302),
.A2(n_1090),
.B(n_872),
.Y(n_2657)
);

INVx3_ASAP7_75t_L g2658 ( 
.A(n_2471),
.Y(n_2658)
);

BUFx6f_ASAP7_75t_L g2659 ( 
.A(n_2275),
.Y(n_2659)
);

HB1xp67_ASAP7_75t_L g2660 ( 
.A(n_2236),
.Y(n_2660)
);

INVx1_ASAP7_75t_SL g2661 ( 
.A(n_2276),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2302),
.Y(n_2662)
);

INVx2_ASAP7_75t_SL g2663 ( 
.A(n_2286),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2339),
.Y(n_2664)
);

INVxp67_ASAP7_75t_SL g2665 ( 
.A(n_2312),
.Y(n_2665)
);

INVx3_ASAP7_75t_L g2666 ( 
.A(n_2471),
.Y(n_2666)
);

AO21x2_ASAP7_75t_L g2667 ( 
.A1(n_2280),
.A2(n_2325),
.B(n_2295),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2339),
.Y(n_2668)
);

BUFx3_ASAP7_75t_L g2669 ( 
.A(n_2349),
.Y(n_2669)
);

NAND2x1p5_ASAP7_75t_L g2670 ( 
.A(n_2491),
.B(n_1204),
.Y(n_2670)
);

INVx3_ASAP7_75t_L g2671 ( 
.A(n_2471),
.Y(n_2671)
);

HB1xp67_ASAP7_75t_L g2672 ( 
.A(n_2247),
.Y(n_2672)
);

CKINVDCx5p33_ASAP7_75t_R g2673 ( 
.A(n_2289),
.Y(n_2673)
);

INVx6_ASAP7_75t_L g2674 ( 
.A(n_2349),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2315),
.B(n_739),
.Y(n_2675)
);

OAI21x1_ASAP7_75t_SL g2676 ( 
.A1(n_2391),
.A2(n_877),
.B(n_871),
.Y(n_2676)
);

BUFx6f_ASAP7_75t_L g2677 ( 
.A(n_2286),
.Y(n_2677)
);

BUFx3_ASAP7_75t_L g2678 ( 
.A(n_2356),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2354),
.Y(n_2679)
);

AO21x2_ASAP7_75t_L g2680 ( 
.A1(n_2280),
.A2(n_877),
.B(n_871),
.Y(n_2680)
);

BUFx6f_ASAP7_75t_L g2681 ( 
.A(n_2328),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2354),
.Y(n_2682)
);

OAI21xp5_ASAP7_75t_L g2683 ( 
.A1(n_2465),
.A2(n_744),
.B(n_741),
.Y(n_2683)
);

OAI21x1_ASAP7_75t_L g2684 ( 
.A1(n_2360),
.A2(n_1034),
.B(n_1018),
.Y(n_2684)
);

AO21x2_ASAP7_75t_L g2685 ( 
.A1(n_2333),
.A2(n_921),
.B(n_920),
.Y(n_2685)
);

OAI21x1_ASAP7_75t_L g2686 ( 
.A1(n_2360),
.A2(n_1034),
.B(n_1018),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2261),
.B(n_745),
.Y(n_2687)
);

INVx1_ASAP7_75t_SL g2688 ( 
.A(n_2494),
.Y(n_2688)
);

OAI21x1_ASAP7_75t_L g2689 ( 
.A1(n_2367),
.A2(n_1034),
.B(n_1018),
.Y(n_2689)
);

AO21x2_ASAP7_75t_L g2690 ( 
.A1(n_2290),
.A2(n_924),
.B(n_923),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2303),
.B(n_2269),
.Y(n_2691)
);

BUFx6f_ASAP7_75t_L g2692 ( 
.A(n_2328),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2367),
.Y(n_2693)
);

INVx1_ASAP7_75t_SL g2694 ( 
.A(n_2272),
.Y(n_2694)
);

BUFx3_ASAP7_75t_L g2695 ( 
.A(n_2356),
.Y(n_2695)
);

HB1xp67_ASAP7_75t_L g2696 ( 
.A(n_2251),
.Y(n_2696)
);

OA21x2_ASAP7_75t_L g2697 ( 
.A1(n_2382),
.A2(n_925),
.B(n_924),
.Y(n_2697)
);

NOR2xp33_ASAP7_75t_L g2698 ( 
.A(n_2493),
.B(n_747),
.Y(n_2698)
);

HB1xp67_ASAP7_75t_L g2699 ( 
.A(n_2253),
.Y(n_2699)
);

AND2x2_ASAP7_75t_SL g2700 ( 
.A(n_2307),
.B(n_925),
.Y(n_2700)
);

INVx2_ASAP7_75t_SL g2701 ( 
.A(n_2444),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2372),
.Y(n_2702)
);

BUFx2_ASAP7_75t_L g2703 ( 
.A(n_2356),
.Y(n_2703)
);

INVxp67_ASAP7_75t_SL g2704 ( 
.A(n_2248),
.Y(n_2704)
);

BUFx2_ASAP7_75t_L g2705 ( 
.A(n_2408),
.Y(n_2705)
);

OAI21x1_ASAP7_75t_L g2706 ( 
.A1(n_2372),
.A2(n_1034),
.B(n_992),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_SL g2707 ( 
.A(n_2244),
.B(n_927),
.Y(n_2707)
);

OAI21x1_ASAP7_75t_L g2708 ( 
.A1(n_2476),
.A2(n_2485),
.B(n_2478),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2248),
.Y(n_2709)
);

INVx3_ASAP7_75t_L g2710 ( 
.A(n_2446),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_2250),
.Y(n_2711)
);

NAND2x1p5_ASAP7_75t_L g2712 ( 
.A(n_2491),
.B(n_1216),
.Y(n_2712)
);

OAI21x1_ASAP7_75t_L g2713 ( 
.A1(n_2476),
.A2(n_992),
.B(n_991),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2250),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2262),
.Y(n_2715)
);

CKINVDCx11_ASAP7_75t_R g2716 ( 
.A(n_2345),
.Y(n_2716)
);

INVx2_ASAP7_75t_SL g2717 ( 
.A(n_2444),
.Y(n_2717)
);

AO21x2_ASAP7_75t_L g2718 ( 
.A1(n_2290),
.A2(n_929),
.B(n_927),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2262),
.Y(n_2719)
);

OAI21x1_ASAP7_75t_L g2720 ( 
.A1(n_2478),
.A2(n_1016),
.B(n_991),
.Y(n_2720)
);

AOI22x1_ASAP7_75t_L g2721 ( 
.A1(n_2437),
.A2(n_757),
.B1(n_759),
.B2(n_755),
.Y(n_2721)
);

INVx2_ASAP7_75t_SL g2722 ( 
.A(n_2444),
.Y(n_2722)
);

INVx1_ASAP7_75t_SL g2723 ( 
.A(n_2277),
.Y(n_2723)
);

AO21x2_ASAP7_75t_L g2724 ( 
.A1(n_2378),
.A2(n_930),
.B(n_929),
.Y(n_2724)
);

OAI21x1_ASAP7_75t_L g2725 ( 
.A1(n_2485),
.A2(n_1028),
.B(n_1016),
.Y(n_2725)
);

OAI21x1_ASAP7_75t_L g2726 ( 
.A1(n_2429),
.A2(n_1029),
.B(n_1028),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2499),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2499),
.Y(n_2728)
);

INVx4_ASAP7_75t_L g2729 ( 
.A(n_2444),
.Y(n_2729)
);

BUFx3_ASAP7_75t_L g2730 ( 
.A(n_2255),
.Y(n_2730)
);

AND2x4_ASAP7_75t_L g2731 ( 
.A(n_2255),
.B(n_365),
.Y(n_2731)
);

INVx3_ASAP7_75t_L g2732 ( 
.A(n_2432),
.Y(n_2732)
);

NAND2x1p5_ASAP7_75t_L g2733 ( 
.A(n_2491),
.B(n_1218),
.Y(n_2733)
);

INVx1_ASAP7_75t_SL g2734 ( 
.A(n_2424),
.Y(n_2734)
);

AO21x2_ASAP7_75t_L g2735 ( 
.A1(n_2443),
.A2(n_932),
.B(n_930),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2384),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2397),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2397),
.Y(n_2738)
);

BUFx6f_ASAP7_75t_L g2739 ( 
.A(n_2242),
.Y(n_2739)
);

INVx1_ASAP7_75t_SL g2740 ( 
.A(n_2424),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2263),
.Y(n_2741)
);

INVx5_ASAP7_75t_SL g2742 ( 
.A(n_2472),
.Y(n_2742)
);

INVx2_ASAP7_75t_SL g2743 ( 
.A(n_2407),
.Y(n_2743)
);

HB1xp67_ASAP7_75t_L g2744 ( 
.A(n_2501),
.Y(n_2744)
);

NAND2x1p5_ASAP7_75t_L g2745 ( 
.A(n_2491),
.B(n_1218),
.Y(n_2745)
);

AND2x2_ASAP7_75t_SL g2746 ( 
.A(n_2497),
.B(n_932),
.Y(n_2746)
);

BUFx2_ASAP7_75t_R g2747 ( 
.A(n_2334),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2358),
.Y(n_2748)
);

AO21x2_ASAP7_75t_L g2749 ( 
.A1(n_2418),
.A2(n_938),
.B(n_935),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2363),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2335),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2343),
.Y(n_2752)
);

BUFx3_ASAP7_75t_L g2753 ( 
.A(n_2353),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2346),
.Y(n_2754)
);

OAI21x1_ASAP7_75t_L g2755 ( 
.A1(n_2429),
.A2(n_1031),
.B(n_1029),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2431),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2431),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2440),
.Y(n_2758)
);

AND2x2_ASAP7_75t_L g2759 ( 
.A(n_2314),
.B(n_935),
.Y(n_2759)
);

AO21x2_ASAP7_75t_L g2760 ( 
.A1(n_2419),
.A2(n_938),
.B(n_971),
.Y(n_2760)
);

OAI21x1_ASAP7_75t_L g2761 ( 
.A1(n_2448),
.A2(n_1054),
.B(n_1031),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2448),
.Y(n_2762)
);

BUFx3_ASAP7_75t_L g2763 ( 
.A(n_2437),
.Y(n_2763)
);

BUFx4_ASAP7_75t_SL g2764 ( 
.A(n_2334),
.Y(n_2764)
);

NOR2xp33_ASAP7_75t_L g2765 ( 
.A(n_2500),
.B(n_761),
.Y(n_2765)
);

AND2x4_ASAP7_75t_L g2766 ( 
.A(n_2242),
.B(n_366),
.Y(n_2766)
);

BUFx4f_ASAP7_75t_SL g2767 ( 
.A(n_2283),
.Y(n_2767)
);

OAI21x1_ASAP7_75t_L g2768 ( 
.A1(n_2450),
.A2(n_1054),
.B(n_976),
.Y(n_2768)
);

INVx6_ASAP7_75t_L g2769 ( 
.A(n_2242),
.Y(n_2769)
);

AOI22xp33_ASAP7_75t_L g2770 ( 
.A1(n_2700),
.A2(n_2265),
.B1(n_2497),
.B2(n_2459),
.Y(n_2770)
);

AOI22xp33_ASAP7_75t_L g2771 ( 
.A1(n_2700),
.A2(n_2595),
.B1(n_2265),
.B2(n_2746),
.Y(n_2771)
);

OAI22xp5_ASAP7_75t_SL g2772 ( 
.A1(n_2700),
.A2(n_2260),
.B1(n_2338),
.B2(n_2341),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2751),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2751),
.Y(n_2774)
);

BUFx4_ASAP7_75t_SL g2775 ( 
.A(n_2641),
.Y(n_2775)
);

INVx6_ASAP7_75t_L g2776 ( 
.A(n_2642),
.Y(n_2776)
);

AOI22xp33_ASAP7_75t_L g2777 ( 
.A1(n_2545),
.A2(n_2365),
.B1(n_2243),
.B2(n_2329),
.Y(n_2777)
);

AOI22xp33_ASAP7_75t_L g2778 ( 
.A1(n_2746),
.A2(n_2317),
.B1(n_2376),
.B2(n_2282),
.Y(n_2778)
);

OAI22xp33_ASAP7_75t_R g2779 ( 
.A1(n_2698),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_2779)
);

INVx8_ASAP7_75t_L g2780 ( 
.A(n_2569),
.Y(n_2780)
);

OAI22xp33_ASAP7_75t_L g2781 ( 
.A1(n_2545),
.A2(n_2338),
.B1(n_2417),
.B2(n_2439),
.Y(n_2781)
);

BUFx6f_ASAP7_75t_L g2782 ( 
.A(n_2626),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2752),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2752),
.Y(n_2784)
);

OAI21xp5_ASAP7_75t_SL g2785 ( 
.A1(n_2631),
.A2(n_2305),
.B(n_2317),
.Y(n_2785)
);

INVx1_ASAP7_75t_SL g2786 ( 
.A(n_2523),
.Y(n_2786)
);

BUFx12f_ASAP7_75t_L g2787 ( 
.A(n_2651),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2754),
.Y(n_2788)
);

OAI22xp5_ASAP7_75t_L g2789 ( 
.A1(n_2577),
.A2(n_2313),
.B1(n_2305),
.B2(n_2376),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2754),
.Y(n_2790)
);

OAI22xp33_ASAP7_75t_L g2791 ( 
.A1(n_2545),
.A2(n_2456),
.B1(n_2252),
.B2(n_2352),
.Y(n_2791)
);

OAI22xp5_ASAP7_75t_L g2792 ( 
.A1(n_2564),
.A2(n_2456),
.B1(n_2375),
.B2(n_2355),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2758),
.Y(n_2793)
);

OAI22xp33_ASAP7_75t_L g2794 ( 
.A1(n_2564),
.A2(n_2457),
.B1(n_2375),
.B2(n_2452),
.Y(n_2794)
);

AND2x2_ASAP7_75t_L g2795 ( 
.A(n_2625),
.B(n_2368),
.Y(n_2795)
);

AOI22xp33_ASAP7_75t_SL g2796 ( 
.A1(n_2631),
.A2(n_2329),
.B1(n_2382),
.B2(n_2492),
.Y(n_2796)
);

AOI22xp33_ASAP7_75t_L g2797 ( 
.A1(n_2746),
.A2(n_2477),
.B1(n_2392),
.B2(n_2414),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2758),
.Y(n_2798)
);

INVx5_ASAP7_75t_L g2799 ( 
.A(n_2674),
.Y(n_2799)
);

CKINVDCx16_ASAP7_75t_R g2800 ( 
.A(n_2615),
.Y(n_2800)
);

AOI22xp5_ASAP7_75t_L g2801 ( 
.A1(n_2511),
.A2(n_2319),
.B1(n_2299),
.B2(n_2398),
.Y(n_2801)
);

INVx2_ASAP7_75t_SL g2802 ( 
.A(n_2764),
.Y(n_2802)
);

AOI22xp33_ASAP7_75t_SL g2803 ( 
.A1(n_2564),
.A2(n_2309),
.B1(n_2503),
.B2(n_2387),
.Y(n_2803)
);

CKINVDCx5p33_ASAP7_75t_R g2804 ( 
.A(n_2517),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2585),
.B(n_2422),
.Y(n_2805)
);

OAI22xp5_ASAP7_75t_L g2806 ( 
.A1(n_2591),
.A2(n_2477),
.B1(n_2392),
.B2(n_2371),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2534),
.Y(n_2807)
);

BUFx2_ASAP7_75t_L g2808 ( 
.A(n_2626),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2578),
.Y(n_2809)
);

INVx8_ASAP7_75t_L g2810 ( 
.A(n_2569),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2534),
.Y(n_2811)
);

INVx4_ASAP7_75t_L g2812 ( 
.A(n_2626),
.Y(n_2812)
);

OAI22x1_ASAP7_75t_L g2813 ( 
.A1(n_2565),
.A2(n_2423),
.B1(n_2293),
.B2(n_2430),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2578),
.Y(n_2814)
);

OAI22xp33_ASAP7_75t_L g2815 ( 
.A1(n_2688),
.A2(n_2274),
.B1(n_2311),
.B2(n_2285),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2582),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2582),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2736),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2736),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2736),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2738),
.Y(n_2821)
);

BUFx2_ASAP7_75t_SL g2822 ( 
.A(n_2763),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2548),
.Y(n_2823)
);

AOI22xp33_ASAP7_75t_L g2824 ( 
.A1(n_2623),
.A2(n_2380),
.B1(n_2496),
.B2(n_2449),
.Y(n_2824)
);

CKINVDCx20_ASAP7_75t_R g2825 ( 
.A(n_2530),
.Y(n_2825)
);

BUFx12f_ASAP7_75t_L g2826 ( 
.A(n_2544),
.Y(n_2826)
);

CKINVDCx11_ASAP7_75t_R g2827 ( 
.A(n_2716),
.Y(n_2827)
);

BUFx10_ASAP7_75t_L g2828 ( 
.A(n_2605),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2738),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2548),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2625),
.B(n_2301),
.Y(n_2831)
);

AOI22xp5_ASAP7_75t_L g2832 ( 
.A1(n_2707),
.A2(n_2319),
.B1(n_2441),
.B2(n_2381),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2571),
.Y(n_2833)
);

AOI22xp33_ASAP7_75t_L g2834 ( 
.A1(n_2623),
.A2(n_2496),
.B1(n_2306),
.B2(n_2472),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2571),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2645),
.B(n_2434),
.Y(n_2836)
);

AOI22xp33_ASAP7_75t_L g2837 ( 
.A1(n_2765),
.A2(n_2753),
.B1(n_2525),
.B2(n_2540),
.Y(n_2837)
);

AOI21xp5_ASAP7_75t_L g2838 ( 
.A1(n_2579),
.A2(n_2270),
.B(n_2336),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2585),
.B(n_2502),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2575),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2738),
.Y(n_2841)
);

CKINVDCx8_ASAP7_75t_R g2842 ( 
.A(n_2635),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2575),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2737),
.Y(n_2844)
);

CKINVDCx20_ASAP7_75t_R g2845 ( 
.A(n_2580),
.Y(n_2845)
);

OAI22x1_ASAP7_75t_SL g2846 ( 
.A1(n_2673),
.A2(n_765),
.B1(n_766),
.B2(n_763),
.Y(n_2846)
);

BUFx12f_ASAP7_75t_L g2847 ( 
.A(n_2646),
.Y(n_2847)
);

AOI22xp33_ASAP7_75t_L g2848 ( 
.A1(n_2753),
.A2(n_2472),
.B1(n_2416),
.B2(n_2373),
.Y(n_2848)
);

BUFx8_ASAP7_75t_SL g2849 ( 
.A(n_2587),
.Y(n_2849)
);

OAI22x1_ASAP7_75t_L g2850 ( 
.A1(n_2705),
.A2(n_2479),
.B1(n_2480),
.B2(n_2473),
.Y(n_2850)
);

CKINVDCx11_ASAP7_75t_R g2851 ( 
.A(n_2615),
.Y(n_2851)
);

AND2x2_ASAP7_75t_L g2852 ( 
.A(n_2705),
.B(n_2436),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2753),
.B(n_2613),
.Y(n_2853)
);

CKINVDCx5p33_ASAP7_75t_R g2854 ( 
.A(n_2529),
.Y(n_2854)
);

BUFx3_ASAP7_75t_L g2855 ( 
.A(n_2593),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2737),
.Y(n_2856)
);

OAI21xp5_ASAP7_75t_SL g2857 ( 
.A1(n_2551),
.A2(n_2366),
.B(n_2383),
.Y(n_2857)
);

AOI22xp33_ASAP7_75t_L g2858 ( 
.A1(n_2543),
.A2(n_2337),
.B1(n_2438),
.B2(n_2409),
.Y(n_2858)
);

INVx1_ASAP7_75t_SL g2859 ( 
.A(n_2661),
.Y(n_2859)
);

CKINVDCx11_ASAP7_75t_R g2860 ( 
.A(n_2638),
.Y(n_2860)
);

AOI22xp33_ASAP7_75t_L g2861 ( 
.A1(n_2543),
.A2(n_2404),
.B1(n_2442),
.B2(n_2390),
.Y(n_2861)
);

CKINVDCx6p67_ASAP7_75t_R g2862 ( 
.A(n_2638),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2573),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2573),
.Y(n_2864)
);

AOI22xp33_ASAP7_75t_SL g2865 ( 
.A1(n_2525),
.A2(n_2400),
.B1(n_2381),
.B2(n_2403),
.Y(n_2865)
);

INVx6_ASAP7_75t_L g2866 ( 
.A(n_2642),
.Y(n_2866)
);

AOI22xp5_ASAP7_75t_L g2867 ( 
.A1(n_2621),
.A2(n_2767),
.B1(n_2525),
.B2(n_2620),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2723),
.B(n_2665),
.Y(n_2868)
);

AOI22xp33_ASAP7_75t_L g2869 ( 
.A1(n_2540),
.A2(n_2472),
.B1(n_2481),
.B2(n_2474),
.Y(n_2869)
);

OAI22xp33_ASAP7_75t_L g2870 ( 
.A1(n_2505),
.A2(n_2298),
.B1(n_2308),
.B2(n_2484),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2573),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2560),
.B(n_2691),
.Y(n_2872)
);

BUFx8_ASAP7_75t_L g2873 ( 
.A(n_2646),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2667),
.B(n_2412),
.Y(n_2874)
);

AOI22xp33_ASAP7_75t_L g2875 ( 
.A1(n_2505),
.A2(n_772),
.B1(n_773),
.B2(n_769),
.Y(n_2875)
);

INVx6_ASAP7_75t_L g2876 ( 
.A(n_2642),
.Y(n_2876)
);

HB1xp67_ASAP7_75t_L g2877 ( 
.A(n_2667),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2667),
.B(n_2413),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2732),
.Y(n_2879)
);

AOI22xp33_ASAP7_75t_L g2880 ( 
.A1(n_2518),
.A2(n_782),
.B1(n_783),
.B2(n_779),
.Y(n_2880)
);

BUFx4f_ASAP7_75t_SL g2881 ( 
.A(n_2593),
.Y(n_2881)
);

AOI22xp33_ASAP7_75t_L g2882 ( 
.A1(n_2540),
.A2(n_2435),
.B1(n_2451),
.B2(n_2486),
.Y(n_2882)
);

BUFx2_ASAP7_75t_L g2883 ( 
.A(n_2626),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2732),
.B(n_2415),
.Y(n_2884)
);

CKINVDCx5p33_ASAP7_75t_R g2885 ( 
.A(n_2507),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2741),
.Y(n_2886)
);

AOI22xp5_ASAP7_75t_L g2887 ( 
.A1(n_2596),
.A2(n_2441),
.B1(n_2487),
.B2(n_2489),
.Y(n_2887)
);

INVx1_ASAP7_75t_SL g2888 ( 
.A(n_2734),
.Y(n_2888)
);

INVx3_ASAP7_75t_L g2889 ( 
.A(n_2540),
.Y(n_2889)
);

AOI22xp33_ASAP7_75t_L g2890 ( 
.A1(n_2540),
.A2(n_2637),
.B1(n_2626),
.B2(n_2596),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2732),
.Y(n_2891)
);

BUFx3_ASAP7_75t_L g2892 ( 
.A(n_2763),
.Y(n_2892)
);

CKINVDCx20_ASAP7_75t_R g2893 ( 
.A(n_2763),
.Y(n_2893)
);

BUFx6f_ASAP7_75t_L g2894 ( 
.A(n_2540),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2732),
.Y(n_2895)
);

BUFx3_ASAP7_75t_L g2896 ( 
.A(n_2654),
.Y(n_2896)
);

AOI22xp33_ASAP7_75t_L g2897 ( 
.A1(n_2637),
.A2(n_2426),
.B1(n_2468),
.B2(n_2454),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2756),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2756),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2756),
.Y(n_2900)
);

INVx3_ASAP7_75t_L g2901 ( 
.A(n_2729),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2757),
.Y(n_2902)
);

AOI21xp5_ASAP7_75t_L g2903 ( 
.A1(n_2617),
.A2(n_2461),
.B(n_2455),
.Y(n_2903)
);

OAI22xp5_ASAP7_75t_SL g2904 ( 
.A1(n_2507),
.A2(n_785),
.B1(n_787),
.B2(n_784),
.Y(n_2904)
);

BUFx3_ASAP7_75t_L g2905 ( 
.A(n_2654),
.Y(n_2905)
);

AOI22xp33_ASAP7_75t_L g2906 ( 
.A1(n_2518),
.A2(n_2469),
.B1(n_2450),
.B2(n_2455),
.Y(n_2906)
);

OAI22xp5_ASAP7_75t_L g2907 ( 
.A1(n_2675),
.A2(n_2466),
.B1(n_2463),
.B2(n_2464),
.Y(n_2907)
);

CKINVDCx11_ASAP7_75t_R g2908 ( 
.A(n_2740),
.Y(n_2908)
);

OAI22xp5_ASAP7_75t_L g2909 ( 
.A1(n_2635),
.A2(n_2467),
.B1(n_2470),
.B2(n_2445),
.Y(n_2909)
);

BUFx3_ASAP7_75t_L g2910 ( 
.A(n_2703),
.Y(n_2910)
);

CKINVDCx20_ASAP7_75t_R g2911 ( 
.A(n_2648),
.Y(n_2911)
);

INVx4_ASAP7_75t_L g2912 ( 
.A(n_2642),
.Y(n_2912)
);

CKINVDCx11_ASAP7_75t_R g2913 ( 
.A(n_2703),
.Y(n_2913)
);

AOI22xp33_ASAP7_75t_SL g2914 ( 
.A1(n_2649),
.A2(n_5),
.B1(n_1),
.B2(n_2),
.Y(n_2914)
);

AOI22xp33_ASAP7_75t_SL g2915 ( 
.A1(n_2649),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2757),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2757),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2762),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2762),
.Y(n_2919)
);

AND2x2_ASAP7_75t_L g2920 ( 
.A(n_2613),
.B(n_9),
.Y(n_2920)
);

AOI22xp33_ASAP7_75t_L g2921 ( 
.A1(n_2596),
.A2(n_1045),
.B1(n_1056),
.B2(n_1040),
.Y(n_2921)
);

CKINVDCx11_ASAP7_75t_R g2922 ( 
.A(n_2694),
.Y(n_2922)
);

AOI21xp33_ASAP7_75t_L g2923 ( 
.A1(n_2649),
.A2(n_1056),
.B(n_1045),
.Y(n_2923)
);

OAI22xp5_ASAP7_75t_L g2924 ( 
.A1(n_2648),
.A2(n_1239),
.B1(n_1262),
.B2(n_1218),
.Y(n_2924)
);

BUFx2_ASAP7_75t_SL g2925 ( 
.A(n_2743),
.Y(n_2925)
);

AOI22xp33_ASAP7_75t_L g2926 ( 
.A1(n_2658),
.A2(n_1056),
.B1(n_1045),
.B2(n_976),
.Y(n_2926)
);

BUFx8_ASAP7_75t_SL g2927 ( 
.A(n_2524),
.Y(n_2927)
);

CKINVDCx20_ASAP7_75t_R g2928 ( 
.A(n_2524),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2762),
.Y(n_2929)
);

BUFx2_ASAP7_75t_L g2930 ( 
.A(n_2601),
.Y(n_2930)
);

AND2x4_ASAP7_75t_SL g2931 ( 
.A(n_2659),
.B(n_1045),
.Y(n_2931)
);

OAI22xp5_ASAP7_75t_L g2932 ( 
.A1(n_2747),
.A2(n_1239),
.B1(n_1262),
.B2(n_1218),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2546),
.Y(n_2933)
);

BUFx2_ASAP7_75t_L g2934 ( 
.A(n_2601),
.Y(n_2934)
);

BUFx10_ASAP7_75t_L g2935 ( 
.A(n_2766),
.Y(n_2935)
);

AND2x2_ASAP7_75t_L g2936 ( 
.A(n_2613),
.B(n_10),
.Y(n_2936)
);

OAI22xp5_ASAP7_75t_L g2937 ( 
.A1(n_2513),
.A2(n_1239),
.B1(n_1262),
.B2(n_1218),
.Y(n_2937)
);

AOI22xp33_ASAP7_75t_SL g2938 ( 
.A1(n_2652),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_2938)
);

BUFx12f_ASAP7_75t_L g2939 ( 
.A(n_2600),
.Y(n_2939)
);

OAI22xp5_ASAP7_75t_L g2940 ( 
.A1(n_2513),
.A2(n_2563),
.B1(n_2663),
.B2(n_2655),
.Y(n_2940)
);

AOI22xp33_ASAP7_75t_L g2941 ( 
.A1(n_2683),
.A2(n_1056),
.B1(n_1045),
.B2(n_13),
.Y(n_2941)
);

BUFx4f_ASAP7_75t_SL g2942 ( 
.A(n_2524),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2546),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2547),
.Y(n_2944)
);

CKINVDCx5p33_ASAP7_75t_R g2945 ( 
.A(n_2743),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2547),
.Y(n_2946)
);

INVx1_ASAP7_75t_SL g2947 ( 
.A(n_2624),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2611),
.Y(n_2948)
);

OAI22xp33_ASAP7_75t_L g2949 ( 
.A1(n_2563),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_2949)
);

INVx2_ASAP7_75t_SL g2950 ( 
.A(n_2701),
.Y(n_2950)
);

AOI22xp33_ASAP7_75t_L g2951 ( 
.A1(n_2759),
.A2(n_1056),
.B1(n_18),
.B2(n_15),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2611),
.Y(n_2952)
);

BUFx12f_ASAP7_75t_L g2953 ( 
.A(n_2600),
.Y(n_2953)
);

OAI22xp33_ASAP7_75t_L g2954 ( 
.A1(n_2563),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2602),
.Y(n_2955)
);

INVx2_ASAP7_75t_SL g2956 ( 
.A(n_2701),
.Y(n_2956)
);

OAI22xp5_ASAP7_75t_SL g2957 ( 
.A1(n_2597),
.A2(n_21),
.B1(n_17),
.B2(n_19),
.Y(n_2957)
);

OAI21xp33_ASAP7_75t_SL g2958 ( 
.A1(n_2559),
.A2(n_21),
.B(n_22),
.Y(n_2958)
);

INVx4_ASAP7_75t_L g2959 ( 
.A(n_2674),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2602),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2741),
.Y(n_2961)
);

OAI22xp33_ASAP7_75t_L g2962 ( 
.A1(n_2563),
.A2(n_26),
.B1(n_22),
.B2(n_25),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2710),
.B(n_25),
.Y(n_2963)
);

AOI22xp33_ASAP7_75t_L g2964 ( 
.A1(n_2759),
.A2(n_1056),
.B1(n_29),
.B2(n_26),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2608),
.Y(n_2965)
);

INVx6_ASAP7_75t_L g2966 ( 
.A(n_2653),
.Y(n_2966)
);

BUFx8_ASAP7_75t_L g2967 ( 
.A(n_2574),
.Y(n_2967)
);

OAI22x1_ASAP7_75t_L g2968 ( 
.A1(n_2513),
.A2(n_32),
.B1(n_28),
.B2(n_30),
.Y(n_2968)
);

OAI22xp33_ASAP7_75t_L g2969 ( 
.A1(n_2563),
.A2(n_34),
.B1(n_28),
.B2(n_33),
.Y(n_2969)
);

CKINVDCx6p67_ASAP7_75t_R g2970 ( 
.A(n_2597),
.Y(n_2970)
);

OAI21xp5_ASAP7_75t_L g2971 ( 
.A1(n_2537),
.A2(n_2541),
.B(n_2531),
.Y(n_2971)
);

BUFx5_ASAP7_75t_L g2972 ( 
.A(n_2516),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2711),
.Y(n_2973)
);

AOI22xp33_ASAP7_75t_SL g2974 ( 
.A1(n_2652),
.A2(n_36),
.B1(n_33),
.B2(n_35),
.Y(n_2974)
);

BUFx2_ASAP7_75t_L g2975 ( 
.A(n_2601),
.Y(n_2975)
);

INVxp67_ASAP7_75t_L g2976 ( 
.A(n_2660),
.Y(n_2976)
);

OAI22xp33_ASAP7_75t_L g2977 ( 
.A1(n_2681),
.A2(n_39),
.B1(n_36),
.B2(n_37),
.Y(n_2977)
);

AOI22xp33_ASAP7_75t_L g2978 ( 
.A1(n_2574),
.A2(n_40),
.B1(n_37),
.B2(n_39),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2711),
.Y(n_2979)
);

INVx4_ASAP7_75t_SL g2980 ( 
.A(n_2674),
.Y(n_2980)
);

BUFx3_ASAP7_75t_L g2981 ( 
.A(n_2624),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2608),
.Y(n_2982)
);

BUFx10_ASAP7_75t_L g2983 ( 
.A(n_2766),
.Y(n_2983)
);

INVx6_ASAP7_75t_L g2984 ( 
.A(n_2653),
.Y(n_2984)
);

CKINVDCx5p33_ASAP7_75t_R g2985 ( 
.A(n_2624),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2672),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2696),
.Y(n_2987)
);

AOI22xp33_ASAP7_75t_L g2988 ( 
.A1(n_2658),
.A2(n_2671),
.B1(n_2666),
.B2(n_2724),
.Y(n_2988)
);

AOI21xp5_ASAP7_75t_L g2989 ( 
.A1(n_2557),
.A2(n_1262),
.B(n_1239),
.Y(n_2989)
);

NAND2x1p5_ASAP7_75t_L g2990 ( 
.A(n_2653),
.B(n_1239),
.Y(n_2990)
);

AOI22xp33_ASAP7_75t_SL g2991 ( 
.A1(n_2652),
.A2(n_2538),
.B1(n_2555),
.B2(n_2539),
.Y(n_2991)
);

CKINVDCx5p33_ASAP7_75t_R g2992 ( 
.A(n_2624),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2699),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2744),
.Y(n_2994)
);

INVx3_ASAP7_75t_L g2995 ( 
.A(n_2729),
.Y(n_2995)
);

OAI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_2655),
.A2(n_1273),
.B1(n_1274),
.B2(n_1262),
.Y(n_2996)
);

OAI22xp33_ASAP7_75t_L g2997 ( 
.A1(n_2681),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_2997)
);

BUFx12f_ASAP7_75t_L g2998 ( 
.A(n_2766),
.Y(n_2998)
);

AOI22xp33_ASAP7_75t_L g2999 ( 
.A1(n_2724),
.A2(n_2735),
.B1(n_2721),
.B2(n_2639),
.Y(n_2999)
);

AOI22xp33_ASAP7_75t_L g3000 ( 
.A1(n_2658),
.A2(n_976),
.B1(n_988),
.B2(n_973),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2874),
.B(n_2878),
.Y(n_3001)
);

AND2x2_ASAP7_75t_L g3002 ( 
.A(n_2930),
.B(n_2613),
.Y(n_3002)
);

OR2x2_ASAP7_75t_L g3003 ( 
.A(n_2879),
.B(n_2710),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2793),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2798),
.Y(n_3005)
);

A2O1A1Ixp33_ASAP7_75t_L g3006 ( 
.A1(n_2796),
.A2(n_2537),
.B(n_2636),
.C(n_2597),
.Y(n_3006)
);

OA21x2_ASAP7_75t_L g3007 ( 
.A1(n_2890),
.A2(n_2521),
.B(n_2708),
.Y(n_3007)
);

NAND2x1_ASAP7_75t_L g3008 ( 
.A(n_2776),
.B(n_2674),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2886),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2774),
.Y(n_3010)
);

AOI22xp33_ASAP7_75t_L g3011 ( 
.A1(n_2779),
.A2(n_2618),
.B1(n_2616),
.B2(n_2724),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2961),
.Y(n_3012)
);

AO31x2_ASAP7_75t_L g3013 ( 
.A1(n_2989),
.A2(n_2559),
.A3(n_2628),
.B(n_2509),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2783),
.Y(n_3014)
);

AND2x4_ASAP7_75t_L g3015 ( 
.A(n_2853),
.B(n_2934),
.Y(n_3015)
);

OA21x2_ASAP7_75t_L g3016 ( 
.A1(n_2923),
.A2(n_2521),
.B(n_2708),
.Y(n_3016)
);

AOI21xp5_ASAP7_75t_L g3017 ( 
.A1(n_2838),
.A2(n_2557),
.B(n_2614),
.Y(n_3017)
);

AOI21xp33_ASAP7_75t_L g3018 ( 
.A1(n_2949),
.A2(n_2735),
.B(n_2687),
.Y(n_3018)
);

NOR2xp33_ASAP7_75t_L g3019 ( 
.A(n_2828),
.B(n_2508),
.Y(n_3019)
);

CKINVDCx20_ASAP7_75t_R g3020 ( 
.A(n_2849),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2784),
.Y(n_3021)
);

BUFx2_ASAP7_75t_L g3022 ( 
.A(n_2889),
.Y(n_3022)
);

OR2x2_ASAP7_75t_L g3023 ( 
.A(n_2891),
.B(n_2710),
.Y(n_3023)
);

INVx3_ASAP7_75t_L g3024 ( 
.A(n_2894),
.Y(n_3024)
);

A2O1A1Ixp33_ASAP7_75t_L g3025 ( 
.A1(n_2796),
.A2(n_2636),
.B(n_2678),
.C(n_2669),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2788),
.Y(n_3026)
);

AO21x2_ASAP7_75t_L g3027 ( 
.A1(n_2989),
.A2(n_2532),
.B(n_2515),
.Y(n_3027)
);

AOI21xp5_ASAP7_75t_L g3028 ( 
.A1(n_2838),
.A2(n_2921),
.B(n_2557),
.Y(n_3028)
);

AOI21xp5_ASAP7_75t_L g3029 ( 
.A1(n_2921),
.A2(n_2614),
.B(n_2555),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2807),
.Y(n_3030)
);

AOI21xp33_ASAP7_75t_L g3031 ( 
.A1(n_2949),
.A2(n_2735),
.B(n_2538),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2976),
.B(n_2710),
.Y(n_3032)
);

AND2x2_ASAP7_75t_L g3033 ( 
.A(n_2975),
.B(n_2616),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2773),
.Y(n_3034)
);

OR2x2_ASAP7_75t_L g3035 ( 
.A(n_2895),
.B(n_2658),
.Y(n_3035)
);

BUFx6f_ASAP7_75t_L g3036 ( 
.A(n_2913),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2790),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_SL g3038 ( 
.A(n_2815),
.B(n_2971),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2811),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2933),
.Y(n_3040)
);

AOI21xp5_ASAP7_75t_L g3041 ( 
.A1(n_2903),
.A2(n_2614),
.B(n_2555),
.Y(n_3041)
);

CKINVDCx11_ASAP7_75t_R g3042 ( 
.A(n_2827),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2976),
.B(n_2748),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2943),
.Y(n_3044)
);

OA21x2_ASAP7_75t_L g3045 ( 
.A1(n_2837),
.A2(n_2512),
.B(n_2606),
.Y(n_3045)
);

OAI21x1_ASAP7_75t_L g3046 ( 
.A1(n_2903),
.A2(n_2512),
.B(n_2532),
.Y(n_3046)
);

NOR2xp33_ASAP7_75t_L g3047 ( 
.A(n_2828),
.B(n_2859),
.Y(n_3047)
);

A2O1A1Ixp33_ASAP7_75t_L g3048 ( 
.A1(n_2785),
.A2(n_2636),
.B(n_2678),
.C(n_2669),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2944),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2986),
.B(n_2748),
.Y(n_3050)
);

OAI21xp5_ASAP7_75t_L g3051 ( 
.A1(n_2771),
.A2(n_2538),
.B(n_2539),
.Y(n_3051)
);

AOI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_2870),
.A2(n_2555),
.B(n_2539),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2987),
.B(n_2748),
.Y(n_3053)
);

AOI21xp5_ASAP7_75t_L g3054 ( 
.A1(n_2870),
.A2(n_2539),
.B(n_2538),
.Y(n_3054)
);

OAI21x1_ASAP7_75t_L g3055 ( 
.A1(n_2937),
.A2(n_2676),
.B(n_2535),
.Y(n_3055)
);

BUFx3_ASAP7_75t_L g3056 ( 
.A(n_2845),
.Y(n_3056)
);

CKINVDCx11_ASAP7_75t_R g3057 ( 
.A(n_2825),
.Y(n_3057)
);

AOI21xp5_ASAP7_75t_L g3058 ( 
.A1(n_2771),
.A2(n_2697),
.B(n_2670),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2946),
.Y(n_3059)
);

OA21x2_ASAP7_75t_L g3060 ( 
.A1(n_2877),
.A2(n_2606),
.B(n_2726),
.Y(n_3060)
);

INVx4_ASAP7_75t_SL g3061 ( 
.A(n_2881),
.Y(n_3061)
);

AND2x4_ASAP7_75t_L g3062 ( 
.A(n_2889),
.B(n_2666),
.Y(n_3062)
);

AND2x4_ASAP7_75t_L g3063 ( 
.A(n_2799),
.B(n_2666),
.Y(n_3063)
);

NOR2x1_ASAP7_75t_SL g3064 ( 
.A(n_2822),
.B(n_2522),
.Y(n_3064)
);

BUFx2_ASAP7_75t_L g3065 ( 
.A(n_2808),
.Y(n_3065)
);

OR2x2_ASAP7_75t_L g3066 ( 
.A(n_2993),
.B(n_2666),
.Y(n_3066)
);

AND2x4_ASAP7_75t_L g3067 ( 
.A(n_2799),
.B(n_2671),
.Y(n_3067)
);

A2O1A1Ixp33_ASAP7_75t_L g3068 ( 
.A1(n_2857),
.A2(n_2678),
.B(n_2695),
.C(n_2669),
.Y(n_3068)
);

BUFx8_ASAP7_75t_L g3069 ( 
.A(n_2847),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2994),
.B(n_2750),
.Y(n_3070)
);

AOI21xp5_ASAP7_75t_L g3071 ( 
.A1(n_2991),
.A2(n_2697),
.B(n_2670),
.Y(n_3071)
);

AOI221xp5_ASAP7_75t_L g3072 ( 
.A1(n_2977),
.A2(n_2607),
.B1(n_2634),
.B2(n_2542),
.C(n_2704),
.Y(n_3072)
);

A2O1A1Ixp33_ASAP7_75t_L g3073 ( 
.A1(n_2867),
.A2(n_2695),
.B(n_2663),
.C(n_2766),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_2809),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2818),
.B(n_2820),
.Y(n_3075)
);

INVx3_ASAP7_75t_L g3076 ( 
.A(n_2894),
.Y(n_3076)
);

OAI21x1_ASAP7_75t_L g3077 ( 
.A1(n_2988),
.A2(n_2676),
.B(n_2535),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2823),
.Y(n_3078)
);

HB1xp67_ASAP7_75t_L g3079 ( 
.A(n_2868),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2814),
.Y(n_3080)
);

OR2x6_ASAP7_75t_L g3081 ( 
.A(n_2940),
.B(n_2671),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2872),
.B(n_2750),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2830),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2816),
.Y(n_3084)
);

OAI21xp5_ASAP7_75t_L g3085 ( 
.A1(n_2941),
.A2(n_2697),
.B(n_2561),
.Y(n_3085)
);

AOI21xp5_ASAP7_75t_L g3086 ( 
.A1(n_2991),
.A2(n_2697),
.B(n_2670),
.Y(n_3086)
);

OAI22xp33_ASAP7_75t_L g3087 ( 
.A1(n_2781),
.A2(n_2681),
.B1(n_2659),
.B2(n_2677),
.Y(n_3087)
);

OAI221xp5_ASAP7_75t_SL g3088 ( 
.A1(n_2978),
.A2(n_2770),
.B1(n_2778),
.B2(n_2997),
.C(n_2977),
.Y(n_3088)
);

BUFx2_ASAP7_75t_L g3089 ( 
.A(n_2883),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2877),
.B(n_2750),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2817),
.Y(n_3091)
);

AOI22xp33_ASAP7_75t_L g3092 ( 
.A1(n_2772),
.A2(n_2618),
.B1(n_2616),
.B2(n_2671),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2833),
.Y(n_3093)
);

OAI21x1_ASAP7_75t_L g3094 ( 
.A1(n_2909),
.A2(n_2768),
.B(n_2572),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2819),
.Y(n_3095)
);

BUFx2_ASAP7_75t_L g3096 ( 
.A(n_2894),
.Y(n_3096)
);

OA21x2_ASAP7_75t_L g3097 ( 
.A1(n_2999),
.A2(n_2755),
.B(n_2726),
.Y(n_3097)
);

AO31x2_ASAP7_75t_L g3098 ( 
.A1(n_2850),
.A2(n_2559),
.A3(n_2509),
.B(n_2549),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2844),
.Y(n_3099)
);

HB1xp67_ASAP7_75t_L g3100 ( 
.A(n_2813),
.Y(n_3100)
);

AND2x2_ASAP7_75t_L g3101 ( 
.A(n_2831),
.B(n_2616),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_L g3102 ( 
.A(n_2839),
.B(n_2939),
.Y(n_3102)
);

OAI221xp5_ASAP7_75t_L g3103 ( 
.A1(n_2941),
.A2(n_2721),
.B1(n_2639),
.B2(n_2695),
.C(n_2542),
.Y(n_3103)
);

INVx2_ASAP7_75t_SL g3104 ( 
.A(n_2945),
.Y(n_3104)
);

OA21x2_ASAP7_75t_L g3105 ( 
.A1(n_2999),
.A2(n_2761),
.B(n_2755),
.Y(n_3105)
);

BUFx3_ASAP7_75t_L g3106 ( 
.A(n_2927),
.Y(n_3106)
);

AOI22xp33_ASAP7_75t_L g3107 ( 
.A1(n_2781),
.A2(n_2618),
.B1(n_2731),
.B2(n_2601),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2863),
.B(n_2603),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2835),
.Y(n_3109)
);

INVx2_ASAP7_75t_SL g3110 ( 
.A(n_2780),
.Y(n_3110)
);

OA21x2_ASAP7_75t_L g3111 ( 
.A1(n_2963),
.A2(n_2761),
.B(n_2572),
.Y(n_3111)
);

OAI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_2887),
.A2(n_2803),
.B(n_2778),
.Y(n_3112)
);

OA21x2_ASAP7_75t_L g3113 ( 
.A1(n_2884),
.A2(n_2720),
.B(n_2713),
.Y(n_3113)
);

BUFx2_ASAP7_75t_L g3114 ( 
.A(n_2812),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_2856),
.Y(n_3115)
);

AOI22xp33_ASAP7_75t_SL g3116 ( 
.A1(n_2957),
.A2(n_2718),
.B1(n_2690),
.B2(n_2522),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_L g3117 ( 
.A(n_2864),
.B(n_2603),
.Y(n_3117)
);

OAI21x1_ASAP7_75t_L g3118 ( 
.A1(n_2990),
.A2(n_2768),
.B(n_2720),
.Y(n_3118)
);

OR2x2_ASAP7_75t_L g3119 ( 
.A(n_2898),
.B(n_2618),
.Y(n_3119)
);

AOI22xp33_ASAP7_75t_L g3120 ( 
.A1(n_2794),
.A2(n_2731),
.B1(n_2528),
.B2(n_2681),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2840),
.Y(n_3121)
);

NAND3xp33_ASAP7_75t_L g3122 ( 
.A(n_2914),
.B(n_2729),
.C(n_2714),
.Y(n_3122)
);

A2O1A1Ixp33_ASAP7_75t_L g3123 ( 
.A1(n_2801),
.A2(n_2731),
.B(n_2681),
.C(n_2659),
.Y(n_3123)
);

BUFx3_ASAP7_75t_L g3124 ( 
.A(n_2802),
.Y(n_3124)
);

BUFx10_ASAP7_75t_L g3125 ( 
.A(n_2804),
.Y(n_3125)
);

INVx2_ASAP7_75t_SL g3126 ( 
.A(n_2780),
.Y(n_3126)
);

A2O1A1Ixp33_ASAP7_75t_L g3127 ( 
.A1(n_2770),
.A2(n_2731),
.B(n_2681),
.C(n_2659),
.Y(n_3127)
);

INVx2_ASAP7_75t_L g3128 ( 
.A(n_2821),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2871),
.B(n_2603),
.Y(n_3129)
);

OA21x2_ASAP7_75t_L g3130 ( 
.A1(n_2843),
.A2(n_2725),
.B(n_2713),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_L g3131 ( 
.A(n_2948),
.B(n_2952),
.Y(n_3131)
);

INVxp67_ASAP7_75t_L g3132 ( 
.A(n_2925),
.Y(n_3132)
);

AOI22xp33_ASAP7_75t_L g3133 ( 
.A1(n_2794),
.A2(n_2528),
.B1(n_2677),
.B2(n_2659),
.Y(n_3133)
);

AOI22xp33_ASAP7_75t_L g3134 ( 
.A1(n_2997),
.A2(n_2528),
.B1(n_2692),
.B2(n_2677),
.Y(n_3134)
);

OAI21x1_ASAP7_75t_L g3135 ( 
.A1(n_2990),
.A2(n_2725),
.B(n_2570),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2955),
.B(n_2664),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2960),
.Y(n_3137)
);

CKINVDCx11_ASAP7_75t_R g3138 ( 
.A(n_2842),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2965),
.Y(n_3139)
);

OAI21xp5_ASAP7_75t_SL g3140 ( 
.A1(n_2978),
.A2(n_2692),
.B(n_2677),
.Y(n_3140)
);

OR2x6_ASAP7_75t_L g3141 ( 
.A(n_2966),
.B(n_2559),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2982),
.B(n_2664),
.Y(n_3142)
);

INVx3_ASAP7_75t_L g3143 ( 
.A(n_2812),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2899),
.Y(n_3144)
);

BUFx3_ASAP7_75t_L g3145 ( 
.A(n_2787),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2829),
.Y(n_3146)
);

AND2x4_ASAP7_75t_L g3147 ( 
.A(n_2799),
.B(n_2509),
.Y(n_3147)
);

AO31x2_ASAP7_75t_L g3148 ( 
.A1(n_2912),
.A2(n_2549),
.A3(n_2558),
.B(n_2533),
.Y(n_3148)
);

OAI21x1_ASAP7_75t_L g3149 ( 
.A1(n_2901),
.A2(n_2570),
.B(n_2567),
.Y(n_3149)
);

BUFx3_ASAP7_75t_L g3150 ( 
.A(n_2873),
.Y(n_3150)
);

AO21x2_ASAP7_75t_L g3151 ( 
.A1(n_2954),
.A2(n_2515),
.B(n_2680),
.Y(n_3151)
);

OAI22x1_ASAP7_75t_L g3152 ( 
.A1(n_2885),
.A2(n_2729),
.B1(n_2717),
.B2(n_2722),
.Y(n_3152)
);

AOI21x1_ASAP7_75t_L g3153 ( 
.A1(n_2907),
.A2(n_2722),
.B(n_2717),
.Y(n_3153)
);

AND2x2_ASAP7_75t_L g3154 ( 
.A(n_2795),
.B(n_2581),
.Y(n_3154)
);

OAI21x1_ASAP7_75t_L g3155 ( 
.A1(n_2901),
.A2(n_2567),
.B(n_2562),
.Y(n_3155)
);

OR2x2_ASAP7_75t_L g3156 ( 
.A(n_2900),
.B(n_2516),
.Y(n_3156)
);

OAI322xp33_ASAP7_75t_L g3157 ( 
.A1(n_2954),
.A2(n_2714),
.A3(n_2728),
.B1(n_2727),
.B2(n_2709),
.C1(n_2527),
.C2(n_2520),
.Y(n_3157)
);

OA21x2_ASAP7_75t_L g3158 ( 
.A1(n_2902),
.A2(n_2592),
.B(n_2590),
.Y(n_3158)
);

AOI21xp5_ASAP7_75t_L g3159 ( 
.A1(n_2815),
.A2(n_2653),
.B(n_2685),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_2841),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2916),
.Y(n_3161)
);

AOI21xp5_ASAP7_75t_L g3162 ( 
.A1(n_2791),
.A2(n_2653),
.B(n_2685),
.Y(n_3162)
);

BUFx2_ASAP7_75t_L g3163 ( 
.A(n_2892),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_L g3164 ( 
.A(n_2917),
.B(n_2664),
.Y(n_3164)
);

INVx2_ASAP7_75t_L g3165 ( 
.A(n_2973),
.Y(n_3165)
);

AOI21xp5_ASAP7_75t_L g3166 ( 
.A1(n_2791),
.A2(n_2653),
.B(n_2685),
.Y(n_3166)
);

BUFx4f_ASAP7_75t_SL g3167 ( 
.A(n_2826),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_2979),
.Y(n_3168)
);

AOI22xp33_ASAP7_75t_SL g3169 ( 
.A1(n_2789),
.A2(n_2718),
.B1(n_2690),
.B2(n_2522),
.Y(n_3169)
);

AOI21xp5_ASAP7_75t_L g3170 ( 
.A1(n_2962),
.A2(n_2506),
.B(n_2690),
.Y(n_3170)
);

AOI21xp5_ASAP7_75t_L g3171 ( 
.A1(n_2962),
.A2(n_2506),
.B(n_2718),
.Y(n_3171)
);

OA21x2_ASAP7_75t_L g3172 ( 
.A1(n_2918),
.A2(n_2592),
.B(n_2590),
.Y(n_3172)
);

AOI21xp5_ASAP7_75t_L g3173 ( 
.A1(n_2969),
.A2(n_2506),
.B(n_2712),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2919),
.B(n_2693),
.Y(n_3174)
);

INVxp67_ASAP7_75t_L g3175 ( 
.A(n_2836),
.Y(n_3175)
);

AOI21xp5_ASAP7_75t_L g3176 ( 
.A1(n_2969),
.A2(n_2915),
.B(n_2914),
.Y(n_3176)
);

AOI22xp33_ASAP7_75t_SL g3177 ( 
.A1(n_2967),
.A2(n_2806),
.B1(n_2792),
.B2(n_2893),
.Y(n_3177)
);

CKINVDCx14_ASAP7_75t_R g3178 ( 
.A(n_2911),
.Y(n_3178)
);

OAI21x1_ASAP7_75t_L g3179 ( 
.A1(n_2995),
.A2(n_2562),
.B(n_2554),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_2852),
.B(n_2896),
.Y(n_3180)
);

AND2x4_ASAP7_75t_L g3181 ( 
.A(n_2799),
.B(n_2520),
.Y(n_3181)
);

OAI22xp5_ASAP7_75t_L g3182 ( 
.A1(n_2915),
.A2(n_2561),
.B1(n_2742),
.B2(n_2692),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_2929),
.B(n_2693),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2972),
.Y(n_3184)
);

OR2x6_ASAP7_75t_L g3185 ( 
.A(n_2966),
.B(n_2677),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2972),
.Y(n_3186)
);

OAI21x1_ASAP7_75t_L g3187 ( 
.A1(n_2995),
.A2(n_2554),
.B(n_2594),
.Y(n_3187)
);

AOI22xp5_ASAP7_75t_L g3188 ( 
.A1(n_2832),
.A2(n_2692),
.B1(n_2566),
.B2(n_2588),
.Y(n_3188)
);

OR2x2_ASAP7_75t_L g3189 ( 
.A(n_2805),
.B(n_2527),
.Y(n_3189)
);

OAI221xp5_ASAP7_75t_L g3190 ( 
.A1(n_2803),
.A2(n_2588),
.B1(n_2604),
.B2(n_2584),
.C(n_2566),
.Y(n_3190)
);

AOI21x1_ASAP7_75t_L g3191 ( 
.A1(n_2968),
.A2(n_2583),
.B(n_2514),
.Y(n_3191)
);

AND2x4_ASAP7_75t_L g3192 ( 
.A(n_2980),
.B(n_2581),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2972),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2972),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2972),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_SL g3196 ( 
.A(n_2800),
.B(n_2692),
.Y(n_3196)
);

BUFx2_ASAP7_75t_L g3197 ( 
.A(n_2782),
.Y(n_3197)
);

OAI21x1_ASAP7_75t_L g3198 ( 
.A1(n_2996),
.A2(n_2599),
.B(n_2594),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_3010),
.Y(n_3199)
);

AND2x2_ASAP7_75t_L g3200 ( 
.A(n_3015),
.B(n_2782),
.Y(n_3200)
);

AOI22xp33_ASAP7_75t_L g3201 ( 
.A1(n_3112),
.A2(n_2967),
.B1(n_2777),
.B2(n_2953),
.Y(n_3201)
);

OAI22xp33_ASAP7_75t_L g3202 ( 
.A1(n_3176),
.A2(n_2942),
.B1(n_2782),
.B2(n_2998),
.Y(n_3202)
);

OR2x6_ASAP7_75t_L g3203 ( 
.A(n_3159),
.B(n_2966),
.Y(n_3203)
);

OAI211xp5_ASAP7_75t_SL g3204 ( 
.A1(n_3038),
.A2(n_2875),
.B(n_2880),
.C(n_2882),
.Y(n_3204)
);

AOI222xp33_ASAP7_75t_L g3205 ( 
.A1(n_3112),
.A2(n_3072),
.B1(n_3103),
.B2(n_3140),
.C1(n_2951),
.C2(n_2964),
.Y(n_3205)
);

OAI21x1_ASAP7_75t_L g3206 ( 
.A1(n_3153),
.A2(n_2647),
.B(n_2640),
.Y(n_3206)
);

INVx3_ASAP7_75t_L g3207 ( 
.A(n_3015),
.Y(n_3207)
);

OAI21xp33_ASAP7_75t_L g3208 ( 
.A1(n_3088),
.A2(n_2964),
.B(n_2951),
.Y(n_3208)
);

AOI221xp5_ASAP7_75t_L g3209 ( 
.A1(n_3088),
.A2(n_3176),
.B1(n_3018),
.B2(n_3103),
.C(n_3006),
.Y(n_3209)
);

NOR2x1p5_ASAP7_75t_L g3210 ( 
.A(n_3106),
.B(n_2862),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_3001),
.B(n_2972),
.Y(n_3211)
);

OR2x2_ASAP7_75t_L g3212 ( 
.A(n_3032),
.B(n_2786),
.Y(n_3212)
);

HB1xp67_ASAP7_75t_L g3213 ( 
.A(n_3079),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3014),
.Y(n_3214)
);

OAI22xp33_ASAP7_75t_L g3215 ( 
.A1(n_3190),
.A2(n_2942),
.B1(n_2959),
.B2(n_2881),
.Y(n_3215)
);

AOI21xp5_ASAP7_75t_L g3216 ( 
.A1(n_3028),
.A2(n_2861),
.B(n_2858),
.Y(n_3216)
);

AND2x4_ASAP7_75t_L g3217 ( 
.A(n_3141),
.B(n_2980),
.Y(n_3217)
);

OR2x2_ASAP7_75t_L g3218 ( 
.A(n_3032),
.B(n_2947),
.Y(n_3218)
);

INVx11_ASAP7_75t_L g3219 ( 
.A(n_3069),
.Y(n_3219)
);

OAI22xp5_ASAP7_75t_L g3220 ( 
.A1(n_3116),
.A2(n_2974),
.B1(n_2938),
.B2(n_2858),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3021),
.Y(n_3221)
);

AOI22xp33_ASAP7_75t_SL g3222 ( 
.A1(n_3182),
.A2(n_2958),
.B1(n_2780),
.B2(n_2810),
.Y(n_3222)
);

CKINVDCx5p33_ASAP7_75t_R g3223 ( 
.A(n_3057),
.Y(n_3223)
);

OAI221xp5_ASAP7_75t_L g3224 ( 
.A1(n_3177),
.A2(n_2861),
.B1(n_2848),
.B2(n_2880),
.C(n_2875),
.Y(n_3224)
);

OAI22xp33_ASAP7_75t_L g3225 ( 
.A1(n_3190),
.A2(n_2959),
.B1(n_2970),
.B2(n_2912),
.Y(n_3225)
);

AND2x4_ASAP7_75t_L g3226 ( 
.A(n_3141),
.B(n_3062),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3026),
.Y(n_3227)
);

AOI221xp5_ASAP7_75t_L g3228 ( 
.A1(n_3018),
.A2(n_2904),
.B1(n_2974),
.B2(n_2938),
.C(n_2846),
.Y(n_3228)
);

OAI22xp33_ASAP7_75t_L g3229 ( 
.A1(n_3122),
.A2(n_2910),
.B1(n_2905),
.B2(n_2984),
.Y(n_3229)
);

OAI21x1_ASAP7_75t_L g3230 ( 
.A1(n_3159),
.A2(n_2647),
.B(n_2640),
.Y(n_3230)
);

INVx2_ASAP7_75t_SL g3231 ( 
.A(n_3036),
.Y(n_3231)
);

AOI221xp5_ASAP7_75t_L g3232 ( 
.A1(n_3072),
.A2(n_2897),
.B1(n_2906),
.B2(n_2936),
.C(n_2920),
.Y(n_3232)
);

NAND3xp33_ASAP7_75t_L g3233 ( 
.A(n_3100),
.B(n_2865),
.C(n_2906),
.Y(n_3233)
);

OAI22xp5_ASAP7_75t_L g3234 ( 
.A1(n_3116),
.A2(n_2797),
.B1(n_2865),
.B2(n_2824),
.Y(n_3234)
);

OAI221xp5_ASAP7_75t_L g3235 ( 
.A1(n_3177),
.A2(n_2869),
.B1(n_2834),
.B2(n_2797),
.C(n_2888),
.Y(n_3235)
);

AOI22xp33_ASAP7_75t_L g3236 ( 
.A1(n_3133),
.A2(n_2922),
.B1(n_2855),
.B2(n_2908),
.Y(n_3236)
);

OAI22xp5_ASAP7_75t_L g3237 ( 
.A1(n_3011),
.A2(n_3134),
.B1(n_3169),
.B2(n_3025),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_3001),
.B(n_3090),
.Y(n_3238)
);

BUFx3_ASAP7_75t_L g3239 ( 
.A(n_3020),
.Y(n_3239)
);

AND2x2_ASAP7_75t_L g3240 ( 
.A(n_3065),
.B(n_2928),
.Y(n_3240)
);

AOI222xp33_ASAP7_75t_L g3241 ( 
.A1(n_3019),
.A2(n_2519),
.B1(n_2851),
.B2(n_2860),
.C1(n_2873),
.C2(n_2810),
.Y(n_3241)
);

AOI211xp5_ASAP7_75t_SL g3242 ( 
.A1(n_3087),
.A2(n_2932),
.B(n_2924),
.C(n_2775),
.Y(n_3242)
);

OAI211xp5_ASAP7_75t_L g3243 ( 
.A1(n_3058),
.A2(n_2810),
.B(n_2992),
.C(n_2985),
.Y(n_3243)
);

OA21x2_ASAP7_75t_L g3244 ( 
.A1(n_3184),
.A2(n_2599),
.B(n_2553),
.Y(n_3244)
);

AOI22xp33_ASAP7_75t_L g3245 ( 
.A1(n_3120),
.A2(n_2981),
.B1(n_2528),
.B2(n_2604),
.Y(n_3245)
);

AOI22xp33_ASAP7_75t_L g3246 ( 
.A1(n_3182),
.A2(n_2528),
.B1(n_2584),
.B2(n_2680),
.Y(n_3246)
);

NAND4xp25_ASAP7_75t_L g3247 ( 
.A(n_3092),
.B(n_2727),
.C(n_2728),
.D(n_2709),
.Y(n_3247)
);

AND2x2_ASAP7_75t_L g3248 ( 
.A(n_3089),
.B(n_3002),
.Y(n_3248)
);

AND2x2_ASAP7_75t_L g3249 ( 
.A(n_3033),
.B(n_2980),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_3004),
.Y(n_3250)
);

OAI21x1_ASAP7_75t_L g3251 ( 
.A1(n_3162),
.A2(n_2552),
.B(n_2684),
.Y(n_3251)
);

AND2x2_ASAP7_75t_L g3252 ( 
.A(n_3101),
.B(n_2776),
.Y(n_3252)
);

OAI22xp5_ASAP7_75t_L g3253 ( 
.A1(n_3169),
.A2(n_2742),
.B1(n_2866),
.B2(n_2776),
.Y(n_3253)
);

BUFx6f_ASAP7_75t_L g3254 ( 
.A(n_3036),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_3090),
.B(n_2680),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_3180),
.B(n_2866),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_3030),
.Y(n_3257)
);

HB1xp67_ASAP7_75t_L g3258 ( 
.A(n_3066),
.Y(n_3258)
);

AND2x2_ASAP7_75t_L g3259 ( 
.A(n_3154),
.B(n_2866),
.Y(n_3259)
);

A2O1A1Ixp33_ASAP7_75t_L g3260 ( 
.A1(n_3068),
.A2(n_2854),
.B(n_2775),
.C(n_2931),
.Y(n_3260)
);

AND2x2_ASAP7_75t_L g3261 ( 
.A(n_3163),
.B(n_2876),
.Y(n_3261)
);

CKINVDCx20_ASAP7_75t_R g3262 ( 
.A(n_3042),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_3005),
.Y(n_3263)
);

AOI221xp5_ASAP7_75t_L g3264 ( 
.A1(n_3058),
.A2(n_2956),
.B1(n_2950),
.B2(n_2719),
.C(n_2715),
.Y(n_3264)
);

AND2x2_ASAP7_75t_L g3265 ( 
.A(n_3022),
.B(n_2876),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3039),
.Y(n_3266)
);

BUFx3_ASAP7_75t_L g3267 ( 
.A(n_3036),
.Y(n_3267)
);

AO21x1_ASAP7_75t_L g3268 ( 
.A1(n_3047),
.A2(n_2733),
.B(n_2712),
.Y(n_3268)
);

BUFx3_ASAP7_75t_L g3269 ( 
.A(n_3056),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3040),
.Y(n_3270)
);

AO31x2_ASAP7_75t_L g3271 ( 
.A1(n_3064),
.A2(n_2549),
.A3(n_2558),
.B(n_2533),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3044),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3049),
.Y(n_3273)
);

AOI221xp5_ASAP7_75t_L g3274 ( 
.A1(n_3031),
.A2(n_2719),
.B1(n_2715),
.B2(n_2711),
.C(n_2644),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3128),
.Y(n_3275)
);

OA21x2_ASAP7_75t_L g3276 ( 
.A1(n_3186),
.A2(n_2553),
.B(n_2526),
.Y(n_3276)
);

INVx4_ASAP7_75t_L g3277 ( 
.A(n_3061),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3059),
.Y(n_3278)
);

HB1xp67_ASAP7_75t_L g3279 ( 
.A(n_3119),
.Y(n_3279)
);

AOI21xp5_ASAP7_75t_L g3280 ( 
.A1(n_3028),
.A2(n_2749),
.B(n_2536),
.Y(n_3280)
);

AND2x2_ASAP7_75t_L g3281 ( 
.A(n_3175),
.B(n_2876),
.Y(n_3281)
);

AOI22xp33_ASAP7_75t_SL g3282 ( 
.A1(n_3178),
.A2(n_2984),
.B1(n_2742),
.B2(n_2983),
.Y(n_3282)
);

INVxp67_ASAP7_75t_SL g3283 ( 
.A(n_3075),
.Y(n_3283)
);

INVxp67_ASAP7_75t_L g3284 ( 
.A(n_3102),
.Y(n_3284)
);

AND2x2_ASAP7_75t_L g3285 ( 
.A(n_3062),
.B(n_2935),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3078),
.Y(n_3286)
);

AOI222xp33_ASAP7_75t_L g3287 ( 
.A1(n_3085),
.A2(n_2519),
.B1(n_45),
.B2(n_47),
.C1(n_42),
.C2(n_44),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3083),
.Y(n_3288)
);

AOI22xp33_ASAP7_75t_L g3289 ( 
.A1(n_3107),
.A2(n_2935),
.B1(n_2983),
.B2(n_2769),
.Y(n_3289)
);

AOI22xp5_ASAP7_75t_L g3290 ( 
.A1(n_3188),
.A2(n_2769),
.B1(n_2984),
.B2(n_2739),
.Y(n_3290)
);

AND2x4_ASAP7_75t_L g3291 ( 
.A(n_3141),
.B(n_2533),
.Y(n_3291)
);

OAI22xp33_ASAP7_75t_L g3292 ( 
.A1(n_3081),
.A2(n_2739),
.B1(n_2769),
.B2(n_2561),
.Y(n_3292)
);

INVx2_ASAP7_75t_L g3293 ( 
.A(n_3146),
.Y(n_3293)
);

AOI22xp33_ASAP7_75t_L g3294 ( 
.A1(n_3081),
.A2(n_3085),
.B1(n_3196),
.B2(n_3031),
.Y(n_3294)
);

AND2x4_ASAP7_75t_L g3295 ( 
.A(n_3181),
.B(n_2558),
.Y(n_3295)
);

AOI22xp33_ASAP7_75t_L g3296 ( 
.A1(n_3081),
.A2(n_2769),
.B1(n_2609),
.B2(n_2581),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3093),
.Y(n_3297)
);

OAI211xp5_ASAP7_75t_SL g3298 ( 
.A1(n_3048),
.A2(n_2609),
.B(n_2581),
.C(n_2550),
.Y(n_3298)
);

AOI222xp33_ASAP7_75t_L g3299 ( 
.A1(n_3051),
.A2(n_47),
.B1(n_49),
.B2(n_44),
.C1(n_46),
.C2(n_48),
.Y(n_3299)
);

OAI22xp5_ASAP7_75t_L g3300 ( 
.A1(n_3127),
.A2(n_2742),
.B1(n_2712),
.B2(n_2733),
.Y(n_3300)
);

OAI211xp5_ASAP7_75t_L g3301 ( 
.A1(n_3051),
.A2(n_2612),
.B(n_2644),
.C(n_2630),
.Y(n_3301)
);

AOI22xp33_ASAP7_75t_L g3302 ( 
.A1(n_3150),
.A2(n_3171),
.B1(n_3170),
.B2(n_3110),
.Y(n_3302)
);

OR2x6_ASAP7_75t_L g3303 ( 
.A(n_3162),
.B(n_2568),
.Y(n_3303)
);

AO31x2_ASAP7_75t_L g3304 ( 
.A1(n_3054),
.A2(n_2568),
.A3(n_2719),
.B(n_2715),
.Y(n_3304)
);

BUFx3_ASAP7_75t_L g3305 ( 
.A(n_3124),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3109),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3121),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_3082),
.B(n_2612),
.Y(n_3308)
);

AOI21xp5_ASAP7_75t_L g3309 ( 
.A1(n_3017),
.A2(n_2749),
.B(n_2536),
.Y(n_3309)
);

AOI22xp5_ASAP7_75t_L g3310 ( 
.A1(n_3123),
.A2(n_2739),
.B1(n_2609),
.B2(n_2514),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3043),
.B(n_2568),
.Y(n_3311)
);

AND2x2_ASAP7_75t_L g3312 ( 
.A(n_3096),
.B(n_2609),
.Y(n_3312)
);

AOI22xp33_ASAP7_75t_SL g3313 ( 
.A1(n_3151),
.A2(n_2742),
.B1(n_2739),
.B2(n_2730),
.Y(n_3313)
);

AOI22xp5_ASAP7_75t_L g3314 ( 
.A1(n_3073),
.A2(n_2739),
.B1(n_2514),
.B2(n_2586),
.Y(n_3314)
);

HB1xp67_ASAP7_75t_L g3315 ( 
.A(n_3003),
.Y(n_3315)
);

AOI211xp5_ASAP7_75t_L g3316 ( 
.A1(n_3170),
.A2(n_3171),
.B(n_3166),
.C(n_3173),
.Y(n_3316)
);

OAI221xp5_ASAP7_75t_L g3317 ( 
.A1(n_3132),
.A2(n_2730),
.B1(n_2550),
.B2(n_2510),
.C(n_3000),
.Y(n_3317)
);

BUFx2_ASAP7_75t_L g3318 ( 
.A(n_3114),
.Y(n_3318)
);

HB1xp67_ASAP7_75t_L g3319 ( 
.A(n_3023),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3137),
.Y(n_3320)
);

OAI22xp5_ASAP7_75t_L g3321 ( 
.A1(n_3173),
.A2(n_2745),
.B1(n_2733),
.B2(n_2643),
.Y(n_3321)
);

INVx3_ASAP7_75t_L g3322 ( 
.A(n_3008),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3139),
.Y(n_3323)
);

AOI221xp5_ASAP7_75t_L g3324 ( 
.A1(n_3157),
.A2(n_2662),
.B1(n_2668),
.B2(n_2650),
.C(n_2630),
.Y(n_3324)
);

AOI221xp5_ASAP7_75t_L g3325 ( 
.A1(n_3082),
.A2(n_2668),
.B1(n_2679),
.B2(n_2662),
.C(n_2650),
.Y(n_3325)
);

AOI22xp5_ASAP7_75t_L g3326 ( 
.A1(n_3132),
.A2(n_2739),
.B1(n_2514),
.B2(n_2586),
.Y(n_3326)
);

OAI22xp33_ASAP7_75t_L g3327 ( 
.A1(n_3191),
.A2(n_3166),
.B1(n_3185),
.B2(n_3152),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3043),
.B(n_2679),
.Y(n_3328)
);

AOI22xp33_ASAP7_75t_L g3329 ( 
.A1(n_3126),
.A2(n_2586),
.B1(n_2583),
.B2(n_2730),
.Y(n_3329)
);

AOI22xp33_ASAP7_75t_L g3330 ( 
.A1(n_3151),
.A2(n_2586),
.B1(n_2583),
.B2(n_2536),
.Y(n_3330)
);

AOI22xp33_ASAP7_75t_L g3331 ( 
.A1(n_3138),
.A2(n_2583),
.B1(n_2610),
.B2(n_2749),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_3160),
.Y(n_3332)
);

AO21x2_ASAP7_75t_L g3333 ( 
.A1(n_3193),
.A2(n_2515),
.B(n_2760),
.Y(n_3333)
);

OAI221xp5_ASAP7_75t_L g3334 ( 
.A1(n_3104),
.A2(n_2550),
.B1(n_2510),
.B2(n_2643),
.C(n_2552),
.Y(n_3334)
);

INVx2_ASAP7_75t_L g3335 ( 
.A(n_3165),
.Y(n_3335)
);

INVx3_ASAP7_75t_L g3336 ( 
.A(n_3143),
.Y(n_3336)
);

AOI22xp33_ASAP7_75t_L g3337 ( 
.A1(n_3069),
.A2(n_2610),
.B1(n_2550),
.B2(n_2510),
.Y(n_3337)
);

A2O1A1Ixp33_ASAP7_75t_L g3338 ( 
.A1(n_3071),
.A2(n_2552),
.B(n_2510),
.C(n_2556),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_3144),
.B(n_2693),
.Y(n_3339)
);

AOI22xp33_ASAP7_75t_L g3340 ( 
.A1(n_3145),
.A2(n_2610),
.B1(n_2598),
.B2(n_2760),
.Y(n_3340)
);

OAI22xp5_ASAP7_75t_L g3341 ( 
.A1(n_3071),
.A2(n_2745),
.B1(n_2643),
.B2(n_2682),
.Y(n_3341)
);

OAI22xp5_ASAP7_75t_L g3342 ( 
.A1(n_3086),
.A2(n_2745),
.B1(n_2682),
.B2(n_2926),
.Y(n_3342)
);

AOI222xp33_ASAP7_75t_L g3343 ( 
.A1(n_3167),
.A2(n_53),
.B1(n_55),
.B2(n_46),
.C1(n_52),
.C2(n_54),
.Y(n_3343)
);

AOI221xp5_ASAP7_75t_L g3344 ( 
.A1(n_3086),
.A2(n_2702),
.B1(n_2552),
.B2(n_54),
.C(n_52),
.Y(n_3344)
);

OAI22xp33_ASAP7_75t_L g3345 ( 
.A1(n_3185),
.A2(n_2702),
.B1(n_2760),
.B2(n_2598),
.Y(n_3345)
);

AOI22xp33_ASAP7_75t_SL g3346 ( 
.A1(n_3052),
.A2(n_3054),
.B1(n_3041),
.B2(n_3017),
.Y(n_3346)
);

OAI22xp5_ASAP7_75t_L g3347 ( 
.A1(n_3052),
.A2(n_2702),
.B1(n_56),
.B2(n_53),
.Y(n_3347)
);

NAND3xp33_ASAP7_75t_L g3348 ( 
.A(n_3050),
.B(n_976),
.C(n_973),
.Y(n_3348)
);

AOI221xp5_ASAP7_75t_L g3349 ( 
.A1(n_3050),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.C(n_58),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3131),
.Y(n_3350)
);

CKINVDCx14_ASAP7_75t_R g3351 ( 
.A(n_3125),
.Y(n_3351)
);

AOI321xp33_ASAP7_75t_L g3352 ( 
.A1(n_3041),
.A2(n_61),
.A3(n_63),
.B1(n_57),
.B2(n_60),
.C(n_62),
.Y(n_3352)
);

AOI22xp33_ASAP7_75t_L g3353 ( 
.A1(n_3185),
.A2(n_2598),
.B1(n_2622),
.B2(n_2627),
.Y(n_3353)
);

AND2x2_ASAP7_75t_L g3354 ( 
.A(n_3197),
.B(n_2684),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3161),
.B(n_2686),
.Y(n_3355)
);

OAI22xp5_ASAP7_75t_L g3356 ( 
.A1(n_3029),
.A2(n_65),
.B1(n_62),
.B2(n_64),
.Y(n_3356)
);

OR2x2_ASAP7_75t_L g3357 ( 
.A(n_3053),
.B(n_2686),
.Y(n_3357)
);

AO22x1_ASAP7_75t_L g3358 ( 
.A1(n_3192),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3131),
.Y(n_3359)
);

AOI22xp33_ASAP7_75t_L g3360 ( 
.A1(n_3077),
.A2(n_2622),
.B1(n_2629),
.B2(n_2627),
.Y(n_3360)
);

AOI22xp33_ASAP7_75t_L g3361 ( 
.A1(n_3063),
.A2(n_2629),
.B1(n_2689),
.B2(n_2619),
.Y(n_3361)
);

BUFx2_ASAP7_75t_L g3362 ( 
.A(n_3322),
.Y(n_3362)
);

OR2x2_ASAP7_75t_L g3363 ( 
.A(n_3211),
.B(n_3053),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3207),
.B(n_3063),
.Y(n_3364)
);

AND2x2_ASAP7_75t_L g3365 ( 
.A(n_3207),
.B(n_3226),
.Y(n_3365)
);

INVx2_ASAP7_75t_L g3366 ( 
.A(n_3271),
.Y(n_3366)
);

BUFx2_ASAP7_75t_L g3367 ( 
.A(n_3322),
.Y(n_3367)
);

AND2x2_ASAP7_75t_L g3368 ( 
.A(n_3226),
.B(n_3067),
.Y(n_3368)
);

AND2x4_ASAP7_75t_L g3369 ( 
.A(n_3217),
.B(n_3143),
.Y(n_3369)
);

INVx2_ASAP7_75t_L g3370 ( 
.A(n_3271),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3199),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_3271),
.Y(n_3372)
);

INVx1_ASAP7_75t_SL g3373 ( 
.A(n_3262),
.Y(n_3373)
);

AND2x4_ASAP7_75t_L g3374 ( 
.A(n_3217),
.B(n_3192),
.Y(n_3374)
);

AND2x2_ASAP7_75t_L g3375 ( 
.A(n_3318),
.B(n_3067),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3213),
.B(n_3070),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3214),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_3200),
.B(n_3181),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_3248),
.B(n_3147),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_3350),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_SL g3381 ( 
.A(n_3229),
.B(n_3061),
.Y(n_3381)
);

INVxp67_ASAP7_75t_R g3382 ( 
.A(n_3300),
.Y(n_3382)
);

OAI221xp5_ASAP7_75t_L g3383 ( 
.A1(n_3209),
.A2(n_3070),
.B1(n_3189),
.B2(n_3035),
.C(n_3075),
.Y(n_3383)
);

AND2x2_ASAP7_75t_L g3384 ( 
.A(n_3265),
.B(n_3147),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3359),
.B(n_3009),
.Y(n_3385)
);

AND2x2_ASAP7_75t_L g3386 ( 
.A(n_3261),
.B(n_3195),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3221),
.Y(n_3387)
);

INVx2_ASAP7_75t_L g3388 ( 
.A(n_3227),
.Y(n_3388)
);

AND2x4_ASAP7_75t_L g3389 ( 
.A(n_3203),
.B(n_3098),
.Y(n_3389)
);

INVx2_ASAP7_75t_L g3390 ( 
.A(n_3257),
.Y(n_3390)
);

OAI22xp5_ASAP7_75t_L g3391 ( 
.A1(n_3220),
.A2(n_3024),
.B1(n_3076),
.B2(n_3029),
.Y(n_3391)
);

INVx2_ASAP7_75t_L g3392 ( 
.A(n_3266),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3270),
.Y(n_3393)
);

BUFx6f_ASAP7_75t_SL g3394 ( 
.A(n_3277),
.Y(n_3394)
);

OR2x2_ASAP7_75t_L g3395 ( 
.A(n_3211),
.B(n_3168),
.Y(n_3395)
);

AND2x2_ASAP7_75t_L g3396 ( 
.A(n_3336),
.B(n_3024),
.Y(n_3396)
);

OR2x2_ASAP7_75t_L g3397 ( 
.A(n_3238),
.B(n_3095),
.Y(n_3397)
);

INVx2_ASAP7_75t_L g3398 ( 
.A(n_3272),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3283),
.B(n_3012),
.Y(n_3399)
);

AO21x2_ASAP7_75t_L g3400 ( 
.A1(n_3347),
.A2(n_3194),
.B(n_3046),
.Y(n_3400)
);

INVx5_ASAP7_75t_SL g3401 ( 
.A(n_3219),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3273),
.Y(n_3402)
);

INVxp67_ASAP7_75t_L g3403 ( 
.A(n_3212),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3238),
.B(n_3034),
.Y(n_3404)
);

AND2x4_ASAP7_75t_L g3405 ( 
.A(n_3203),
.B(n_3098),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3278),
.Y(n_3406)
);

HB1xp67_ASAP7_75t_L g3407 ( 
.A(n_3258),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3286),
.Y(n_3408)
);

INVx3_ASAP7_75t_L g3409 ( 
.A(n_3336),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3288),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_SL g3411 ( 
.A(n_3202),
.B(n_3061),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_3297),
.Y(n_3412)
);

AND2x2_ASAP7_75t_L g3413 ( 
.A(n_3256),
.B(n_3281),
.Y(n_3413)
);

INVx2_ASAP7_75t_R g3414 ( 
.A(n_3305),
.Y(n_3414)
);

BUFx4f_ASAP7_75t_L g3415 ( 
.A(n_3254),
.Y(n_3415)
);

AND2x4_ASAP7_75t_L g3416 ( 
.A(n_3203),
.B(n_3098),
.Y(n_3416)
);

NAND3xp33_ASAP7_75t_L g3417 ( 
.A(n_3316),
.B(n_3007),
.C(n_3099),
.Y(n_3417)
);

AND2x2_ASAP7_75t_L g3418 ( 
.A(n_3259),
.B(n_3076),
.Y(n_3418)
);

AND2x4_ASAP7_75t_L g3419 ( 
.A(n_3303),
.B(n_3037),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_3306),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3307),
.Y(n_3421)
);

INVx2_ASAP7_75t_L g3422 ( 
.A(n_3320),
.Y(n_3422)
);

INVx1_ASAP7_75t_SL g3423 ( 
.A(n_3223),
.Y(n_3423)
);

NAND2xp33_ASAP7_75t_SL g3424 ( 
.A(n_3277),
.B(n_3074),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3216),
.B(n_3315),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_3323),
.Y(n_3426)
);

HB1xp67_ASAP7_75t_L g3427 ( 
.A(n_3279),
.Y(n_3427)
);

AOI221xp5_ASAP7_75t_L g3428 ( 
.A1(n_3220),
.A2(n_3091),
.B1(n_3084),
.B2(n_3080),
.C(n_3115),
.Y(n_3428)
);

INVx2_ASAP7_75t_L g3429 ( 
.A(n_3250),
.Y(n_3429)
);

INVx3_ASAP7_75t_L g3430 ( 
.A(n_3295),
.Y(n_3430)
);

INVx3_ASAP7_75t_L g3431 ( 
.A(n_3295),
.Y(n_3431)
);

INVx2_ASAP7_75t_L g3432 ( 
.A(n_3263),
.Y(n_3432)
);

AND2x4_ASAP7_75t_L g3433 ( 
.A(n_3303),
.B(n_3148),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3339),
.Y(n_3434)
);

BUFx6f_ASAP7_75t_L g3435 ( 
.A(n_3254),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3339),
.Y(n_3436)
);

AND2x4_ASAP7_75t_L g3437 ( 
.A(n_3303),
.B(n_3148),
.Y(n_3437)
);

NOR2xp67_ASAP7_75t_L g3438 ( 
.A(n_3243),
.B(n_3164),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_3275),
.Y(n_3439)
);

NAND2x1_ASAP7_75t_L g3440 ( 
.A(n_3253),
.B(n_3007),
.Y(n_3440)
);

INVxp67_ASAP7_75t_L g3441 ( 
.A(n_3311),
.Y(n_3441)
);

BUFx6f_ASAP7_75t_L g3442 ( 
.A(n_3254),
.Y(n_3442)
);

INVx3_ASAP7_75t_L g3443 ( 
.A(n_3291),
.Y(n_3443)
);

INVxp67_ASAP7_75t_SL g3444 ( 
.A(n_3268),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_3311),
.Y(n_3445)
);

NOR2x1_ASAP7_75t_L g3446 ( 
.A(n_3210),
.B(n_3136),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3293),
.Y(n_3447)
);

HB1xp67_ASAP7_75t_L g3448 ( 
.A(n_3319),
.Y(n_3448)
);

AND2x4_ASAP7_75t_SL g3449 ( 
.A(n_3240),
.B(n_3125),
.Y(n_3449)
);

INVx3_ASAP7_75t_L g3450 ( 
.A(n_3291),
.Y(n_3450)
);

AND2x2_ASAP7_75t_L g3451 ( 
.A(n_3252),
.B(n_3148),
.Y(n_3451)
);

NOR2xp33_ASAP7_75t_L g3452 ( 
.A(n_3351),
.B(n_3136),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3355),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3328),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3355),
.Y(n_3455)
);

HB1xp67_ASAP7_75t_L g3456 ( 
.A(n_3332),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3335),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_3285),
.B(n_3045),
.Y(n_3458)
);

HB1xp67_ASAP7_75t_L g3459 ( 
.A(n_3218),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3308),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_3304),
.Y(n_3461)
);

HB1xp67_ASAP7_75t_L g3462 ( 
.A(n_3357),
.Y(n_3462)
);

AND2x2_ASAP7_75t_L g3463 ( 
.A(n_3249),
.B(n_3045),
.Y(n_3463)
);

INVx2_ASAP7_75t_L g3464 ( 
.A(n_3304),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3304),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3255),
.Y(n_3466)
);

BUFx2_ASAP7_75t_L g3467 ( 
.A(n_3267),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3255),
.Y(n_3468)
);

OR2x2_ASAP7_75t_L g3469 ( 
.A(n_3302),
.B(n_3164),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3312),
.Y(n_3470)
);

INVx2_ASAP7_75t_L g3471 ( 
.A(n_3354),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_3333),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3313),
.B(n_3111),
.Y(n_3473)
);

OR2x2_ASAP7_75t_L g3474 ( 
.A(n_3253),
.B(n_3174),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3347),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3333),
.Y(n_3476)
);

AND2x2_ASAP7_75t_L g3477 ( 
.A(n_3294),
.B(n_3111),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3301),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3233),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3325),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3356),
.Y(n_3481)
);

AND2x2_ASAP7_75t_L g3482 ( 
.A(n_3296),
.B(n_3174),
.Y(n_3482)
);

INVx3_ASAP7_75t_L g3483 ( 
.A(n_3231),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_3206),
.Y(n_3484)
);

OR2x2_ASAP7_75t_L g3485 ( 
.A(n_3327),
.B(n_3183),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3251),
.Y(n_3486)
);

OR2x2_ASAP7_75t_L g3487 ( 
.A(n_3341),
.B(n_3183),
.Y(n_3487)
);

AND2x2_ASAP7_75t_L g3488 ( 
.A(n_3284),
.B(n_3108),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3274),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_3264),
.B(n_3234),
.Y(n_3490)
);

AND2x2_ASAP7_75t_L g3491 ( 
.A(n_3282),
.B(n_3108),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_3234),
.B(n_3142),
.Y(n_3492)
);

BUFx2_ASAP7_75t_L g3493 ( 
.A(n_3338),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3356),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3324),
.Y(n_3495)
);

INVx2_ASAP7_75t_L g3496 ( 
.A(n_3366),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3371),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3371),
.Y(n_3498)
);

AND2x2_ASAP7_75t_L g3499 ( 
.A(n_3368),
.B(n_3290),
.Y(n_3499)
);

INVxp67_ASAP7_75t_SL g3500 ( 
.A(n_3461),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_SL g3501 ( 
.A(n_3493),
.B(n_3352),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3368),
.B(n_3289),
.Y(n_3502)
);

OAI22xp5_ASAP7_75t_L g3503 ( 
.A1(n_3490),
.A2(n_3237),
.B1(n_3222),
.B2(n_3201),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3480),
.B(n_3237),
.Y(n_3504)
);

AOI22xp33_ASAP7_75t_L g3505 ( 
.A1(n_3479),
.A2(n_3208),
.B1(n_3205),
.B2(n_3204),
.Y(n_3505)
);

OAI22xp5_ASAP7_75t_L g3506 ( 
.A1(n_3493),
.A2(n_3224),
.B1(n_3344),
.B2(n_3314),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3374),
.B(n_3241),
.Y(n_3507)
);

INVx2_ASAP7_75t_L g3508 ( 
.A(n_3366),
.Y(n_3508)
);

AOI22xp33_ASAP7_75t_SL g3509 ( 
.A1(n_3391),
.A2(n_3235),
.B1(n_3287),
.B2(n_3205),
.Y(n_3509)
);

AOI22xp33_ASAP7_75t_L g3510 ( 
.A1(n_3495),
.A2(n_3287),
.B1(n_3228),
.B2(n_3299),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3387),
.Y(n_3511)
);

AND2x4_ASAP7_75t_L g3512 ( 
.A(n_3446),
.B(n_3260),
.Y(n_3512)
);

BUFx6f_ASAP7_75t_L g3513 ( 
.A(n_3435),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3387),
.Y(n_3514)
);

AOI21xp33_ASAP7_75t_L g3515 ( 
.A1(n_3489),
.A2(n_3299),
.B(n_3343),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_3495),
.B(n_3232),
.Y(n_3516)
);

BUFx2_ASAP7_75t_L g3517 ( 
.A(n_3467),
.Y(n_3517)
);

OAI21x1_ASAP7_75t_L g3518 ( 
.A1(n_3440),
.A2(n_3409),
.B(n_3486),
.Y(n_3518)
);

OA21x2_ASAP7_75t_L g3519 ( 
.A1(n_3417),
.A2(n_3309),
.B(n_3280),
.Y(n_3519)
);

INVx2_ASAP7_75t_SL g3520 ( 
.A(n_3449),
.Y(n_3520)
);

AO21x2_ASAP7_75t_L g3521 ( 
.A1(n_3444),
.A2(n_3225),
.B(n_3215),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3370),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3393),
.Y(n_3523)
);

INVx4_ASAP7_75t_L g3524 ( 
.A(n_3435),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3393),
.Y(n_3525)
);

HB1xp67_ASAP7_75t_L g3526 ( 
.A(n_3407),
.Y(n_3526)
);

AO31x2_ASAP7_75t_L g3527 ( 
.A1(n_3489),
.A2(n_3341),
.A3(n_3321),
.B(n_3342),
.Y(n_3527)
);

HB1xp67_ASAP7_75t_L g3528 ( 
.A(n_3427),
.Y(n_3528)
);

OA21x2_ASAP7_75t_L g3529 ( 
.A1(n_3370),
.A2(n_3230),
.B(n_3330),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3402),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3402),
.Y(n_3531)
);

AO21x2_ASAP7_75t_L g3532 ( 
.A1(n_3381),
.A2(n_3292),
.B(n_3345),
.Y(n_3532)
);

OAI21x1_ASAP7_75t_L g3533 ( 
.A1(n_3440),
.A2(n_3321),
.B(n_3342),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3372),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_3372),
.Y(n_3535)
);

OR2x6_ASAP7_75t_L g3536 ( 
.A(n_3411),
.B(n_3358),
.Y(n_3536)
);

INVx2_ASAP7_75t_L g3537 ( 
.A(n_3461),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_3464),
.Y(n_3538)
);

AOI22xp33_ASAP7_75t_SL g3539 ( 
.A1(n_3494),
.A2(n_3300),
.B1(n_3343),
.B2(n_3269),
.Y(n_3539)
);

BUFx6f_ASAP7_75t_L g3540 ( 
.A(n_3435),
.Y(n_3540)
);

INVx2_ASAP7_75t_L g3541 ( 
.A(n_3464),
.Y(n_3541)
);

A2O1A1Ixp33_ASAP7_75t_L g3542 ( 
.A1(n_3494),
.A2(n_3242),
.B(n_3349),
.C(n_3298),
.Y(n_3542)
);

OAI211xp5_ASAP7_75t_L g3543 ( 
.A1(n_3481),
.A2(n_3346),
.B(n_3246),
.C(n_3242),
.Y(n_3543)
);

OR2x2_ASAP7_75t_L g3544 ( 
.A(n_3425),
.B(n_3247),
.Y(n_3544)
);

AOI21xp5_ASAP7_75t_L g3545 ( 
.A1(n_3492),
.A2(n_3241),
.B(n_3334),
.Y(n_3545)
);

OA21x2_ASAP7_75t_L g3546 ( 
.A1(n_3465),
.A2(n_3236),
.B(n_3360),
.Y(n_3546)
);

HB1xp67_ASAP7_75t_L g3547 ( 
.A(n_3448),
.Y(n_3547)
);

NAND4xp25_ASAP7_75t_L g3548 ( 
.A(n_3428),
.B(n_3310),
.C(n_3331),
.D(n_3337),
.Y(n_3548)
);

AND2x2_ASAP7_75t_L g3549 ( 
.A(n_3374),
.B(n_3365),
.Y(n_3549)
);

AND2x4_ASAP7_75t_L g3550 ( 
.A(n_3374),
.B(n_3326),
.Y(n_3550)
);

AOI21xp33_ASAP7_75t_L g3551 ( 
.A1(n_3478),
.A2(n_3245),
.B(n_3317),
.Y(n_3551)
);

AND2x4_ASAP7_75t_L g3552 ( 
.A(n_3483),
.B(n_3239),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3406),
.Y(n_3553)
);

INVx2_ASAP7_75t_L g3554 ( 
.A(n_3465),
.Y(n_3554)
);

AND2x4_ASAP7_75t_L g3555 ( 
.A(n_3483),
.B(n_3329),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3488),
.B(n_3142),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3406),
.Y(n_3557)
);

INVx2_ASAP7_75t_SL g3558 ( 
.A(n_3449),
.Y(n_3558)
);

AND2x2_ASAP7_75t_L g3559 ( 
.A(n_3365),
.B(n_3156),
.Y(n_3559)
);

AND4x1_ASAP7_75t_L g3560 ( 
.A(n_3475),
.B(n_3348),
.C(n_3340),
.D(n_3353),
.Y(n_3560)
);

BUFx3_ASAP7_75t_L g3561 ( 
.A(n_3467),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3408),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3408),
.Y(n_3563)
);

AOI22xp33_ASAP7_75t_L g3564 ( 
.A1(n_3477),
.A2(n_3016),
.B1(n_3027),
.B2(n_3113),
.Y(n_3564)
);

A2O1A1Ixp33_ASAP7_75t_L g3565 ( 
.A1(n_3438),
.A2(n_3055),
.B(n_3094),
.C(n_3361),
.Y(n_3565)
);

AOI221xp5_ASAP7_75t_L g3566 ( 
.A1(n_3477),
.A2(n_3129),
.B1(n_3117),
.B2(n_69),
.C(n_67),
.Y(n_3566)
);

AOI21xp5_ASAP7_75t_L g3567 ( 
.A1(n_3382),
.A2(n_3129),
.B(n_3117),
.Y(n_3567)
);

A2O1A1Ixp33_ASAP7_75t_L g3568 ( 
.A1(n_3485),
.A2(n_3424),
.B(n_3415),
.C(n_3469),
.Y(n_3568)
);

OAI21x1_ASAP7_75t_L g3569 ( 
.A1(n_3409),
.A2(n_3149),
.B(n_3155),
.Y(n_3569)
);

INVx2_ASAP7_75t_SL g3570 ( 
.A(n_3415),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3410),
.Y(n_3571)
);

INVx4_ASAP7_75t_L g3572 ( 
.A(n_3435),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3410),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3377),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_3433),
.Y(n_3575)
);

NAND3xp33_ASAP7_75t_L g3576 ( 
.A(n_3485),
.B(n_3016),
.C(n_3097),
.Y(n_3576)
);

INVx5_ASAP7_75t_SL g3577 ( 
.A(n_3435),
.Y(n_3577)
);

AOI22xp33_ASAP7_75t_SL g3578 ( 
.A1(n_3383),
.A2(n_3097),
.B1(n_3105),
.B2(n_3027),
.Y(n_3578)
);

BUFx3_ASAP7_75t_L g3579 ( 
.A(n_3415),
.Y(n_3579)
);

AND2x2_ASAP7_75t_L g3580 ( 
.A(n_3364),
.B(n_3013),
.Y(n_3580)
);

AND2x2_ASAP7_75t_L g3581 ( 
.A(n_3364),
.B(n_3013),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3421),
.Y(n_3582)
);

OR2x2_ASAP7_75t_L g3583 ( 
.A(n_3469),
.B(n_3013),
.Y(n_3583)
);

OAI221xp5_ASAP7_75t_L g3584 ( 
.A1(n_3474),
.A2(n_3105),
.B1(n_3113),
.B2(n_3060),
.C(n_3276),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3388),
.Y(n_3585)
);

NAND4xp25_ASAP7_75t_SL g3586 ( 
.A(n_3473),
.B(n_70),
.C(n_68),
.D(n_69),
.Y(n_3586)
);

AOI211xp5_ASAP7_75t_L g3587 ( 
.A1(n_3382),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3488),
.B(n_3060),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3388),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_3433),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3433),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3390),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3390),
.Y(n_3593)
);

OA21x2_ASAP7_75t_L g3594 ( 
.A1(n_3472),
.A2(n_3187),
.B(n_3179),
.Y(n_3594)
);

OAI22xp5_ASAP7_75t_L g3595 ( 
.A1(n_3452),
.A2(n_3276),
.B1(n_3244),
.B2(n_3158),
.Y(n_3595)
);

INVx2_ASAP7_75t_SL g3596 ( 
.A(n_3442),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3424),
.A2(n_3244),
.B(n_3118),
.Y(n_3597)
);

AOI22xp5_ASAP7_75t_L g3598 ( 
.A1(n_3394),
.A2(n_3172),
.B1(n_3158),
.B2(n_3130),
.Y(n_3598)
);

BUFx3_ASAP7_75t_L g3599 ( 
.A(n_3442),
.Y(n_3599)
);

INVx2_ASAP7_75t_L g3600 ( 
.A(n_3437),
.Y(n_3600)
);

BUFx3_ASAP7_75t_L g3601 ( 
.A(n_3442),
.Y(n_3601)
);

BUFx3_ASAP7_75t_L g3602 ( 
.A(n_3442),
.Y(n_3602)
);

INVxp67_ASAP7_75t_SL g3603 ( 
.A(n_3472),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3437),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3392),
.Y(n_3605)
);

AND2x2_ASAP7_75t_L g3606 ( 
.A(n_3369),
.B(n_3172),
.Y(n_3606)
);

OAI22xp33_ASAP7_75t_L g3607 ( 
.A1(n_3442),
.A2(n_3130),
.B1(n_74),
.B2(n_71),
.Y(n_3607)
);

AOI21xp5_ASAP7_75t_L g3608 ( 
.A1(n_3373),
.A2(n_3400),
.B(n_3473),
.Y(n_3608)
);

BUFx3_ASAP7_75t_L g3609 ( 
.A(n_3483),
.Y(n_3609)
);

INVx2_ASAP7_75t_L g3610 ( 
.A(n_3437),
.Y(n_3610)
);

BUFx2_ASAP7_75t_L g3611 ( 
.A(n_3362),
.Y(n_3611)
);

BUFx6f_ASAP7_75t_L g3612 ( 
.A(n_3362),
.Y(n_3612)
);

O2A1O1Ixp33_ASAP7_75t_L g3613 ( 
.A1(n_3474),
.A2(n_76),
.B(n_73),
.C(n_74),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3392),
.Y(n_3614)
);

OA21x2_ASAP7_75t_L g3615 ( 
.A1(n_3476),
.A2(n_3135),
.B(n_3198),
.Y(n_3615)
);

OAI21x1_ASAP7_75t_L g3616 ( 
.A1(n_3409),
.A2(n_2689),
.B(n_2706),
.Y(n_3616)
);

AOI211xp5_ASAP7_75t_L g3617 ( 
.A1(n_3491),
.A2(n_79),
.B(n_76),
.C(n_78),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3398),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3398),
.Y(n_3619)
);

AOI22xp33_ASAP7_75t_L g3620 ( 
.A1(n_3400),
.A2(n_2619),
.B1(n_2633),
.B2(n_2632),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3412),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3412),
.Y(n_3622)
);

HB1xp67_ASAP7_75t_L g3623 ( 
.A(n_3526),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3507),
.B(n_3369),
.Y(n_3624)
);

AND2x2_ASAP7_75t_L g3625 ( 
.A(n_3549),
.B(n_3369),
.Y(n_3625)
);

OAI221xp5_ASAP7_75t_L g3626 ( 
.A1(n_3509),
.A2(n_3403),
.B1(n_3468),
.B2(n_3466),
.C(n_3367),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3497),
.Y(n_3627)
);

NAND3xp33_ASAP7_75t_L g3628 ( 
.A(n_3509),
.B(n_3484),
.C(n_3455),
.Y(n_3628)
);

AOI22xp5_ASAP7_75t_L g3629 ( 
.A1(n_3501),
.A2(n_3394),
.B1(n_3491),
.B2(n_3482),
.Y(n_3629)
);

HB1xp67_ASAP7_75t_L g3630 ( 
.A(n_3526),
.Y(n_3630)
);

AOI22xp33_ASAP7_75t_L g3631 ( 
.A1(n_3501),
.A2(n_3414),
.B1(n_3400),
.B2(n_3394),
.Y(n_3631)
);

AND2x2_ASAP7_75t_L g3632 ( 
.A(n_3520),
.B(n_3414),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3498),
.Y(n_3633)
);

HB1xp67_ASAP7_75t_L g3634 ( 
.A(n_3528),
.Y(n_3634)
);

AND2x2_ASAP7_75t_L g3635 ( 
.A(n_3558),
.B(n_3378),
.Y(n_3635)
);

INVx2_ASAP7_75t_L g3636 ( 
.A(n_3612),
.Y(n_3636)
);

AND2x4_ASAP7_75t_L g3637 ( 
.A(n_3561),
.B(n_3367),
.Y(n_3637)
);

AND2x2_ASAP7_75t_L g3638 ( 
.A(n_3499),
.B(n_3502),
.Y(n_3638)
);

AND2x2_ASAP7_75t_L g3639 ( 
.A(n_3550),
.B(n_3378),
.Y(n_3639)
);

HB1xp67_ASAP7_75t_L g3640 ( 
.A(n_3528),
.Y(n_3640)
);

OAI221xp5_ASAP7_75t_L g3641 ( 
.A1(n_3510),
.A2(n_3423),
.B1(n_3462),
.B2(n_3455),
.C(n_3453),
.Y(n_3641)
);

AOI31xp33_ASAP7_75t_L g3642 ( 
.A1(n_3539),
.A2(n_3401),
.A3(n_3459),
.B(n_3375),
.Y(n_3642)
);

OR2x2_ASAP7_75t_L g3643 ( 
.A(n_3544),
.B(n_3556),
.Y(n_3643)
);

NAND4xp25_ASAP7_75t_SL g3644 ( 
.A(n_3510),
.B(n_3463),
.C(n_3375),
.D(n_3487),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3505),
.B(n_3482),
.Y(n_3645)
);

AND2x2_ASAP7_75t_L g3646 ( 
.A(n_3550),
.B(n_3413),
.Y(n_3646)
);

AND2x2_ASAP7_75t_L g3647 ( 
.A(n_3555),
.B(n_3413),
.Y(n_3647)
);

NAND4xp25_ASAP7_75t_L g3648 ( 
.A(n_3505),
.B(n_3484),
.C(n_3486),
.D(n_3453),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_3612),
.Y(n_3649)
);

INVx2_ASAP7_75t_L g3650 ( 
.A(n_3612),
.Y(n_3650)
);

AND2x2_ASAP7_75t_L g3651 ( 
.A(n_3555),
.B(n_3430),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3511),
.Y(n_3652)
);

NOR2xp67_ASAP7_75t_L g3653 ( 
.A(n_3512),
.B(n_3430),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3514),
.Y(n_3654)
);

AO21x2_ASAP7_75t_L g3655 ( 
.A1(n_3608),
.A2(n_3476),
.B(n_3405),
.Y(n_3655)
);

INVx3_ASAP7_75t_L g3656 ( 
.A(n_3612),
.Y(n_3656)
);

AND2x4_ASAP7_75t_SL g3657 ( 
.A(n_3552),
.B(n_3443),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3561),
.Y(n_3658)
);

OR2x2_ASAP7_75t_L g3659 ( 
.A(n_3547),
.B(n_3517),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3523),
.Y(n_3660)
);

AND2x2_ASAP7_75t_L g3661 ( 
.A(n_3552),
.B(n_3430),
.Y(n_3661)
);

INVx3_ASAP7_75t_L g3662 ( 
.A(n_3609),
.Y(n_3662)
);

OA21x2_ASAP7_75t_L g3663 ( 
.A1(n_3504),
.A2(n_3405),
.B(n_3389),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3525),
.Y(n_3664)
);

AND2x2_ASAP7_75t_L g3665 ( 
.A(n_3559),
.B(n_3431),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3611),
.Y(n_3666)
);

NAND4xp25_ASAP7_75t_L g3667 ( 
.A(n_3539),
.B(n_3487),
.C(n_3399),
.D(n_3376),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_3570),
.B(n_3431),
.Y(n_3668)
);

INVx1_ASAP7_75t_SL g3669 ( 
.A(n_3512),
.Y(n_3669)
);

OR2x2_ASAP7_75t_L g3670 ( 
.A(n_3547),
.B(n_3363),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3513),
.Y(n_3671)
);

INVx5_ASAP7_75t_SL g3672 ( 
.A(n_3536),
.Y(n_3672)
);

AOI22xp33_ASAP7_75t_L g3673 ( 
.A1(n_3515),
.A2(n_3401),
.B1(n_3471),
.B2(n_3454),
.Y(n_3673)
);

AND2x4_ASAP7_75t_L g3674 ( 
.A(n_3609),
.B(n_3389),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3530),
.Y(n_3675)
);

NAND2xp33_ASAP7_75t_L g3676 ( 
.A(n_3542),
.B(n_3401),
.Y(n_3676)
);

NAND3xp33_ASAP7_75t_L g3677 ( 
.A(n_3560),
.B(n_3460),
.C(n_3441),
.Y(n_3677)
);

AOI22xp33_ASAP7_75t_L g3678 ( 
.A1(n_3503),
.A2(n_3401),
.B1(n_3471),
.B2(n_3405),
.Y(n_3678)
);

AO21x2_ASAP7_75t_L g3679 ( 
.A1(n_3568),
.A2(n_3416),
.B(n_3389),
.Y(n_3679)
);

NAND2x1_ASAP7_75t_SL g3680 ( 
.A(n_3524),
.B(n_3416),
.Y(n_3680)
);

XNOR2xp5_ASAP7_75t_L g3681 ( 
.A(n_3617),
.B(n_3418),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3531),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3506),
.B(n_3460),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3553),
.Y(n_3684)
);

NAND3xp33_ASAP7_75t_L g3685 ( 
.A(n_3587),
.B(n_3445),
.C(n_3436),
.Y(n_3685)
);

BUFx2_ASAP7_75t_L g3686 ( 
.A(n_3536),
.Y(n_3686)
);

AND2x4_ASAP7_75t_L g3687 ( 
.A(n_3599),
.B(n_3416),
.Y(n_3687)
);

AOI21xp5_ASAP7_75t_L g3688 ( 
.A1(n_3516),
.A2(n_3385),
.B(n_3404),
.Y(n_3688)
);

OAI21x1_ASAP7_75t_L g3689 ( 
.A1(n_3518),
.A2(n_3450),
.B(n_3443),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3557),
.Y(n_3690)
);

OAI22xp5_ASAP7_75t_L g3691 ( 
.A1(n_3536),
.A2(n_3542),
.B1(n_3543),
.B2(n_3566),
.Y(n_3691)
);

AND2x2_ASAP7_75t_L g3692 ( 
.A(n_3579),
.B(n_3431),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3562),
.Y(n_3693)
);

AND2x4_ASAP7_75t_L g3694 ( 
.A(n_3599),
.B(n_3443),
.Y(n_3694)
);

INVx3_ASAP7_75t_L g3695 ( 
.A(n_3524),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3563),
.Y(n_3696)
);

AOI211xp5_ASAP7_75t_L g3697 ( 
.A1(n_3586),
.A2(n_3458),
.B(n_3463),
.C(n_3445),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3571),
.Y(n_3698)
);

INVx2_ASAP7_75t_L g3699 ( 
.A(n_3513),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3573),
.Y(n_3700)
);

INVx2_ASAP7_75t_L g3701 ( 
.A(n_3513),
.Y(n_3701)
);

BUFx2_ASAP7_75t_L g3702 ( 
.A(n_3579),
.Y(n_3702)
);

AND2x4_ASAP7_75t_SL g3703 ( 
.A(n_3572),
.B(n_3450),
.Y(n_3703)
);

AND2x4_ASAP7_75t_L g3704 ( 
.A(n_3601),
.B(n_3450),
.Y(n_3704)
);

AND2x2_ASAP7_75t_L g3705 ( 
.A(n_3577),
.B(n_3384),
.Y(n_3705)
);

AND2x4_ASAP7_75t_L g3706 ( 
.A(n_3601),
.B(n_3420),
.Y(n_3706)
);

AOI221xp5_ASAP7_75t_L g3707 ( 
.A1(n_3613),
.A2(n_3434),
.B1(n_3380),
.B2(n_3457),
.C(n_3456),
.Y(n_3707)
);

HB1xp67_ASAP7_75t_L g3708 ( 
.A(n_3585),
.Y(n_3708)
);

OR2x2_ASAP7_75t_L g3709 ( 
.A(n_3546),
.B(n_3363),
.Y(n_3709)
);

AOI221xp5_ASAP7_75t_L g3710 ( 
.A1(n_3551),
.A2(n_3380),
.B1(n_3457),
.B2(n_3420),
.C(n_3426),
.Y(n_3710)
);

HB1xp67_ASAP7_75t_L g3711 ( 
.A(n_3589),
.Y(n_3711)
);

OAI33xp33_ASAP7_75t_L g3712 ( 
.A1(n_3607),
.A2(n_3395),
.A3(n_3426),
.B1(n_3422),
.B2(n_3397),
.B3(n_3429),
.Y(n_3712)
);

OAI22xp5_ASAP7_75t_L g3713 ( 
.A1(n_3568),
.A2(n_3470),
.B1(n_3397),
.B2(n_3379),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3574),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3577),
.B(n_3384),
.Y(n_3715)
);

INVx5_ASAP7_75t_L g3716 ( 
.A(n_3513),
.Y(n_3716)
);

AOI22xp33_ASAP7_75t_L g3717 ( 
.A1(n_3545),
.A2(n_3439),
.B1(n_3447),
.B2(n_3422),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3582),
.Y(n_3718)
);

OAI22xp5_ASAP7_75t_SL g3719 ( 
.A1(n_3578),
.A2(n_3419),
.B1(n_3432),
.B2(n_3429),
.Y(n_3719)
);

NOR3xp33_ASAP7_75t_L g3720 ( 
.A(n_3607),
.B(n_3447),
.C(n_3439),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3567),
.B(n_3432),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3592),
.Y(n_3722)
);

INVxp67_ASAP7_75t_L g3723 ( 
.A(n_3602),
.Y(n_3723)
);

AND2x2_ASAP7_75t_L g3724 ( 
.A(n_3577),
.B(n_3379),
.Y(n_3724)
);

NOR2xp33_ASAP7_75t_SL g3725 ( 
.A(n_3572),
.B(n_3396),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_3596),
.B(n_3451),
.Y(n_3726)
);

AOI33xp33_ASAP7_75t_L g3727 ( 
.A1(n_3578),
.A2(n_3458),
.A3(n_3419),
.B1(n_3451),
.B2(n_3396),
.B3(n_81),
.Y(n_3727)
);

OR2x2_ASAP7_75t_L g3728 ( 
.A(n_3546),
.B(n_3395),
.Y(n_3728)
);

INVx2_ASAP7_75t_L g3729 ( 
.A(n_3540),
.Y(n_3729)
);

OAI22xp5_ASAP7_75t_L g3730 ( 
.A1(n_3565),
.A2(n_3576),
.B1(n_3519),
.B2(n_3564),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3593),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3602),
.B(n_3386),
.Y(n_3732)
);

AND2x4_ASAP7_75t_L g3733 ( 
.A(n_3540),
.B(n_3419),
.Y(n_3733)
);

AND2x4_ASAP7_75t_L g3734 ( 
.A(n_3540),
.B(n_3386),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3521),
.B(n_3418),
.Y(n_3735)
);

AND2x2_ASAP7_75t_L g3736 ( 
.A(n_3521),
.B(n_2633),
.Y(n_3736)
);

HB1xp67_ASAP7_75t_L g3737 ( 
.A(n_3605),
.Y(n_3737)
);

AND2x2_ASAP7_75t_L g3738 ( 
.A(n_3672),
.B(n_3532),
.Y(n_3738)
);

HB1xp67_ASAP7_75t_L g3739 ( 
.A(n_3623),
.Y(n_3739)
);

AND2x2_ASAP7_75t_L g3740 ( 
.A(n_3672),
.B(n_3532),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3623),
.Y(n_3741)
);

AND2x2_ASAP7_75t_L g3742 ( 
.A(n_3672),
.B(n_3540),
.Y(n_3742)
);

AND2x2_ASAP7_75t_L g3743 ( 
.A(n_3624),
.B(n_3533),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3630),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3630),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3656),
.Y(n_3746)
);

CKINVDCx20_ASAP7_75t_R g3747 ( 
.A(n_3686),
.Y(n_3747)
);

AND2x2_ASAP7_75t_L g3748 ( 
.A(n_3632),
.B(n_3575),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3634),
.Y(n_3749)
);

INVx1_ASAP7_75t_SL g3750 ( 
.A(n_3669),
.Y(n_3750)
);

AOI22xp33_ASAP7_75t_L g3751 ( 
.A1(n_3676),
.A2(n_3519),
.B1(n_3548),
.B2(n_3546),
.Y(n_3751)
);

AND2x2_ASAP7_75t_L g3752 ( 
.A(n_3657),
.B(n_3575),
.Y(n_3752)
);

AND2x2_ASAP7_75t_L g3753 ( 
.A(n_3657),
.B(n_3590),
.Y(n_3753)
);

AND2x2_ASAP7_75t_L g3754 ( 
.A(n_3647),
.B(n_3590),
.Y(n_3754)
);

INVx1_ASAP7_75t_SL g3755 ( 
.A(n_3659),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3634),
.Y(n_3756)
);

OR2x2_ASAP7_75t_L g3757 ( 
.A(n_3640),
.B(n_3670),
.Y(n_3757)
);

NOR2xp67_ASAP7_75t_SL g3758 ( 
.A(n_3716),
.B(n_3519),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_SL g3759 ( 
.A(n_3642),
.B(n_3565),
.Y(n_3759)
);

OR2x2_ASAP7_75t_L g3760 ( 
.A(n_3640),
.B(n_3614),
.Y(n_3760)
);

AND2x2_ASAP7_75t_L g3761 ( 
.A(n_3646),
.B(n_3591),
.Y(n_3761)
);

OR2x6_ASAP7_75t_L g3762 ( 
.A(n_3691),
.B(n_3591),
.Y(n_3762)
);

AND2x2_ASAP7_75t_L g3763 ( 
.A(n_3639),
.B(n_3600),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3708),
.Y(n_3764)
);

AND2x2_ASAP7_75t_L g3765 ( 
.A(n_3625),
.B(n_3638),
.Y(n_3765)
);

AND2x4_ASAP7_75t_SL g3766 ( 
.A(n_3637),
.B(n_3662),
.Y(n_3766)
);

HB1xp67_ASAP7_75t_L g3767 ( 
.A(n_3666),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3708),
.Y(n_3768)
);

AND2x2_ASAP7_75t_L g3769 ( 
.A(n_3705),
.B(n_3600),
.Y(n_3769)
);

OR2x2_ASAP7_75t_L g3770 ( 
.A(n_3643),
.B(n_3618),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_3715),
.B(n_3604),
.Y(n_3771)
);

NOR2x1_ASAP7_75t_L g3772 ( 
.A(n_3676),
.B(n_3619),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3711),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3711),
.Y(n_3774)
);

AND2x2_ASAP7_75t_L g3775 ( 
.A(n_3724),
.B(n_3604),
.Y(n_3775)
);

NOR2xp33_ASAP7_75t_L g3776 ( 
.A(n_3645),
.B(n_3583),
.Y(n_3776)
);

NOR2x1_ASAP7_75t_L g3777 ( 
.A(n_3695),
.B(n_3621),
.Y(n_3777)
);

AND2x4_ASAP7_75t_L g3778 ( 
.A(n_3653),
.B(n_3610),
.Y(n_3778)
);

AND2x2_ASAP7_75t_L g3779 ( 
.A(n_3635),
.B(n_3610),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3702),
.B(n_3580),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_3658),
.B(n_3622),
.Y(n_3781)
);

HB1xp67_ASAP7_75t_L g3782 ( 
.A(n_3666),
.Y(n_3782)
);

AND2x2_ASAP7_75t_L g3783 ( 
.A(n_3661),
.B(n_3581),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3737),
.Y(n_3784)
);

NOR2xp67_ASAP7_75t_L g3785 ( 
.A(n_3716),
.B(n_3597),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3737),
.Y(n_3786)
);

HB1xp67_ASAP7_75t_L g3787 ( 
.A(n_3636),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_3658),
.B(n_3527),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3681),
.B(n_3527),
.Y(n_3789)
);

INVx1_ASAP7_75t_SL g3790 ( 
.A(n_3637),
.Y(n_3790)
);

INVx1_ASAP7_75t_SL g3791 ( 
.A(n_3703),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3656),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3627),
.Y(n_3793)
);

AND2x2_ASAP7_75t_L g3794 ( 
.A(n_3703),
.B(n_3606),
.Y(n_3794)
);

AND2x2_ASAP7_75t_L g3795 ( 
.A(n_3651),
.B(n_3527),
.Y(n_3795)
);

NOR3xp33_ASAP7_75t_L g3796 ( 
.A(n_3628),
.B(n_3595),
.C(n_3584),
.Y(n_3796)
);

AND2x2_ASAP7_75t_L g3797 ( 
.A(n_3735),
.B(n_3527),
.Y(n_3797)
);

A2O1A1Ixp33_ASAP7_75t_L g3798 ( 
.A1(n_3727),
.A2(n_3564),
.B(n_3598),
.C(n_3588),
.Y(n_3798)
);

XNOR2xp5_ASAP7_75t_L g3799 ( 
.A(n_3629),
.B(n_78),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_3727),
.B(n_3529),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3662),
.B(n_3537),
.Y(n_3801)
);

BUFx2_ASAP7_75t_L g3802 ( 
.A(n_3680),
.Y(n_3802)
);

OAI321xp33_ASAP7_75t_L g3803 ( 
.A1(n_3730),
.A2(n_3541),
.A3(n_3538),
.B1(n_3554),
.B2(n_3537),
.C(n_3603),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3633),
.Y(n_3804)
);

AND2x4_ASAP7_75t_L g3805 ( 
.A(n_3716),
.B(n_3695),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3679),
.B(n_3538),
.Y(n_3806)
);

NAND2x1_ASAP7_75t_L g3807 ( 
.A(n_3631),
.B(n_3541),
.Y(n_3807)
);

INVx2_ASAP7_75t_L g3808 ( 
.A(n_3716),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3652),
.Y(n_3809)
);

HB1xp67_ASAP7_75t_L g3810 ( 
.A(n_3636),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3697),
.B(n_3529),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3654),
.Y(n_3812)
);

NOR3xp33_ASAP7_75t_L g3813 ( 
.A(n_3626),
.B(n_3603),
.C(n_3554),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3660),
.Y(n_3814)
);

HB1xp67_ASAP7_75t_L g3815 ( 
.A(n_3649),
.Y(n_3815)
);

INVx2_ASAP7_75t_L g3816 ( 
.A(n_3649),
.Y(n_3816)
);

AND2x2_ASAP7_75t_L g3817 ( 
.A(n_3679),
.B(n_3500),
.Y(n_3817)
);

INVxp67_ASAP7_75t_SL g3818 ( 
.A(n_3723),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3664),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3675),
.Y(n_3820)
);

INVx2_ASAP7_75t_L g3821 ( 
.A(n_3650),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3682),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3723),
.B(n_3529),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_SL g3824 ( 
.A(n_3725),
.B(n_3620),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3684),
.Y(n_3825)
);

AND2x2_ASAP7_75t_L g3826 ( 
.A(n_3692),
.B(n_3500),
.Y(n_3826)
);

AND2x2_ASAP7_75t_L g3827 ( 
.A(n_3732),
.B(n_3496),
.Y(n_3827)
);

OR2x2_ASAP7_75t_L g3828 ( 
.A(n_3709),
.B(n_3496),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3690),
.Y(n_3829)
);

AND2x2_ASAP7_75t_L g3830 ( 
.A(n_3668),
.B(n_3508),
.Y(n_3830)
);

AND2x2_ASAP7_75t_L g3831 ( 
.A(n_3765),
.B(n_3678),
.Y(n_3831)
);

INVx2_ASAP7_75t_SL g3832 ( 
.A(n_3766),
.Y(n_3832)
);

INVx1_ASAP7_75t_SL g3833 ( 
.A(n_3747),
.Y(n_3833)
);

INVx2_ASAP7_75t_L g3834 ( 
.A(n_3766),
.Y(n_3834)
);

NOR3xp33_ASAP7_75t_SL g3835 ( 
.A(n_3759),
.B(n_3644),
.C(n_3648),
.Y(n_3835)
);

AND2x2_ASAP7_75t_L g3836 ( 
.A(n_3765),
.B(n_3678),
.Y(n_3836)
);

AOI22xp5_ASAP7_75t_L g3837 ( 
.A1(n_3796),
.A2(n_3720),
.B1(n_3719),
.B2(n_3717),
.Y(n_3837)
);

NOR4xp25_ASAP7_75t_L g3838 ( 
.A(n_3803),
.B(n_3631),
.C(n_3717),
.D(n_3641),
.Y(n_3838)
);

NAND3xp33_ASAP7_75t_L g3839 ( 
.A(n_3751),
.B(n_3720),
.C(n_3673),
.Y(n_3839)
);

HB1xp67_ASAP7_75t_L g3840 ( 
.A(n_3739),
.Y(n_3840)
);

XNOR2xp5_ASAP7_75t_L g3841 ( 
.A(n_3747),
.B(n_3667),
.Y(n_3841)
);

AND2x4_ASAP7_75t_L g3842 ( 
.A(n_3805),
.B(n_3742),
.Y(n_3842)
);

NOR4xp25_ASAP7_75t_L g3843 ( 
.A(n_3750),
.B(n_3677),
.C(n_3683),
.D(n_3707),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_3818),
.B(n_3688),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3741),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3741),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3744),
.Y(n_3847)
);

XNOR2xp5_ASAP7_75t_L g3848 ( 
.A(n_3799),
.B(n_3713),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3744),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3745),
.Y(n_3850)
);

NOR3xp33_ASAP7_75t_SL g3851 ( 
.A(n_3799),
.B(n_3712),
.C(n_3710),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3745),
.Y(n_3852)
);

AOI22xp5_ASAP7_75t_L g3853 ( 
.A1(n_3762),
.A2(n_3712),
.B1(n_3673),
.B2(n_3685),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3756),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3805),
.Y(n_3855)
);

INVx2_ASAP7_75t_SL g3856 ( 
.A(n_3805),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3755),
.B(n_3714),
.Y(n_3857)
);

BUFx3_ASAP7_75t_L g3858 ( 
.A(n_3742),
.Y(n_3858)
);

XOR2x2_ASAP7_75t_L g3859 ( 
.A(n_3772),
.B(n_3655),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3756),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3764),
.Y(n_3861)
);

XOR2x2_ASAP7_75t_L g3862 ( 
.A(n_3807),
.B(n_3655),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3764),
.Y(n_3863)
);

NAND4xp75_ASAP7_75t_L g3864 ( 
.A(n_3738),
.B(n_3650),
.C(n_3663),
.D(n_3671),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3768),
.Y(n_3865)
);

XNOR2xp5_ASAP7_75t_L g3866 ( 
.A(n_3791),
.B(n_3694),
.Y(n_3866)
);

AND2x2_ASAP7_75t_L g3867 ( 
.A(n_3769),
.B(n_3665),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3768),
.Y(n_3868)
);

OR2x2_ASAP7_75t_L g3869 ( 
.A(n_3762),
.B(n_3721),
.Y(n_3869)
);

XNOR2xp5_ASAP7_75t_L g3870 ( 
.A(n_3762),
.B(n_3694),
.Y(n_3870)
);

OR2x2_ASAP7_75t_L g3871 ( 
.A(n_3762),
.B(n_3728),
.Y(n_3871)
);

XOR2x2_ASAP7_75t_L g3872 ( 
.A(n_3807),
.B(n_3694),
.Y(n_3872)
);

XOR2x2_ASAP7_75t_L g3873 ( 
.A(n_3789),
.B(n_3704),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3773),
.Y(n_3874)
);

INVx2_ASAP7_75t_L g3875 ( 
.A(n_3778),
.Y(n_3875)
);

AND2x2_ASAP7_75t_L g3876 ( 
.A(n_3769),
.B(n_3704),
.Y(n_3876)
);

INVx2_ASAP7_75t_SL g3877 ( 
.A(n_3778),
.Y(n_3877)
);

NAND4xp75_ASAP7_75t_SL g3878 ( 
.A(n_3758),
.B(n_3663),
.C(n_3736),
.D(n_3615),
.Y(n_3878)
);

AND2x2_ASAP7_75t_L g3879 ( 
.A(n_3771),
.B(n_3704),
.Y(n_3879)
);

AND2x2_ASAP7_75t_L g3880 ( 
.A(n_3771),
.B(n_3671),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_3749),
.B(n_3718),
.Y(n_3881)
);

NOR3xp33_ASAP7_75t_L g3882 ( 
.A(n_3738),
.B(n_3701),
.C(n_3699),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3773),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3774),
.Y(n_3884)
);

AND2x2_ASAP7_75t_L g3885 ( 
.A(n_3775),
.B(n_3699),
.Y(n_3885)
);

NOR4xp75_ASAP7_75t_L g3886 ( 
.A(n_3800),
.B(n_3726),
.C(n_3729),
.D(n_3701),
.Y(n_3886)
);

NOR3xp33_ASAP7_75t_SL g3887 ( 
.A(n_3798),
.B(n_3696),
.C(n_3693),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_3767),
.B(n_3698),
.Y(n_3888)
);

BUFx2_ASAP7_75t_L g3889 ( 
.A(n_3802),
.Y(n_3889)
);

CKINVDCx5p33_ASAP7_75t_R g3890 ( 
.A(n_3740),
.Y(n_3890)
);

INVxp67_ASAP7_75t_SL g3891 ( 
.A(n_3758),
.Y(n_3891)
);

OR2x2_ASAP7_75t_L g3892 ( 
.A(n_3782),
.B(n_3729),
.Y(n_3892)
);

HB1xp67_ASAP7_75t_L g3893 ( 
.A(n_3757),
.Y(n_3893)
);

INVx2_ASAP7_75t_L g3894 ( 
.A(n_3778),
.Y(n_3894)
);

OR2x2_ASAP7_75t_L g3895 ( 
.A(n_3757),
.B(n_3770),
.Y(n_3895)
);

AND2x2_ASAP7_75t_L g3896 ( 
.A(n_3775),
.B(n_3734),
.Y(n_3896)
);

NAND4xp75_ASAP7_75t_L g3897 ( 
.A(n_3740),
.B(n_3663),
.C(n_3731),
.D(n_3722),
.Y(n_3897)
);

INVxp67_ASAP7_75t_SL g3898 ( 
.A(n_3817),
.Y(n_3898)
);

INVxp67_ASAP7_75t_SL g3899 ( 
.A(n_3817),
.Y(n_3899)
);

OA22x2_ASAP7_75t_L g3900 ( 
.A1(n_3811),
.A2(n_3733),
.B1(n_3734),
.B2(n_3687),
.Y(n_3900)
);

NAND4xp75_ASAP7_75t_L g3901 ( 
.A(n_3777),
.B(n_3700),
.C(n_3615),
.D(n_3594),
.Y(n_3901)
);

AND2x2_ASAP7_75t_L g3902 ( 
.A(n_3754),
.B(n_3734),
.Y(n_3902)
);

AND2x2_ASAP7_75t_L g3903 ( 
.A(n_3754),
.B(n_3733),
.Y(n_3903)
);

BUFx3_ASAP7_75t_L g3904 ( 
.A(n_3746),
.Y(n_3904)
);

NAND4xp75_ASAP7_75t_L g3905 ( 
.A(n_3797),
.B(n_3785),
.C(n_3824),
.D(n_3795),
.Y(n_3905)
);

HB1xp67_ASAP7_75t_L g3906 ( 
.A(n_3774),
.Y(n_3906)
);

NOR3xp33_ASAP7_75t_L g3907 ( 
.A(n_3813),
.B(n_3689),
.C(n_3706),
.Y(n_3907)
);

INVx2_ASAP7_75t_L g3908 ( 
.A(n_3802),
.Y(n_3908)
);

INVx2_ASAP7_75t_SL g3909 ( 
.A(n_3752),
.Y(n_3909)
);

NAND4xp75_ASAP7_75t_SL g3910 ( 
.A(n_3797),
.B(n_3776),
.C(n_3795),
.D(n_3826),
.Y(n_3910)
);

INVx1_ASAP7_75t_SL g3911 ( 
.A(n_3790),
.Y(n_3911)
);

XNOR2x2_ASAP7_75t_L g3912 ( 
.A(n_3784),
.B(n_3508),
.Y(n_3912)
);

XOR2x2_ASAP7_75t_L g3913 ( 
.A(n_3781),
.B(n_3733),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3787),
.Y(n_3914)
);

AOI22xp5_ASAP7_75t_L g3915 ( 
.A1(n_3743),
.A2(n_3674),
.B1(n_3687),
.B2(n_3706),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3810),
.Y(n_3916)
);

AND2x2_ASAP7_75t_L g3917 ( 
.A(n_3763),
.B(n_3674),
.Y(n_3917)
);

INVxp67_ASAP7_75t_L g3918 ( 
.A(n_3815),
.Y(n_3918)
);

BUFx3_ASAP7_75t_L g3919 ( 
.A(n_3746),
.Y(n_3919)
);

AND2x2_ASAP7_75t_L g3920 ( 
.A(n_3763),
.B(n_3674),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3760),
.Y(n_3921)
);

NAND4xp75_ASAP7_75t_SL g3922 ( 
.A(n_3826),
.B(n_3615),
.C(n_3594),
.D(n_3687),
.Y(n_3922)
);

OR2x2_ASAP7_75t_L g3923 ( 
.A(n_3833),
.B(n_3770),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_L g3924 ( 
.A(n_3851),
.B(n_3786),
.Y(n_3924)
);

AND2x2_ASAP7_75t_L g3925 ( 
.A(n_3833),
.B(n_3761),
.Y(n_3925)
);

AND2x2_ASAP7_75t_L g3926 ( 
.A(n_3876),
.B(n_3761),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3893),
.Y(n_3927)
);

A2O1A1Ixp33_ASAP7_75t_L g3928 ( 
.A1(n_3887),
.A2(n_3806),
.B(n_3743),
.C(n_3788),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3879),
.B(n_3779),
.Y(n_3929)
);

INVx2_ASAP7_75t_L g3930 ( 
.A(n_3877),
.Y(n_3930)
);

OR2x2_ASAP7_75t_L g3931 ( 
.A(n_3911),
.B(n_3792),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_L g3932 ( 
.A(n_3851),
.B(n_3816),
.Y(n_3932)
);

NOR2xp33_ASAP7_75t_L g3933 ( 
.A(n_3858),
.B(n_3792),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3893),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3906),
.Y(n_3935)
);

INVx2_ASAP7_75t_L g3936 ( 
.A(n_3904),
.Y(n_3936)
);

AOI22xp33_ASAP7_75t_L g3937 ( 
.A1(n_3839),
.A2(n_3806),
.B1(n_3804),
.B2(n_3793),
.Y(n_3937)
);

AND2x2_ASAP7_75t_L g3938 ( 
.A(n_3896),
.B(n_3779),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3906),
.Y(n_3939)
);

AND2x2_ASAP7_75t_L g3940 ( 
.A(n_3903),
.B(n_3752),
.Y(n_3940)
);

INVx2_ASAP7_75t_L g3941 ( 
.A(n_3904),
.Y(n_3941)
);

OR2x2_ASAP7_75t_L g3942 ( 
.A(n_3911),
.B(n_3816),
.Y(n_3942)
);

OR2x2_ASAP7_75t_L g3943 ( 
.A(n_3844),
.B(n_3821),
.Y(n_3943)
);

AND2x2_ASAP7_75t_L g3944 ( 
.A(n_3867),
.B(n_3753),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_3887),
.B(n_3821),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3840),
.Y(n_3946)
);

INVxp67_ASAP7_75t_L g3947 ( 
.A(n_3840),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3898),
.Y(n_3948)
);

INVx2_ASAP7_75t_L g3949 ( 
.A(n_3856),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_3843),
.B(n_3918),
.Y(n_3950)
);

OR2x2_ASAP7_75t_L g3951 ( 
.A(n_3844),
.B(n_3760),
.Y(n_3951)
);

OR2x2_ASAP7_75t_L g3952 ( 
.A(n_3895),
.B(n_3808),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3918),
.B(n_3829),
.Y(n_3953)
);

NOR2xp33_ASAP7_75t_L g3954 ( 
.A(n_3890),
.B(n_3808),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3898),
.B(n_3829),
.Y(n_3955)
);

AND2x4_ASAP7_75t_L g3956 ( 
.A(n_3832),
.B(n_3753),
.Y(n_3956)
);

INVx2_ASAP7_75t_L g3957 ( 
.A(n_3842),
.Y(n_3957)
);

OR2x2_ASAP7_75t_L g3958 ( 
.A(n_3871),
.B(n_3809),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3899),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3899),
.Y(n_3960)
);

INVx2_ASAP7_75t_SL g3961 ( 
.A(n_3842),
.Y(n_3961)
);

AND2x2_ASAP7_75t_L g3962 ( 
.A(n_3902),
.B(n_3748),
.Y(n_3962)
);

AOI21xp33_ASAP7_75t_L g3963 ( 
.A1(n_3891),
.A2(n_3823),
.B(n_3828),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_L g3964 ( 
.A(n_3914),
.B(n_3812),
.Y(n_3964)
);

NAND2xp67_ASAP7_75t_SL g3965 ( 
.A(n_3880),
.B(n_3801),
.Y(n_3965)
);

OR2x2_ASAP7_75t_L g3966 ( 
.A(n_3857),
.B(n_3814),
.Y(n_3966)
);

OAI21xp33_ASAP7_75t_L g3967 ( 
.A1(n_3835),
.A2(n_3748),
.B(n_3780),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3921),
.Y(n_3968)
);

INVx1_ASAP7_75t_SL g3969 ( 
.A(n_3912),
.Y(n_3969)
);

OAI21xp33_ASAP7_75t_L g3970 ( 
.A1(n_3835),
.A2(n_3780),
.B(n_3794),
.Y(n_3970)
);

AND2x2_ASAP7_75t_L g3971 ( 
.A(n_3834),
.B(n_3794),
.Y(n_3971)
);

INVx2_ASAP7_75t_SL g3972 ( 
.A(n_3875),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3916),
.Y(n_3973)
);

INVx2_ASAP7_75t_L g3974 ( 
.A(n_3894),
.Y(n_3974)
);

OAI21xp5_ASAP7_75t_L g3975 ( 
.A1(n_3848),
.A2(n_3820),
.B(n_3819),
.Y(n_3975)
);

OR2x2_ASAP7_75t_L g3976 ( 
.A(n_3857),
.B(n_3822),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3837),
.B(n_3825),
.Y(n_3977)
);

INVx2_ASAP7_75t_L g3978 ( 
.A(n_3855),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3845),
.Y(n_3979)
);

INVx2_ASAP7_75t_L g3980 ( 
.A(n_3917),
.Y(n_3980)
);

NAND2xp33_ASAP7_75t_L g3981 ( 
.A(n_3870),
.B(n_3827),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3846),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3847),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_3853),
.B(n_3801),
.Y(n_3984)
);

AND2x2_ASAP7_75t_L g3985 ( 
.A(n_3920),
.B(n_3783),
.Y(n_3985)
);

INVxp67_ASAP7_75t_L g3986 ( 
.A(n_3891),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_3882),
.B(n_3827),
.Y(n_3987)
);

OR2x2_ASAP7_75t_L g3988 ( 
.A(n_3908),
.B(n_3828),
.Y(n_3988)
);

OR2x2_ASAP7_75t_L g3989 ( 
.A(n_3892),
.B(n_3830),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3849),
.Y(n_3990)
);

AND2x2_ASAP7_75t_L g3991 ( 
.A(n_3909),
.B(n_3783),
.Y(n_3991)
);

AND2x2_ASAP7_75t_SL g3992 ( 
.A(n_3838),
.B(n_3830),
.Y(n_3992)
);

NOR2x1_ASAP7_75t_L g3993 ( 
.A(n_3897),
.B(n_3706),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3882),
.B(n_3522),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3850),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3852),
.Y(n_3996)
);

INVx2_ASAP7_75t_L g3997 ( 
.A(n_3919),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_3885),
.B(n_3522),
.Y(n_3998)
);

AND2x4_ASAP7_75t_L g3999 ( 
.A(n_3889),
.B(n_3534),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3854),
.Y(n_4000)
);

NAND2xp33_ASAP7_75t_R g4001 ( 
.A(n_3869),
.B(n_80),
.Y(n_4001)
);

INVx2_ASAP7_75t_SL g4002 ( 
.A(n_3866),
.Y(n_4002)
);

AND2x2_ASAP7_75t_L g4003 ( 
.A(n_3831),
.B(n_3836),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3860),
.Y(n_4004)
);

NOR2xp33_ASAP7_75t_L g4005 ( 
.A(n_3841),
.B(n_3534),
.Y(n_4005)
);

AND2x2_ASAP7_75t_L g4006 ( 
.A(n_3915),
.B(n_3535),
.Y(n_4006)
);

AND2x2_ASAP7_75t_L g4007 ( 
.A(n_3913),
.B(n_3535),
.Y(n_4007)
);

OR2x2_ASAP7_75t_L g4008 ( 
.A(n_3888),
.B(n_3881),
.Y(n_4008)
);

NOR3xp33_ASAP7_75t_L g4009 ( 
.A(n_3905),
.B(n_80),
.C(n_82),
.Y(n_4009)
);

AND2x2_ASAP7_75t_L g4010 ( 
.A(n_3872),
.B(n_3569),
.Y(n_4010)
);

INVxp67_ASAP7_75t_L g4011 ( 
.A(n_3864),
.Y(n_4011)
);

INVx2_ASAP7_75t_SL g4012 ( 
.A(n_3956),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_4003),
.B(n_3873),
.Y(n_4013)
);

AOI21xp33_ASAP7_75t_L g4014 ( 
.A1(n_3969),
.A2(n_3900),
.B(n_3888),
.Y(n_4014)
);

AOI221xp5_ASAP7_75t_L g4015 ( 
.A1(n_3969),
.A2(n_3907),
.B1(n_3861),
.B2(n_3868),
.C(n_3865),
.Y(n_4015)
);

AOI22xp5_ASAP7_75t_L g4016 ( 
.A1(n_3992),
.A2(n_3859),
.B1(n_3862),
.B2(n_3907),
.Y(n_4016)
);

INVx2_ASAP7_75t_L g4017 ( 
.A(n_3956),
.Y(n_4017)
);

XNOR2xp5_ASAP7_75t_L g4018 ( 
.A(n_3925),
.B(n_3910),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3927),
.Y(n_4019)
);

AOI22xp5_ASAP7_75t_L g4020 ( 
.A1(n_4009),
.A2(n_3900),
.B1(n_3901),
.B2(n_3874),
.Y(n_4020)
);

AOI31xp33_ASAP7_75t_L g4021 ( 
.A1(n_3950),
.A2(n_3863),
.A3(n_3884),
.B(n_3883),
.Y(n_4021)
);

O2A1O1Ixp33_ASAP7_75t_L g4022 ( 
.A1(n_4009),
.A2(n_3881),
.B(n_3910),
.C(n_3886),
.Y(n_4022)
);

OR2x2_ASAP7_75t_L g4023 ( 
.A(n_3931),
.B(n_3878),
.Y(n_4023)
);

OAI21xp5_ASAP7_75t_L g4024 ( 
.A1(n_4011),
.A2(n_3878),
.B(n_3922),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3934),
.Y(n_4025)
);

INVx1_ASAP7_75t_SL g4026 ( 
.A(n_3923),
.Y(n_4026)
);

AO21x1_ASAP7_75t_L g4027 ( 
.A1(n_3950),
.A2(n_3922),
.B(n_82),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3935),
.Y(n_4028)
);

OAI21xp5_ASAP7_75t_L g4029 ( 
.A1(n_4011),
.A2(n_3594),
.B(n_3620),
.Y(n_4029)
);

AOI22xp5_ASAP7_75t_L g4030 ( 
.A1(n_3924),
.A2(n_3616),
.B1(n_2632),
.B2(n_85),
.Y(n_4030)
);

INVxp33_ASAP7_75t_L g4031 ( 
.A(n_3954),
.Y(n_4031)
);

NAND3xp33_ASAP7_75t_L g4032 ( 
.A(n_3932),
.B(n_83),
.C(n_84),
.Y(n_4032)
);

NAND3xp33_ASAP7_75t_L g4033 ( 
.A(n_3932),
.B(n_84),
.C(n_85),
.Y(n_4033)
);

OAI21xp33_ASAP7_75t_L g4034 ( 
.A1(n_3924),
.A2(n_87),
.B(n_89),
.Y(n_4034)
);

NAND3xp33_ASAP7_75t_L g4035 ( 
.A(n_3986),
.B(n_87),
.C(n_90),
.Y(n_4035)
);

A2O1A1Ixp33_ASAP7_75t_L g4036 ( 
.A1(n_3993),
.A2(n_93),
.B(n_90),
.C(n_92),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_3961),
.B(n_92),
.Y(n_4037)
);

NAND3xp33_ASAP7_75t_L g4038 ( 
.A(n_3937),
.B(n_96),
.C(n_97),
.Y(n_4038)
);

AOI21xp33_ASAP7_75t_L g4039 ( 
.A1(n_4001),
.A2(n_4002),
.B(n_3981),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_3939),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_3942),
.Y(n_4041)
);

NAND2x1_ASAP7_75t_L g4042 ( 
.A(n_3999),
.B(n_96),
.Y(n_4042)
);

NOR3xp33_ASAP7_75t_L g4043 ( 
.A(n_3954),
.B(n_98),
.C(n_99),
.Y(n_4043)
);

OAI21xp33_ASAP7_75t_L g4044 ( 
.A1(n_3970),
.A2(n_98),
.B(n_99),
.Y(n_4044)
);

OAI21xp5_ASAP7_75t_L g4045 ( 
.A1(n_3937),
.A2(n_100),
.B(n_101),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3947),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3947),
.Y(n_4047)
);

OAI22xp33_ASAP7_75t_SL g4048 ( 
.A1(n_3945),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_4048)
);

AND2x2_ASAP7_75t_L g4049 ( 
.A(n_3940),
.B(n_103),
.Y(n_4049)
);

NOR2xp67_ASAP7_75t_SL g4050 ( 
.A(n_3997),
.B(n_973),
.Y(n_4050)
);

NOR2xp33_ASAP7_75t_L g4051 ( 
.A(n_3986),
.B(n_105),
.Y(n_4051)
);

OR2x2_ASAP7_75t_L g4052 ( 
.A(n_3989),
.B(n_105),
.Y(n_4052)
);

OAI21xp5_ASAP7_75t_L g4053 ( 
.A1(n_3928),
.A2(n_106),
.B(n_107),
.Y(n_4053)
);

INVxp67_ASAP7_75t_L g4054 ( 
.A(n_3933),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3948),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_3957),
.B(n_108),
.Y(n_4056)
);

OAI22xp5_ASAP7_75t_L g4057 ( 
.A1(n_3984),
.A2(n_115),
.B1(n_112),
.B2(n_113),
.Y(n_4057)
);

INVx2_ASAP7_75t_L g4058 ( 
.A(n_3944),
.Y(n_4058)
);

OAI21xp5_ASAP7_75t_L g4059 ( 
.A1(n_3945),
.A2(n_112),
.B(n_116),
.Y(n_4059)
);

OAI21xp5_ASAP7_75t_L g4060 ( 
.A1(n_3984),
.A2(n_116),
.B(n_117),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_3962),
.Y(n_4061)
);

AOI21xp33_ASAP7_75t_SL g4062 ( 
.A1(n_3951),
.A2(n_118),
.B(n_119),
.Y(n_4062)
);

O2A1O1Ixp33_ASAP7_75t_L g4063 ( 
.A1(n_3987),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_4063)
);

NOR2xp33_ASAP7_75t_L g4064 ( 
.A(n_3952),
.B(n_120),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3959),
.Y(n_4065)
);

AOI32xp33_ASAP7_75t_L g4066 ( 
.A1(n_3967),
.A2(n_124),
.A3(n_122),
.B1(n_123),
.B2(n_125),
.Y(n_4066)
);

OAI22xp5_ASAP7_75t_L g4067 ( 
.A1(n_3977),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_4067)
);

OAI21xp5_ASAP7_75t_SL g4068 ( 
.A1(n_3975),
.A2(n_126),
.B(n_127),
.Y(n_4068)
);

INVx1_ASAP7_75t_SL g4069 ( 
.A(n_3991),
.Y(n_4069)
);

NOR2xp33_ASAP7_75t_L g4070 ( 
.A(n_3980),
.B(n_3933),
.Y(n_4070)
);

OAI211xp5_ASAP7_75t_L g4071 ( 
.A1(n_3975),
.A2(n_129),
.B(n_127),
.C(n_128),
.Y(n_4071)
);

AOI22xp5_ASAP7_75t_L g4072 ( 
.A1(n_3971),
.A2(n_132),
.B1(n_129),
.B2(n_131),
.Y(n_4072)
);

AOI22xp33_ASAP7_75t_L g4073 ( 
.A1(n_3977),
.A2(n_988),
.B1(n_973),
.B2(n_2656),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3960),
.Y(n_4074)
);

AOI22xp5_ASAP7_75t_L g4075 ( 
.A1(n_3985),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3988),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_L g4077 ( 
.A(n_3938),
.B(n_135),
.Y(n_4077)
);

AOI21xp33_ASAP7_75t_SL g4078 ( 
.A1(n_3987),
.A2(n_136),
.B(n_137),
.Y(n_4078)
);

OAI211xp5_ASAP7_75t_SL g4079 ( 
.A1(n_3963),
.A2(n_140),
.B(n_138),
.C(n_139),
.Y(n_4079)
);

AOI22xp33_ASAP7_75t_L g4080 ( 
.A1(n_4005),
.A2(n_988),
.B1(n_2657),
.B2(n_2656),
.Y(n_4080)
);

XOR2x2_ASAP7_75t_L g4081 ( 
.A(n_3929),
.B(n_138),
.Y(n_4081)
);

OAI21xp5_ASAP7_75t_L g4082 ( 
.A1(n_3963),
.A2(n_141),
.B(n_142),
.Y(n_4082)
);

OAI21xp5_ASAP7_75t_L g4083 ( 
.A1(n_4010),
.A2(n_143),
.B(n_144),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3946),
.Y(n_4084)
);

AND2x4_ASAP7_75t_L g4085 ( 
.A(n_3936),
.B(n_145),
.Y(n_4085)
);

AOI22xp5_ASAP7_75t_L g4086 ( 
.A1(n_3926),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_4086)
);

AOI21xp33_ASAP7_75t_SL g4087 ( 
.A1(n_4008),
.A2(n_3958),
.B(n_3943),
.Y(n_4087)
);

BUFx2_ASAP7_75t_L g4088 ( 
.A(n_3965),
.Y(n_4088)
);

AOI211x1_ASAP7_75t_L g4089 ( 
.A1(n_4007),
.A2(n_149),
.B(n_146),
.C(n_147),
.Y(n_4089)
);

NAND4xp25_ASAP7_75t_SL g4090 ( 
.A(n_3949),
.B(n_152),
.C(n_149),
.D(n_150),
.Y(n_4090)
);

INVx2_ASAP7_75t_L g4091 ( 
.A(n_3941),
.Y(n_4091)
);

AOI221xp5_ASAP7_75t_L g4092 ( 
.A1(n_3973),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.C(n_155),
.Y(n_4092)
);

AOI31xp33_ASAP7_75t_L g4093 ( 
.A1(n_3930),
.A2(n_157),
.A3(n_154),
.B(n_156),
.Y(n_4093)
);

OAI22xp33_ASAP7_75t_R g4094 ( 
.A1(n_3978),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_4094)
);

OR2x2_ASAP7_75t_L g4095 ( 
.A(n_4012),
.B(n_3972),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_4017),
.Y(n_4096)
);

OAI21xp33_ASAP7_75t_L g4097 ( 
.A1(n_4016),
.A2(n_4006),
.B(n_3974),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_4041),
.Y(n_4098)
);

AOI221xp5_ASAP7_75t_L g4099 ( 
.A1(n_4014),
.A2(n_3968),
.B1(n_3953),
.B2(n_3994),
.C(n_3955),
.Y(n_4099)
);

INVxp67_ASAP7_75t_L g4100 ( 
.A(n_4070),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_L g4101 ( 
.A(n_4026),
.B(n_3999),
.Y(n_4101)
);

OAI21xp5_ASAP7_75t_L g4102 ( 
.A1(n_4022),
.A2(n_3994),
.B(n_3964),
.Y(n_4102)
);

AOI21xp5_ASAP7_75t_SL g4103 ( 
.A1(n_4036),
.A2(n_3955),
.B(n_3953),
.Y(n_4103)
);

OAI31xp33_ASAP7_75t_L g4104 ( 
.A1(n_4071),
.A2(n_3966),
.A3(n_3976),
.B(n_3979),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_L g4105 ( 
.A(n_4069),
.B(n_3964),
.Y(n_4105)
);

OAI22xp5_ASAP7_75t_L g4106 ( 
.A1(n_4020),
.A2(n_3983),
.B1(n_3990),
.B2(n_3982),
.Y(n_4106)
);

AND2x2_ASAP7_75t_L g4107 ( 
.A(n_4058),
.B(n_3998),
.Y(n_4107)
);

OAI21xp33_ASAP7_75t_SL g4108 ( 
.A1(n_4015),
.A2(n_3996),
.B(n_3995),
.Y(n_4108)
);

AND2x2_ASAP7_75t_L g4109 ( 
.A(n_4031),
.B(n_4000),
.Y(n_4109)
);

AND2x2_ASAP7_75t_L g4110 ( 
.A(n_4061),
.B(n_4004),
.Y(n_4110)
);

O2A1O1Ixp33_ASAP7_75t_L g4111 ( 
.A1(n_4021),
.A2(n_4048),
.B(n_4045),
.C(n_4068),
.Y(n_4111)
);

OR2x6_ASAP7_75t_L g4112 ( 
.A(n_4054),
.B(n_158),
.Y(n_4112)
);

AOI222xp33_ASAP7_75t_L g4113 ( 
.A1(n_4053),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.C1(n_164),
.C2(n_167),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_4049),
.B(n_4088),
.Y(n_4114)
);

AOI21xp33_ASAP7_75t_L g4115 ( 
.A1(n_4013),
.A2(n_161),
.B(n_162),
.Y(n_4115)
);

AND2x2_ASAP7_75t_L g4116 ( 
.A(n_4076),
.B(n_168),
.Y(n_4116)
);

OAI22xp33_ASAP7_75t_SL g4117 ( 
.A1(n_4023),
.A2(n_4042),
.B1(n_4024),
.B2(n_4046),
.Y(n_4117)
);

OAI21xp5_ASAP7_75t_SL g4118 ( 
.A1(n_4018),
.A2(n_168),
.B(n_169),
.Y(n_4118)
);

INVx2_ASAP7_75t_SL g4119 ( 
.A(n_4085),
.Y(n_4119)
);

INVxp67_ASAP7_75t_SL g4120 ( 
.A(n_4027),
.Y(n_4120)
);

OAI322xp33_ASAP7_75t_L g4121 ( 
.A1(n_4047),
.A2(n_171),
.A3(n_172),
.B1(n_174),
.B2(n_175),
.C1(n_176),
.C2(n_177),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_4089),
.B(n_4066),
.Y(n_4122)
);

O2A1O1Ixp33_ASAP7_75t_SL g4123 ( 
.A1(n_4032),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_4085),
.Y(n_4124)
);

NOR2x1_ASAP7_75t_L g4125 ( 
.A(n_4032),
.B(n_4033),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_4037),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_4052),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_SL g4128 ( 
.A(n_4039),
.B(n_988),
.Y(n_4128)
);

INVx2_ASAP7_75t_L g4129 ( 
.A(n_4091),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_4077),
.Y(n_4130)
);

NAND2xp33_ASAP7_75t_SL g4131 ( 
.A(n_4050),
.B(n_177),
.Y(n_4131)
);

O2A1O1Ixp33_ASAP7_75t_L g4132 ( 
.A1(n_4048),
.A2(n_180),
.B(n_178),
.C(n_179),
.Y(n_4132)
);

NAND3xp33_ASAP7_75t_L g4133 ( 
.A(n_4038),
.B(n_178),
.C(n_179),
.Y(n_4133)
);

AND2x2_ASAP7_75t_L g4134 ( 
.A(n_4083),
.B(n_181),
.Y(n_4134)
);

NAND3xp33_ASAP7_75t_L g4135 ( 
.A(n_4033),
.B(n_4087),
.C(n_4082),
.Y(n_4135)
);

NAND3xp33_ASAP7_75t_SL g4136 ( 
.A(n_4063),
.B(n_181),
.C(n_182),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_4056),
.Y(n_4137)
);

HB1xp67_ASAP7_75t_L g4138 ( 
.A(n_4081),
.Y(n_4138)
);

OAI22xp33_ASAP7_75t_L g4139 ( 
.A1(n_4035),
.A2(n_186),
.B1(n_183),
.B2(n_184),
.Y(n_4139)
);

INVx2_ASAP7_75t_L g4140 ( 
.A(n_4019),
.Y(n_4140)
);

OAI311xp33_ASAP7_75t_L g4141 ( 
.A1(n_4044),
.A2(n_183),
.A3(n_184),
.B1(n_186),
.C1(n_187),
.Y(n_4141)
);

AOI222xp33_ASAP7_75t_L g4142 ( 
.A1(n_4029),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.C1(n_190),
.C2(n_191),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_4025),
.Y(n_4143)
);

OAI21xp5_ASAP7_75t_SL g4144 ( 
.A1(n_4079),
.A2(n_188),
.B(n_189),
.Y(n_4144)
);

OAI22xp33_ASAP7_75t_L g4145 ( 
.A1(n_4035),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_4055),
.Y(n_4146)
);

OAI21xp33_ASAP7_75t_L g4147 ( 
.A1(n_4084),
.A2(n_192),
.B(n_193),
.Y(n_4147)
);

AOI21xp5_ASAP7_75t_L g4148 ( 
.A1(n_4059),
.A2(n_4060),
.B(n_4057),
.Y(n_4148)
);

AOI21xp5_ASAP7_75t_L g4149 ( 
.A1(n_4034),
.A2(n_193),
.B(n_194),
.Y(n_4149)
);

AOI22xp5_ASAP7_75t_L g4150 ( 
.A1(n_4094),
.A2(n_198),
.B1(n_195),
.B2(n_196),
.Y(n_4150)
);

INVxp67_ASAP7_75t_SL g4151 ( 
.A(n_4051),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_4065),
.Y(n_4152)
);

NOR2xp33_ASAP7_75t_L g4153 ( 
.A(n_4062),
.B(n_195),
.Y(n_4153)
);

AOI32xp33_ASAP7_75t_L g4154 ( 
.A1(n_4043),
.A2(n_199),
.A3(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_4074),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_4028),
.Y(n_4156)
);

AOI21xp5_ASAP7_75t_L g4157 ( 
.A1(n_4067),
.A2(n_199),
.B(n_201),
.Y(n_4157)
);

HB1xp67_ASAP7_75t_L g4158 ( 
.A(n_4090),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_L g4159 ( 
.A(n_4078),
.B(n_202),
.Y(n_4159)
);

AND2x2_ASAP7_75t_L g4160 ( 
.A(n_4107),
.B(n_4064),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_4101),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4095),
.Y(n_4162)
);

NAND3xp33_ASAP7_75t_L g4163 ( 
.A(n_4099),
.B(n_4040),
.C(n_4092),
.Y(n_4163)
);

INVxp67_ASAP7_75t_SL g4164 ( 
.A(n_4125),
.Y(n_4164)
);

NOR2xp33_ASAP7_75t_L g4165 ( 
.A(n_4119),
.B(n_4093),
.Y(n_4165)
);

INVxp67_ASAP7_75t_L g4166 ( 
.A(n_4138),
.Y(n_4166)
);

AOI321xp33_ASAP7_75t_L g4167 ( 
.A1(n_4120),
.A2(n_4030),
.A3(n_4073),
.B1(n_4086),
.B2(n_4072),
.C(n_4075),
.Y(n_4167)
);

OAI22xp5_ASAP7_75t_L g4168 ( 
.A1(n_4135),
.A2(n_4080),
.B1(n_205),
.B2(n_203),
.Y(n_4168)
);

OR2x2_ASAP7_75t_L g4169 ( 
.A(n_4124),
.B(n_204),
.Y(n_4169)
);

AOI221xp5_ASAP7_75t_L g4170 ( 
.A1(n_4102),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.C(n_207),
.Y(n_4170)
);

AOI22xp5_ASAP7_75t_L g4171 ( 
.A1(n_4097),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_4171)
);

OAI22xp33_ASAP7_75t_L g4172 ( 
.A1(n_4118),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_4172)
);

HB1xp67_ASAP7_75t_L g4173 ( 
.A(n_4112),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4112),
.Y(n_4174)
);

AOI21xp5_ASAP7_75t_L g4175 ( 
.A1(n_4111),
.A2(n_211),
.B(n_214),
.Y(n_4175)
);

AOI221xp5_ASAP7_75t_L g4176 ( 
.A1(n_4106),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.C(n_219),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_4112),
.Y(n_4177)
);

O2A1O1Ixp33_ASAP7_75t_L g4178 ( 
.A1(n_4141),
.A2(n_219),
.B(n_216),
.C(n_218),
.Y(n_4178)
);

AOI222xp33_ASAP7_75t_L g4179 ( 
.A1(n_4108),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.C1(n_223),
.C2(n_224),
.Y(n_4179)
);

OAI21xp5_ASAP7_75t_L g4180 ( 
.A1(n_4103),
.A2(n_221),
.B(n_222),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_L g4181 ( 
.A(n_4158),
.B(n_223),
.Y(n_4181)
);

AND2x4_ASAP7_75t_L g4182 ( 
.A(n_4096),
.B(n_224),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_4116),
.Y(n_4183)
);

NAND3xp33_ASAP7_75t_L g4184 ( 
.A(n_4104),
.B(n_226),
.C(n_227),
.Y(n_4184)
);

BUFx2_ASAP7_75t_L g4185 ( 
.A(n_4131),
.Y(n_4185)
);

NOR4xp25_ASAP7_75t_L g4186 ( 
.A(n_4118),
.B(n_229),
.C(n_227),
.D(n_228),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4105),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4110),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_4109),
.Y(n_4189)
);

AOI211xp5_ASAP7_75t_L g4190 ( 
.A1(n_4117),
.A2(n_231),
.B(n_229),
.C(n_230),
.Y(n_4190)
);

INVxp67_ASAP7_75t_SL g4191 ( 
.A(n_4114),
.Y(n_4191)
);

AOI21xp33_ASAP7_75t_L g4192 ( 
.A1(n_4104),
.A2(n_230),
.B(n_232),
.Y(n_4192)
);

HB1xp67_ASAP7_75t_L g4193 ( 
.A(n_4098),
.Y(n_4193)
);

OAI22xp33_ASAP7_75t_L g4194 ( 
.A1(n_4144),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_4150),
.B(n_4153),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_4129),
.Y(n_4196)
);

AOI22xp33_ASAP7_75t_L g4197 ( 
.A1(n_4122),
.A2(n_2657),
.B1(n_2589),
.B2(n_2576),
.Y(n_4197)
);

OAI32xp33_ASAP7_75t_L g4198 ( 
.A1(n_4143),
.A2(n_236),
.A3(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_4198)
);

AND2x2_ASAP7_75t_L g4199 ( 
.A(n_4100),
.B(n_236),
.Y(n_4199)
);

AOI211xp5_ASAP7_75t_L g4200 ( 
.A1(n_4115),
.A2(n_239),
.B(n_240),
.C(n_241),
.Y(n_4200)
);

NOR4xp25_ASAP7_75t_SL g4201 ( 
.A(n_4123),
.B(n_240),
.C(n_241),
.D(n_242),
.Y(n_4201)
);

OAI322xp33_ASAP7_75t_L g4202 ( 
.A1(n_4156),
.A2(n_4146),
.A3(n_4155),
.B1(n_4152),
.B2(n_4140),
.C1(n_4148),
.C2(n_4145),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_4127),
.Y(n_4203)
);

INVx2_ASAP7_75t_L g4204 ( 
.A(n_4130),
.Y(n_4204)
);

AND2x2_ASAP7_75t_L g4205 ( 
.A(n_4134),
.B(n_243),
.Y(n_4205)
);

INVx2_ASAP7_75t_L g4206 ( 
.A(n_4126),
.Y(n_4206)
);

AOI21xp5_ASAP7_75t_L g4207 ( 
.A1(n_4132),
.A2(n_243),
.B(n_244),
.Y(n_4207)
);

AOI22xp5_ASAP7_75t_L g4208 ( 
.A1(n_4136),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_4208)
);

OAI21xp5_ASAP7_75t_SL g4209 ( 
.A1(n_4142),
.A2(n_245),
.B(n_246),
.Y(n_4209)
);

OAI221xp5_ASAP7_75t_L g4210 ( 
.A1(n_4151),
.A2(n_4154),
.B1(n_4133),
.B2(n_4137),
.C(n_4157),
.Y(n_4210)
);

OR2x2_ASAP7_75t_L g4211 ( 
.A(n_4159),
.B(n_247),
.Y(n_4211)
);

AOI221xp5_ASAP7_75t_L g4212 ( 
.A1(n_4141),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.C(n_250),
.Y(n_4212)
);

AOI21xp33_ASAP7_75t_SL g4213 ( 
.A1(n_4139),
.A2(n_249),
.B(n_250),
.Y(n_4213)
);

AOI221xp5_ASAP7_75t_L g4214 ( 
.A1(n_4121),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.C(n_254),
.Y(n_4214)
);

OAI21xp5_ASAP7_75t_L g4215 ( 
.A1(n_4149),
.A2(n_251),
.B(n_252),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_L g4216 ( 
.A(n_4113),
.B(n_253),
.Y(n_4216)
);

OAI22xp5_ASAP7_75t_L g4217 ( 
.A1(n_4147),
.A2(n_254),
.B1(n_255),
.B2(n_258),
.Y(n_4217)
);

A2O1A1Ixp33_ASAP7_75t_L g4218 ( 
.A1(n_4128),
.A2(n_255),
.B(n_259),
.C(n_260),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_4101),
.Y(n_4219)
);

AOI221xp5_ASAP7_75t_SL g4220 ( 
.A1(n_4099),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.C(n_263),
.Y(n_4220)
);

NOR3xp33_ASAP7_75t_L g4221 ( 
.A(n_4210),
.B(n_261),
.C(n_262),
.Y(n_4221)
);

OR2x2_ASAP7_75t_L g4222 ( 
.A(n_4186),
.B(n_263),
.Y(n_4222)
);

NAND3x1_ASAP7_75t_L g4223 ( 
.A(n_4180),
.B(n_264),
.C(n_265),
.Y(n_4223)
);

INVx1_ASAP7_75t_SL g4224 ( 
.A(n_4185),
.Y(n_4224)
);

AOI211xp5_ASAP7_75t_L g4225 ( 
.A1(n_4192),
.A2(n_265),
.B(n_266),
.C(n_269),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4173),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_4186),
.B(n_270),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_SL g4228 ( 
.A(n_4212),
.B(n_271),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_4174),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_SL g4230 ( 
.A(n_4178),
.B(n_271),
.Y(n_4230)
);

HB1xp67_ASAP7_75t_L g4231 ( 
.A(n_4177),
.Y(n_4231)
);

NOR4xp25_ASAP7_75t_L g4232 ( 
.A(n_4184),
.B(n_272),
.C(n_273),
.D(n_274),
.Y(n_4232)
);

AOI21xp5_ASAP7_75t_L g4233 ( 
.A1(n_4164),
.A2(n_4175),
.B(n_4191),
.Y(n_4233)
);

CKINVDCx20_ASAP7_75t_R g4234 ( 
.A(n_4166),
.Y(n_4234)
);

AOI21xp5_ASAP7_75t_L g4235 ( 
.A1(n_4207),
.A2(n_274),
.B(n_275),
.Y(n_4235)
);

AOI21xp5_ASAP7_75t_L g4236 ( 
.A1(n_4165),
.A2(n_275),
.B(n_276),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_L g4237 ( 
.A(n_4179),
.B(n_277),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_SL g4238 ( 
.A(n_4172),
.B(n_277),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_L g4239 ( 
.A(n_4162),
.B(n_278),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_L g4240 ( 
.A(n_4182),
.B(n_279),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_4169),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4181),
.Y(n_4242)
);

AOI21xp5_ASAP7_75t_L g4243 ( 
.A1(n_4163),
.A2(n_4201),
.B(n_4195),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_SL g4244 ( 
.A(n_4190),
.B(n_279),
.Y(n_4244)
);

INVx1_ASAP7_75t_SL g4245 ( 
.A(n_4205),
.Y(n_4245)
);

NAND2xp33_ASAP7_75t_L g4246 ( 
.A(n_4193),
.B(n_280),
.Y(n_4246)
);

BUFx2_ASAP7_75t_L g4247 ( 
.A(n_4182),
.Y(n_4247)
);

NOR3x1_ASAP7_75t_L g4248 ( 
.A(n_4209),
.B(n_280),
.C(n_281),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_4160),
.Y(n_4249)
);

NOR2xp33_ASAP7_75t_L g4250 ( 
.A(n_4202),
.B(n_282),
.Y(n_4250)
);

OAI21xp33_ASAP7_75t_SL g4251 ( 
.A1(n_4161),
.A2(n_282),
.B(n_283),
.Y(n_4251)
);

AOI211xp5_ASAP7_75t_L g4252 ( 
.A1(n_4209),
.A2(n_284),
.B(n_285),
.C(n_286),
.Y(n_4252)
);

NOR2xp33_ASAP7_75t_L g4253 ( 
.A(n_4219),
.B(n_284),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_4220),
.B(n_285),
.Y(n_4254)
);

NAND3xp33_ASAP7_75t_L g4255 ( 
.A(n_4220),
.B(n_287),
.C(n_288),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_L g4256 ( 
.A(n_4201),
.B(n_287),
.Y(n_4256)
);

AOI21xp5_ASAP7_75t_L g4257 ( 
.A1(n_4216),
.A2(n_290),
.B(n_292),
.Y(n_4257)
);

OAI221xp5_ASAP7_75t_L g4258 ( 
.A1(n_4167),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.C(n_296),
.Y(n_4258)
);

NAND3xp33_ASAP7_75t_SL g4259 ( 
.A(n_4170),
.B(n_293),
.C(n_294),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_4199),
.Y(n_4260)
);

NOR2xp33_ASAP7_75t_L g4261 ( 
.A(n_4194),
.B(n_295),
.Y(n_4261)
);

NAND3xp33_ASAP7_75t_SL g4262 ( 
.A(n_4176),
.B(n_296),
.C(n_297),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4188),
.Y(n_4263)
);

NAND3xp33_ASAP7_75t_SL g4264 ( 
.A(n_4171),
.B(n_297),
.C(n_298),
.Y(n_4264)
);

AOI21xp5_ASAP7_75t_L g4265 ( 
.A1(n_4215),
.A2(n_4203),
.B(n_4189),
.Y(n_4265)
);

HB1xp67_ASAP7_75t_L g4266 ( 
.A(n_4183),
.Y(n_4266)
);

NOR3xp33_ASAP7_75t_L g4267 ( 
.A(n_4187),
.B(n_298),
.C(n_299),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_4214),
.B(n_300),
.Y(n_4268)
);

AOI21xp5_ASAP7_75t_L g4269 ( 
.A1(n_4204),
.A2(n_300),
.B(n_301),
.Y(n_4269)
);

XNOR2xp5_ASAP7_75t_L g4270 ( 
.A(n_4208),
.B(n_4200),
.Y(n_4270)
);

OAI22xp5_ASAP7_75t_L g4271 ( 
.A1(n_4234),
.A2(n_4196),
.B1(n_4211),
.B2(n_4206),
.Y(n_4271)
);

AOI21xp33_ASAP7_75t_L g4272 ( 
.A1(n_4224),
.A2(n_4226),
.B(n_4231),
.Y(n_4272)
);

NAND2x1_ASAP7_75t_L g4273 ( 
.A(n_4247),
.B(n_4217),
.Y(n_4273)
);

AOI221xp5_ASAP7_75t_L g4274 ( 
.A1(n_4250),
.A2(n_4213),
.B1(n_4168),
.B2(n_4198),
.C(n_4218),
.Y(n_4274)
);

AOI211x1_ASAP7_75t_L g4275 ( 
.A1(n_4243),
.A2(n_4197),
.B(n_302),
.C(n_303),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_L g4276 ( 
.A(n_4245),
.B(n_301),
.Y(n_4276)
);

OAI21xp33_ASAP7_75t_L g4277 ( 
.A1(n_4249),
.A2(n_4270),
.B(n_4230),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_SL g4278 ( 
.A(n_4232),
.B(n_302),
.Y(n_4278)
);

OR2x2_ASAP7_75t_L g4279 ( 
.A(n_4256),
.B(n_304),
.Y(n_4279)
);

OAI221xp5_ASAP7_75t_L g4280 ( 
.A1(n_4258),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.C(n_307),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_4266),
.B(n_4229),
.Y(n_4281)
);

NOR3x1_ASAP7_75t_L g4282 ( 
.A(n_4255),
.B(n_305),
.C(n_307),
.Y(n_4282)
);

NAND2xp5_ASAP7_75t_SL g4283 ( 
.A(n_4251),
.B(n_308),
.Y(n_4283)
);

OAI211xp5_ASAP7_75t_SL g4284 ( 
.A1(n_4265),
.A2(n_308),
.B(n_309),
.C(n_310),
.Y(n_4284)
);

NOR2x1_ASAP7_75t_L g4285 ( 
.A(n_4222),
.B(n_310),
.Y(n_4285)
);

NOR4xp25_ASAP7_75t_SL g4286 ( 
.A(n_4228),
.B(n_4244),
.C(n_4238),
.D(n_4241),
.Y(n_4286)
);

OAI221xp5_ASAP7_75t_L g4287 ( 
.A1(n_4252),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.C(n_314),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_SL g4288 ( 
.A(n_4233),
.B(n_311),
.Y(n_4288)
);

O2A1O1Ixp33_ASAP7_75t_L g4289 ( 
.A1(n_4227),
.A2(n_312),
.B(n_316),
.C(n_317),
.Y(n_4289)
);

AOI21xp33_ASAP7_75t_SL g4290 ( 
.A1(n_4254),
.A2(n_319),
.B(n_320),
.Y(n_4290)
);

AOI221x1_ASAP7_75t_L g4291 ( 
.A1(n_4221),
.A2(n_321),
.B1(n_322),
.B2(n_323),
.C(n_324),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_4223),
.Y(n_4292)
);

NOR2xp33_ASAP7_75t_L g4293 ( 
.A(n_4264),
.B(n_323),
.Y(n_4293)
);

XNOR2x1_ASAP7_75t_L g4294 ( 
.A(n_4260),
.B(n_325),
.Y(n_4294)
);

NAND4xp25_ASAP7_75t_L g4295 ( 
.A(n_4248),
.B(n_327),
.C(n_332),
.D(n_333),
.Y(n_4295)
);

AOI221xp5_ASAP7_75t_L g4296 ( 
.A1(n_4259),
.A2(n_327),
.B1(n_333),
.B2(n_335),
.C(n_336),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_4236),
.B(n_335),
.Y(n_4297)
);

OAI21xp33_ASAP7_75t_L g4298 ( 
.A1(n_4263),
.A2(n_337),
.B(n_338),
.Y(n_4298)
);

AOI221xp5_ASAP7_75t_L g4299 ( 
.A1(n_4259),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.C(n_341),
.Y(n_4299)
);

NAND2xp5_ASAP7_75t_L g4300 ( 
.A(n_4225),
.B(n_341),
.Y(n_4300)
);

AOI21xp33_ASAP7_75t_L g4301 ( 
.A1(n_4242),
.A2(n_342),
.B(n_343),
.Y(n_4301)
);

OAI21xp5_ASAP7_75t_L g4302 ( 
.A1(n_4235),
.A2(n_4257),
.B(n_4237),
.Y(n_4302)
);

AOI211xp5_ASAP7_75t_SL g4303 ( 
.A1(n_4246),
.A2(n_344),
.B(n_345),
.C(n_346),
.Y(n_4303)
);

AOI21xp5_ASAP7_75t_L g4304 ( 
.A1(n_4269),
.A2(n_345),
.B(n_347),
.Y(n_4304)
);

NOR3xp33_ASAP7_75t_L g4305 ( 
.A(n_4268),
.B(n_348),
.C(n_350),
.Y(n_4305)
);

AOI22xp33_ASAP7_75t_L g4306 ( 
.A1(n_4262),
.A2(n_4264),
.B1(n_4239),
.B2(n_4261),
.Y(n_4306)
);

AOI21xp5_ASAP7_75t_SL g4307 ( 
.A1(n_4240),
.A2(n_350),
.B(n_351),
.Y(n_4307)
);

NAND3xp33_ASAP7_75t_L g4308 ( 
.A(n_4267),
.B(n_4253),
.C(n_4262),
.Y(n_4308)
);

AOI22xp33_ASAP7_75t_SL g4309 ( 
.A1(n_4281),
.A2(n_351),
.B1(n_352),
.B2(n_353),
.Y(n_4309)
);

AOI22xp5_ASAP7_75t_L g4310 ( 
.A1(n_4277),
.A2(n_352),
.B1(n_354),
.B2(n_355),
.Y(n_4310)
);

BUFx3_ASAP7_75t_L g4311 ( 
.A(n_4292),
.Y(n_4311)
);

INVx2_ASAP7_75t_L g4312 ( 
.A(n_4294),
.Y(n_4312)
);

HB1xp67_ASAP7_75t_L g4313 ( 
.A(n_4285),
.Y(n_4313)
);

OAI22x1_ASAP7_75t_L g4314 ( 
.A1(n_4283),
.A2(n_354),
.B1(n_355),
.B2(n_357),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_4279),
.Y(n_4315)
);

OAI22xp5_ASAP7_75t_L g4316 ( 
.A1(n_4306),
.A2(n_4280),
.B1(n_4308),
.B2(n_4287),
.Y(n_4316)
);

AOI22xp5_ASAP7_75t_L g4317 ( 
.A1(n_4271),
.A2(n_357),
.B1(n_2589),
.B2(n_2576),
.Y(n_4317)
);

OAI22xp5_ASAP7_75t_L g4318 ( 
.A1(n_4273),
.A2(n_367),
.B1(n_368),
.B2(n_369),
.Y(n_4318)
);

AOI22xp5_ASAP7_75t_SL g4319 ( 
.A1(n_4293),
.A2(n_370),
.B1(n_371),
.B2(n_372),
.Y(n_4319)
);

OAI211xp5_ASAP7_75t_L g4320 ( 
.A1(n_4272),
.A2(n_373),
.B(n_374),
.C(n_376),
.Y(n_4320)
);

AOI22xp5_ASAP7_75t_L g4321 ( 
.A1(n_4274),
.A2(n_4305),
.B1(n_4295),
.B2(n_4284),
.Y(n_4321)
);

OAI22x1_ASAP7_75t_L g4322 ( 
.A1(n_4278),
.A2(n_379),
.B1(n_381),
.B2(n_382),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4276),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4297),
.Y(n_4324)
);

OAI22xp5_ASAP7_75t_L g4325 ( 
.A1(n_4300),
.A2(n_384),
.B1(n_386),
.B2(n_391),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4288),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4298),
.Y(n_4327)
);

INVx1_ASAP7_75t_SL g4328 ( 
.A(n_4304),
.Y(n_4328)
);

OAI22xp5_ASAP7_75t_L g4329 ( 
.A1(n_4275),
.A2(n_394),
.B1(n_395),
.B2(n_396),
.Y(n_4329)
);

AO22x2_ASAP7_75t_L g4330 ( 
.A1(n_4291),
.A2(n_403),
.B1(n_404),
.B2(n_410),
.Y(n_4330)
);

INVx1_ASAP7_75t_SL g4331 ( 
.A(n_4301),
.Y(n_4331)
);

AOI22x1_ASAP7_75t_L g4332 ( 
.A1(n_4303),
.A2(n_4302),
.B1(n_4282),
.B2(n_4307),
.Y(n_4332)
);

AND2x2_ASAP7_75t_L g4333 ( 
.A(n_4311),
.B(n_4286),
.Y(n_4333)
);

NAND2xp33_ASAP7_75t_SL g4334 ( 
.A(n_4314),
.B(n_4303),
.Y(n_4334)
);

AOI32xp33_ASAP7_75t_L g4335 ( 
.A1(n_4328),
.A2(n_4296),
.A3(n_4299),
.B1(n_4290),
.B2(n_4289),
.Y(n_4335)
);

NOR2xp33_ASAP7_75t_L g4336 ( 
.A(n_4313),
.B(n_412),
.Y(n_4336)
);

AOI22xp5_ASAP7_75t_L g4337 ( 
.A1(n_4316),
.A2(n_2526),
.B1(n_2706),
.B2(n_1289),
.Y(n_4337)
);

NAND3xp33_ASAP7_75t_SL g4338 ( 
.A(n_4321),
.B(n_414),
.C(n_417),
.Y(n_4338)
);

OAI22xp33_ASAP7_75t_L g4339 ( 
.A1(n_4310),
.A2(n_418),
.B1(n_419),
.B2(n_422),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4330),
.Y(n_4340)
);

AOI221xp5_ASAP7_75t_L g4341 ( 
.A1(n_4318),
.A2(n_424),
.B1(n_425),
.B2(n_427),
.C(n_428),
.Y(n_4341)
);

O2A1O1Ixp33_ASAP7_75t_L g4342 ( 
.A1(n_4329),
.A2(n_429),
.B(n_431),
.C(n_435),
.Y(n_4342)
);

AOI221xp5_ASAP7_75t_L g4343 ( 
.A1(n_4322),
.A2(n_436),
.B1(n_437),
.B2(n_438),
.C(n_440),
.Y(n_4343)
);

AND2x2_ASAP7_75t_L g4344 ( 
.A(n_4312),
.B(n_441),
.Y(n_4344)
);

AOI221xp5_ASAP7_75t_L g4345 ( 
.A1(n_4330),
.A2(n_444),
.B1(n_445),
.B2(n_448),
.C(n_451),
.Y(n_4345)
);

OAI22xp33_ASAP7_75t_SL g4346 ( 
.A1(n_4332),
.A2(n_453),
.B1(n_454),
.B2(n_455),
.Y(n_4346)
);

O2A1O1Ixp5_ASAP7_75t_L g4347 ( 
.A1(n_4327),
.A2(n_456),
.B(n_458),
.C(n_460),
.Y(n_4347)
);

O2A1O1Ixp33_ASAP7_75t_SL g4348 ( 
.A1(n_4326),
.A2(n_461),
.B(n_462),
.C(n_464),
.Y(n_4348)
);

OAI221xp5_ASAP7_75t_L g4349 ( 
.A1(n_4335),
.A2(n_4331),
.B1(n_4309),
.B2(n_4323),
.C(n_4320),
.Y(n_4349)
);

A2O1A1Ixp33_ASAP7_75t_L g4350 ( 
.A1(n_4334),
.A2(n_4319),
.B(n_4315),
.C(n_4324),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4333),
.Y(n_4351)
);

AOI31xp33_ASAP7_75t_L g4352 ( 
.A1(n_4340),
.A2(n_4325),
.A3(n_4317),
.B(n_471),
.Y(n_4352)
);

OAI221xp5_ASAP7_75t_SL g4353 ( 
.A1(n_4342),
.A2(n_468),
.B1(n_470),
.B2(n_473),
.C(n_474),
.Y(n_4353)
);

INVx1_ASAP7_75t_SL g4354 ( 
.A(n_4344),
.Y(n_4354)
);

O2A1O1Ixp33_ASAP7_75t_L g4355 ( 
.A1(n_4346),
.A2(n_475),
.B(n_477),
.C(n_478),
.Y(n_4355)
);

NOR4xp25_ASAP7_75t_L g4356 ( 
.A(n_4338),
.B(n_1281),
.C(n_1289),
.D(n_1287),
.Y(n_4356)
);

OA211x2_ASAP7_75t_L g4357 ( 
.A1(n_4345),
.A2(n_1281),
.B(n_1289),
.C(n_1287),
.Y(n_4357)
);

O2A1O1Ixp5_ASAP7_75t_L g4358 ( 
.A1(n_4336),
.A2(n_1281),
.B(n_1289),
.C(n_1287),
.Y(n_4358)
);

AOI221xp5_ASAP7_75t_L g4359 ( 
.A1(n_4339),
.A2(n_1281),
.B1(n_1289),
.B2(n_1287),
.C(n_1273),
.Y(n_4359)
);

AOI211xp5_ASAP7_75t_L g4360 ( 
.A1(n_4349),
.A2(n_4348),
.B(n_4343),
.C(n_4341),
.Y(n_4360)
);

AOI311xp33_ASAP7_75t_L g4361 ( 
.A1(n_4351),
.A2(n_4347),
.A3(n_4337),
.B(n_1191),
.C(n_1185),
.Y(n_4361)
);

AOI21xp5_ASAP7_75t_L g4362 ( 
.A1(n_4350),
.A2(n_1281),
.B(n_1287),
.Y(n_4362)
);

OR2x2_ASAP7_75t_L g4363 ( 
.A(n_4354),
.B(n_4356),
.Y(n_4363)
);

NOR2xp33_ASAP7_75t_L g4364 ( 
.A(n_4352),
.B(n_1274),
.Y(n_4364)
);

NAND2x1_ASAP7_75t_SL g4365 ( 
.A(n_4357),
.B(n_1274),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_4355),
.B(n_1274),
.Y(n_4366)
);

NOR3xp33_ASAP7_75t_L g4367 ( 
.A(n_4364),
.B(n_4353),
.C(n_4359),
.Y(n_4367)
);

AND2x2_ASAP7_75t_L g4368 ( 
.A(n_4360),
.B(n_4361),
.Y(n_4368)
);

AOI21xp5_ASAP7_75t_L g4369 ( 
.A1(n_4366),
.A2(n_4358),
.B(n_1274),
.Y(n_4369)
);

NOR3x1_ASAP7_75t_L g4370 ( 
.A(n_4363),
.B(n_1273),
.C(n_1191),
.Y(n_4370)
);

AND2x2_ASAP7_75t_SL g4371 ( 
.A(n_4365),
.B(n_1273),
.Y(n_4371)
);

NAND3xp33_ASAP7_75t_L g4372 ( 
.A(n_4367),
.B(n_4362),
.C(n_1273),
.Y(n_4372)
);

NAND3xp33_ASAP7_75t_L g4373 ( 
.A(n_4368),
.B(n_4369),
.C(n_4371),
.Y(n_4373)
);

CKINVDCx20_ASAP7_75t_R g4374 ( 
.A(n_4373),
.Y(n_4374)
);

OR2x2_ASAP7_75t_L g4375 ( 
.A(n_4372),
.B(n_4370),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4374),
.Y(n_4376)
);

BUFx8_ASAP7_75t_L g4377 ( 
.A(n_4376),
.Y(n_4377)
);

OR4x1_ASAP7_75t_L g4378 ( 
.A(n_4377),
.B(n_4375),
.C(n_1134),
.D(n_1144),
.Y(n_4378)
);

AOI31xp33_ASAP7_75t_L g4379 ( 
.A1(n_4378),
.A2(n_1191),
.A3(n_1134),
.B(n_1144),
.Y(n_4379)
);

XNOR2xp5_ASAP7_75t_L g4380 ( 
.A(n_4379),
.B(n_1191),
.Y(n_4380)
);

AOI21xp5_ASAP7_75t_L g4381 ( 
.A1(n_4380),
.A2(n_1191),
.B(n_1134),
.Y(n_4381)
);

OAI21xp5_ASAP7_75t_L g4382 ( 
.A1(n_4381),
.A2(n_1333),
.B(n_1365),
.Y(n_4382)
);

XNOR2xp5_ASAP7_75t_L g4383 ( 
.A(n_4382),
.B(n_1121),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_4383),
.Y(n_4384)
);

AND2x4_ASAP7_75t_L g4385 ( 
.A(n_4383),
.B(n_1121),
.Y(n_4385)
);

AOI21xp33_ASAP7_75t_SL g4386 ( 
.A1(n_4384),
.A2(n_1121),
.B(n_1134),
.Y(n_4386)
);

AOI211xp5_ASAP7_75t_L g4387 ( 
.A1(n_4386),
.A2(n_4385),
.B(n_1144),
.C(n_1121),
.Y(n_4387)
);


endmodule