module fake_jpeg_24485_n_219 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_219);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_154;
wire n_76;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_35),
.Y(n_48)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_23),
.A2(n_18),
.B1(n_26),
.B2(n_16),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_23),
.B1(n_18),
.B2(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_28),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_43),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_46),
.A2(n_66),
.B1(n_22),
.B2(n_1),
.Y(n_86)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_61),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_53),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_24),
.C(n_31),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_18),
.B1(n_32),
.B2(n_17),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_57),
.A2(n_28),
.B1(n_29),
.B2(n_2),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_24),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_62),
.Y(n_89)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_70),
.Y(n_78)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_34),
.A2(n_21),
.B1(n_31),
.B2(n_30),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

OR2x4_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_19),
.Y(n_68)
);

OR2x2_ASAP7_75t_SL g102 ( 
.A(n_68),
.B(n_3),
.Y(n_102)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_35),
.B(n_38),
.C(n_21),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_71),
.B1(n_50),
.B2(n_47),
.Y(n_108)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_102),
.C(n_72),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_27),
.B(n_22),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_87),
.C(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_94),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_38),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_84),
.B(n_85),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_32),
.B(n_29),
.C(n_27),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_95),
.B1(n_99),
.B2(n_3),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_28),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_28),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_51),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_45),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_49),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_125)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_104),
.B(n_116),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_107),
.Y(n_133)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_108),
.A2(n_123),
.B1(n_126),
.B2(n_101),
.Y(n_149)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_112),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_71),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_114),
.B1(n_125),
.B2(n_127),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_13),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_51),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_121),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_13),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_51),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_75),
.A2(n_58),
.B1(n_8),
.B2(n_10),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_85),
.B(n_12),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_128),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_81),
.A2(n_14),
.B1(n_15),
.B2(n_11),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_79),
.A2(n_11),
.B1(n_102),
.B2(n_84),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_84),
.Y(n_128)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_132),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_98),
.C(n_91),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_136),
.Y(n_151)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_139),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_116),
.C(n_104),
.Y(n_136)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_92),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_82),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_128),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_148),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_149),
.A2(n_123),
.B1(n_121),
.B2(n_82),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_125),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_150),
.A2(n_124),
.B(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_155),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_154),
.A2(n_164),
.B(n_165),
.Y(n_178)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_119),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_147),
.C(n_130),
.Y(n_169)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_163),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_165),
.B1(n_150),
.B2(n_142),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_146),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_123),
.B(n_97),
.Y(n_165)
);

AOI22x1_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_96),
.B1(n_97),
.B2(n_115),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_139),
.B1(n_96),
.B2(n_132),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_175),
.C(n_180),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_173),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_147),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_160),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_148),
.C(n_133),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_149),
.B1(n_167),
.B2(n_162),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_141),
.C(n_107),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

BUFx2_ASAP7_75t_SL g184 ( 
.A(n_181),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_182),
.A2(n_187),
.B1(n_169),
.B2(n_157),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_144),
.C(n_164),
.Y(n_198)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_190),
.Y(n_199)
);

OA21x2_ASAP7_75t_SL g186 ( 
.A1(n_175),
.A2(n_180),
.B(n_172),
.Y(n_186)
);

NAND4xp25_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_183),
.C(n_192),
.D(n_190),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_163),
.B1(n_160),
.B2(n_167),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_133),
.C(n_154),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_188),
.A2(n_176),
.B(n_170),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_194),
.A2(n_196),
.B1(n_197),
.B2(n_185),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_191),
.B(n_137),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_138),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_168),
.B1(n_153),
.B2(n_171),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_200),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_137),
.B(n_158),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_201),
.A2(n_192),
.B(n_89),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_189),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_204),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_203),
.A2(n_135),
.B1(n_138),
.B2(n_74),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_207),
.A2(n_193),
.B(n_201),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_209),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_198),
.C(n_129),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_205),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_210),
.B(n_202),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_SL g215 ( 
.A1(n_212),
.A2(n_214),
.B(n_205),
.C(n_209),
.Y(n_215)
);

OAI221xp5_ASAP7_75t_SL g217 ( 
.A1(n_215),
.A2(n_216),
.B1(n_212),
.B2(n_83),
.C(n_89),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_213),
.A2(n_122),
.B(n_83),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_217),
.B(n_76),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_76),
.Y(n_219)
);


endmodule