module fake_jpeg_2905_n_199 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_199);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_2),
.B(n_12),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_8),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_17),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_79),
.Y(n_91)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_80),
.A2(n_74),
.B1(n_65),
.B2(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_82),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_83),
.A2(n_88),
.B1(n_94),
.B2(n_82),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_81),
.B(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_84),
.B(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_72),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_91),
.C(n_68),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_79),
.A2(n_64),
.B1(n_51),
.B2(n_77),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_69),
.B(n_57),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_59),
.B1(n_62),
.B2(n_52),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_95),
.B1(n_63),
.B2(n_74),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_51),
.B1(n_74),
.B2(n_61),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_63),
.B1(n_62),
.B2(n_54),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_92),
.A2(n_75),
.B1(n_76),
.B2(n_82),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_101),
.B1(n_110),
.B2(n_111),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_100),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_75),
.B1(n_85),
.B2(n_91),
.Y(n_101)
);

OR2x6_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_70),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_102),
.Y(n_130)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_73),
.B1(n_60),
.B2(n_66),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_71),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_112),
.B(n_0),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_5),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_61),
.B(n_55),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_129),
.B(n_10),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_109),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_118),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_71),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_102),
.B(n_22),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_127),
.B(n_132),
.C(n_16),
.D(n_18),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_21),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_24),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_102),
.A2(n_1),
.B(n_3),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_28),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_113),
.B(n_4),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_134),
.B(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_137),
.Y(n_159)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_136),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_30),
.B1(n_48),
.B2(n_47),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_146),
.B1(n_39),
.B2(n_42),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_131),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_144),
.B1(n_137),
.B2(n_146),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_9),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_141),
.B(n_132),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_131),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_36),
.B1(n_44),
.B2(n_43),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_128),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_150),
.Y(n_155)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_13),
.Y(n_150)
);

AOI32xp33_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_15),
.A3(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_152),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_142),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_157),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_129),
.B(n_126),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_163),
.A2(n_164),
.B(n_38),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_150),
.A2(n_124),
.B(n_127),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_167),
.Y(n_176)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_163),
.A2(n_138),
.B1(n_152),
.B2(n_140),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_19),
.B1(n_20),
.B2(n_23),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_171),
.A2(n_165),
.B1(n_166),
.B2(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_156),
.B(n_20),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_173),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_34),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_174),
.A2(n_40),
.B(n_41),
.Y(n_181)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

INVxp67_ASAP7_75t_SL g177 ( 
.A(n_175),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_181),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_176),
.A2(n_160),
.B1(n_158),
.B2(n_167),
.Y(n_179)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_182),
.A2(n_174),
.B1(n_169),
.B2(n_171),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_180),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_170),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_187),
.C(n_177),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_177),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_190),
.Y(n_193)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_187),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_184),
.B1(n_188),
.B2(n_186),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_192),
.B(n_189),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_194),
.B(n_193),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g197 ( 
.A(n_196),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_192),
.Y(n_198)
);

BUFx24_ASAP7_75t_SL g199 ( 
.A(n_198),
.Y(n_199)
);


endmodule