module fake_jpeg_26765_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_63),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_24),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_54),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_43),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_52),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_24),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_31),
.B1(n_29),
.B2(n_34),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_22),
.CON(n_59),
.SN(n_59)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_64),
.Y(n_103)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_65),
.Y(n_102)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_38),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_70),
.A2(n_20),
.B1(n_35),
.B2(n_36),
.Y(n_111)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_29),
.B1(n_19),
.B2(n_30),
.Y(n_74)
);

OAI22x1_ASAP7_75t_L g114 ( 
.A1(n_74),
.A2(n_86),
.B1(n_93),
.B2(n_23),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_22),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_79),
.Y(n_118)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_37),
.B1(n_45),
.B2(n_41),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_78),
.A2(n_99),
.B1(n_25),
.B2(n_21),
.Y(n_134)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_88),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_42),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_84),
.A2(n_17),
.B(n_23),
.C(n_28),
.Y(n_126)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_29),
.B1(n_19),
.B2(n_30),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_89),
.Y(n_110)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_45),
.B1(n_41),
.B2(n_37),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_92),
.A2(n_16),
.B1(n_32),
.B2(n_25),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_48),
.A2(n_19),
.B1(n_30),
.B2(n_35),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_95),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_42),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_42),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_53),
.A2(n_35),
.B1(n_20),
.B2(n_27),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_67),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_104),
.Y(n_113)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_106),
.B1(n_16),
.B2(n_32),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_96),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_116),
.Y(n_144)
);

AO22x1_ASAP7_75t_SL g112 ( 
.A1(n_70),
.A2(n_35),
.B1(n_17),
.B2(n_36),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_112),
.A2(n_81),
.B1(n_72),
.B2(n_102),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_114),
.A2(n_7),
.B1(n_13),
.B2(n_11),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_98),
.C(n_71),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_123),
.C(n_104),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g116 ( 
.A1(n_73),
.A2(n_16),
.A3(n_32),
.B1(n_34),
.B2(n_21),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_134),
.B1(n_92),
.B2(n_105),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_102),
.B1(n_33),
.B2(n_17),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_17),
.C(n_33),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_137),
.B(n_103),
.Y(n_145)
);

XNOR2x1_ASAP7_75t_L g131 ( 
.A(n_73),
.B(n_33),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_88),
.Y(n_147)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_84),
.B(n_107),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_160),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_139),
.A2(n_159),
.B1(n_161),
.B2(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_142),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_141),
.B(n_6),
.Y(n_204)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_75),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_143),
.B(n_158),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_145),
.A2(n_125),
.B(n_1),
.Y(n_192)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_146),
.B(n_149),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_147),
.B(n_133),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_137),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_151),
.B(n_153),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_77),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_114),
.A2(n_90),
.B1(n_85),
.B2(n_101),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_154),
.A2(n_157),
.B1(n_149),
.B2(n_170),
.Y(n_202)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_97),
.C(n_103),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_164),
.C(n_130),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_82),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_81),
.B1(n_102),
.B2(n_82),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_168),
.B1(n_136),
.B2(n_110),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_33),
.B1(n_23),
.B2(n_83),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_112),
.C(n_111),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_7),
.Y(n_165)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_112),
.A2(n_87),
.B(n_1),
.C(n_3),
.Y(n_166)
);

OAI31xp33_ASAP7_75t_L g187 ( 
.A1(n_166),
.A2(n_121),
.A3(n_1),
.B(n_3),
.Y(n_187)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_117),
.Y(n_182)
);

NOR2x1_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_6),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_177),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_186),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_130),
.C(n_117),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_159),
.B(n_144),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_178),
.A2(n_192),
.B(n_0),
.Y(n_231)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_188),
.Y(n_213)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_138),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_183),
.B(n_194),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_121),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_202),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_124),
.C(n_109),
.Y(n_188)
);

OAI22x1_ASAP7_75t_SL g189 ( 
.A1(n_166),
.A2(n_109),
.B1(n_136),
.B2(n_129),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_189),
.A2(n_191),
.B1(n_157),
.B2(n_155),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_8),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_199),
.Y(n_215)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_153),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_198),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_145),
.B(n_0),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_200),
.Y(n_229)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_144),
.A2(n_8),
.A3(n_13),
.B1(n_11),
.B2(n_9),
.Y(n_203)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g219 ( 
.A(n_204),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_184),
.Y(n_235)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_208),
.B(n_218),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_200),
.A2(n_164),
.B1(n_162),
.B2(n_169),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_209),
.A2(n_222),
.B1(n_232),
.B2(n_190),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_210),
.A2(n_220),
.B1(n_199),
.B2(n_178),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_173),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_6),
.B1(n_13),
.B2(n_9),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_221),
.B(n_224),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_180),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_179),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_226),
.B(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_177),
.Y(n_228)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_175),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_231),
.B(n_192),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_201),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_232)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_174),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_176),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_171),
.Y(n_240)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_242),
.Y(n_275)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

AO22x2_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_189),
.B1(n_187),
.B2(n_201),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_254),
.B1(n_232),
.B2(n_212),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_171),
.Y(n_244)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_246),
.Y(n_276)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_210),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_247),
.A2(n_248),
.B(n_212),
.Y(n_269)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_186),
.C(n_204),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_217),
.C(n_195),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_253),
.B(n_231),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_207),
.B(n_194),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_255),
.Y(n_257)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_256),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_262),
.Y(n_280)
);

NOR3xp33_ASAP7_75t_SL g260 ( 
.A(n_250),
.B(n_238),
.C(n_203),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_273),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_234),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_211),
.C(n_215),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_239),
.C(n_241),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_268),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_215),
.Y(n_268)
);

AO21x1_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_235),
.B(n_255),
.Y(n_283)
);

XNOR2x1_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_211),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_270),
.A2(n_256),
.B1(n_243),
.B2(n_242),
.Y(n_277)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_206),
.B1(n_223),
.B2(n_172),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_277),
.A2(n_279),
.B(n_267),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_270),
.A2(n_243),
.B(n_223),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_276),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_281),
.B(n_286),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_288),
.C(n_290),
.Y(n_298)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_260),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_291),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_258),
.C(n_262),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_259),
.C(n_268),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_266),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_264),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_300),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_294),
.A2(n_285),
.B(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_252),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_284),
.A2(n_267),
.B1(n_265),
.B2(n_271),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_301),
.A2(n_305),
.B1(n_306),
.B2(n_253),
.Y(n_310)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_283),
.Y(n_302)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_289),
.B(n_261),
.Y(n_304)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_277),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_279),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_303),
.A2(n_236),
.B(n_249),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_307),
.A2(n_15),
.B(n_4),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_311),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_300),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_293),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_296),
.A2(n_285),
.B1(n_172),
.B2(n_280),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_314),
.A2(n_295),
.B1(n_301),
.B2(n_297),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_280),
.C(n_219),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_315),
.B(n_298),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_317),
.B(n_322),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_319),
.B(n_321),
.Y(n_325)
);

NAND2xp33_ASAP7_75t_R g319 ( 
.A(n_313),
.B(n_294),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_297),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_323),
.B(n_15),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_326),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_320),
.B(n_316),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_323),
.B(n_308),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_328),
.A2(n_324),
.B(n_325),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_312),
.B(n_309),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_329),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_315),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_15),
.B(n_4),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_5),
.Y(n_335)
);


endmodule