module fake_jpeg_10594_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

OR2x2_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_16),
.Y(n_60)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_45),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_47),
.Y(n_59)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_31),
.B1(n_27),
.B2(n_23),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_51),
.B1(n_70),
.B2(n_26),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_50),
.B(n_58),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_31),
.B1(n_35),
.B2(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_57),
.Y(n_76)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_20),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_62),
.B(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_28),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_66),
.C(n_34),
.Y(n_111)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_28),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_21),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_35),
.B1(n_32),
.B2(n_28),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_17),
.B1(n_24),
.B2(n_29),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_31),
.B1(n_35),
.B2(n_23),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_20),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_26),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_77),
.B(n_79),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_78),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_92),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_35),
.B1(n_25),
.B2(n_32),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_56),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_19),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_96),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_63),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_89),
.Y(n_136)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_72),
.A2(n_25),
.B1(n_24),
.B2(n_33),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_102),
.B1(n_108),
.B2(n_113),
.Y(n_118)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_94),
.Y(n_140)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_19),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_66),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_99),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_104),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_44),
.B1(n_34),
.B2(n_19),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_61),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_74),
.C(n_48),
.Y(n_139)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

AO22x1_ASAP7_75t_SL g105 ( 
.A1(n_51),
.A2(n_34),
.B1(n_19),
.B2(n_21),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_69),
.B1(n_58),
.B2(n_62),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_67),
.A2(n_29),
.B1(n_17),
.B2(n_68),
.Y(n_108)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_75),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_48),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_34),
.B1(n_8),
.B2(n_10),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_117),
.A2(n_99),
.B1(n_106),
.B2(n_109),
.Y(n_145)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_53),
.A3(n_59),
.B1(n_50),
.B2(n_65),
.Y(n_121)
);

AOI32xp33_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_110),
.A3(n_75),
.B1(n_52),
.B2(n_112),
.Y(n_165)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_125),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_96),
.B(n_77),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_102),
.B(n_85),
.Y(n_157)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_130),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_74),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_128),
.B(n_79),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_141),
.B1(n_101),
.B2(n_89),
.Y(n_173)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_83),
.Y(n_162)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_60),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_139),
.C(n_142),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_105),
.A2(n_52),
.B1(n_75),
.B2(n_48),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_106),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_145),
.B(n_148),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_147),
.B(n_162),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_142),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_103),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_149),
.A2(n_157),
.B(n_163),
.Y(n_193)
);

CKINVDCx6p67_ASAP7_75t_R g151 ( 
.A(n_140),
.Y(n_151)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_78),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_164),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_143),
.A2(n_83),
.B1(n_98),
.B2(n_95),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_153),
.Y(n_210)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_161),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_104),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_156),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_94),
.B(n_48),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_98),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_88),
.C(n_116),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_131),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_132),
.C(n_125),
.Y(n_179)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_170),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_121),
.B(n_0),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_120),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_119),
.B(n_112),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_114),
.A2(n_1),
.B(n_3),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_SL g207 ( 
.A(n_171),
.B(n_176),
.C(n_163),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_11),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_175),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_8),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_114),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_128),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_118),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_190),
.C(n_169),
.Y(n_214)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_180),
.B(n_184),
.Y(n_213)
);

AND2x6_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_120),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_181),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_177),
.B(n_134),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_186),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_159),
.B(n_134),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_189),
.A2(n_208),
.B(n_146),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_129),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_196),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_135),
.Y(n_195)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_198),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_147),
.B(n_117),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_149),
.B(n_118),
.Y(n_200)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_207),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_136),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_204),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_149),
.B(n_145),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_226),
.C(n_179),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_200),
.A2(n_174),
.B1(n_173),
.B2(n_165),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_222),
.B1(n_180),
.B2(n_193),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_178),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_221),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_194),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_189),
.A2(n_168),
.B1(n_152),
.B2(n_160),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_194),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_230),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_190),
.B(n_148),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_233),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_158),
.C(n_168),
.Y(n_225)
);

OAI21xp33_ASAP7_75t_L g241 ( 
.A1(n_225),
.A2(n_195),
.B(n_209),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_169),
.Y(n_226)
);

A2O1A1O1Ixp25_ASAP7_75t_L g228 ( 
.A1(n_187),
.A2(n_144),
.B(n_157),
.C(n_155),
.D(n_171),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_186),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_183),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_146),
.B1(n_154),
.B2(n_150),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_236),
.B1(n_202),
.B2(n_192),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_188),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_206),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_144),
.Y(n_234)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_238),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_198),
.A2(n_150),
.B1(n_116),
.B2(n_167),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

OAI22x1_ASAP7_75t_SL g242 ( 
.A1(n_227),
.A2(n_208),
.B1(n_193),
.B2(n_207),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_242),
.A2(n_246),
.B1(n_259),
.B2(n_219),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_237),
.C(n_223),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_182),
.Y(n_247)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_247),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_181),
.C(n_191),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_249),
.C(n_233),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_196),
.C(n_185),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_254),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_253),
.Y(n_273)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_212),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_255),
.Y(n_276)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_256),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_218),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_229),
.B1(n_236),
.B2(n_234),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_182),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_258),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_216),
.A2(n_210),
.B1(n_202),
.B2(n_184),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_206),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_224),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_211),
.B(n_197),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_218),
.B(n_211),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_272),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_281),
.C(n_249),
.Y(n_285)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_242),
.A2(n_227),
.B(n_229),
.Y(n_269)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

XOR2x2_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_228),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_278),
.B(n_10),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_240),
.A2(n_235),
.B1(n_219),
.B2(n_222),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_275),
.A2(n_259),
.B1(n_244),
.B2(n_262),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_217),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_238),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_284),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_247),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_288),
.C(n_290),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_286),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_239),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_7),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_243),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_245),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_243),
.C(n_251),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_293),
.C(n_263),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_261),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_276),
.A2(n_250),
.B1(n_244),
.B2(n_258),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_295),
.A2(n_296),
.B1(n_278),
.B2(n_277),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_250),
.B1(n_161),
.B2(n_136),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_6),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_294),
.A2(n_268),
.B1(n_267),
.B2(n_273),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_298),
.A2(n_292),
.B1(n_290),
.B2(n_288),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_274),
.B(n_266),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_307),
.C(n_291),
.Y(n_311)
);

AND2x4_ASAP7_75t_SL g300 ( 
.A(n_295),
.B(n_274),
.Y(n_300)
);

AOI21x1_ASAP7_75t_SL g313 ( 
.A1(n_300),
.A2(n_303),
.B(n_289),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g302 ( 
.A(n_289),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_308),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_306),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_282),
.A2(n_7),
.B(n_15),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_293),
.B(n_6),
.Y(n_309)
);

AOI211xp5_ASAP7_75t_L g312 ( 
.A1(n_309),
.A2(n_310),
.B(n_300),
.C(n_305),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_310),
.A2(n_6),
.B1(n_13),
.B2(n_12),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_311),
.A2(n_317),
.B1(n_3),
.B2(n_4),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_312),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_319),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_306),
.B1(n_12),
.B2(n_13),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_136),
.C(n_3),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_1),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_14),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_301),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_316),
.C(n_4),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_325),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_324),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_3),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_313),
.B1(n_319),
.B2(n_315),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_329),
.B(n_330),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_327),
.C(n_328),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_320),
.B1(n_332),
.B2(n_5),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_5),
.B(n_317),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_5),
.Y(n_336)
);


endmodule