module fake_jpeg_9757_n_139 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

INVx6_ASAP7_75t_SL g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_33),
.Y(n_38)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_19),
.Y(n_44)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_49),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_31),
.A2(n_26),
.B1(n_25),
.B2(n_17),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_51),
.B1(n_20),
.B2(n_25),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_20),
.B1(n_19),
.B2(n_23),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_30),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_30),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_63),
.B1(n_66),
.B2(n_16),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_29),
.B1(n_37),
.B2(n_33),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_59),
.A2(n_42),
.B1(n_28),
.B2(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_16),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_0),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_0),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_37),
.B1(n_23),
.B2(n_17),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_35),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_28),
.B1(n_32),
.B2(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_68),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_67),
.A2(n_43),
.B(n_45),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_70),
.A2(n_57),
.B(n_24),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_84),
.C(n_24),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_79),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_82),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_62),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_59),
.B1(n_58),
.B2(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_30),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_92),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_54),
.B1(n_68),
.B2(n_56),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_76),
.B(n_69),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_90),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

BUFx24_ASAP7_75t_SL g90 ( 
.A(n_75),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_60),
.B1(n_57),
.B2(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_81),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_92),
.C(n_74),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_18),
.B1(n_27),
.B2(n_15),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_71),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_70),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_97),
.B(n_80),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_101),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_93),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_102),
.A2(n_98),
.B1(n_76),
.B2(n_104),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_105),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_107),
.C(n_85),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_73),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_111),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_73),
.C(n_88),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_86),
.B1(n_96),
.B2(n_72),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_86),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_72),
.A3(n_27),
.B1(n_15),
.B2(n_13),
.C1(n_50),
.C2(n_8),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_118),
.B(n_11),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_103),
.B1(n_102),
.B2(n_94),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_119),
.A2(n_27),
.B1(n_15),
.B2(n_13),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_103),
.C(n_81),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_122),
.Y(n_124)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_1),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_125),
.A2(n_126),
.B(n_119),
.Y(n_131)
);

AOI31xp67_ASAP7_75t_L g127 ( 
.A1(n_120),
.A2(n_1),
.A3(n_2),
.B(n_3),
.Y(n_127)
);

AOI21x1_ASAP7_75t_SL g130 ( 
.A1(n_127),
.A2(n_9),
.B(n_10),
.Y(n_130)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_129),
.B(n_131),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_124),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_132),
.A2(n_129),
.B1(n_2),
.B2(n_4),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_117),
.C(n_121),
.Y(n_135)
);

NAND2xp33_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_136),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_133),
.B1(n_1),
.B2(n_5),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_133),
.Y(n_139)
);


endmodule