module fake_netlist_5_1986_n_883 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_883);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_883;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_785;
wire n_316;
wire n_855;
wire n_389;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_523;
wire n_268;
wire n_315;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_525;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_501;
wire n_284;
wire n_245;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_443;
wire n_372;
wire n_293;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_854;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_385;
wire n_516;
wire n_498;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_820;
wire n_757;
wire n_307;
wire n_633;
wire n_530;
wire n_439;
wire n_556;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_804;
wire n_867;
wire n_537;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_399;
wire n_579;
wire n_394;
wire n_250;
wire n_341;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_519;
wire n_406;
wire n_470;
wire n_782;
wire n_325;
wire n_449;
wire n_862;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_831;
wire n_826;
wire n_335;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_570;
wire n_457;
wire n_514;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_218;
wire n_400;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_680;
wire n_432;
wire n_395;
wire n_553;
wire n_727;
wire n_839;
wire n_311;
wire n_813;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_477;
wire n_571;
wire n_461;
wire n_338;
wire n_693;
wire n_333;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_345;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_557;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_710;
wire n_707;
wire n_795;
wire n_695;
wire n_832;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_520;
wire n_426;
wire n_808;
wire n_409;
wire n_797;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_599;
wire n_334;
wire n_766;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_32),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_170),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_49),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_144),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_136),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_195),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_7),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_157),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_139),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_25),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_74),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_178),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_80),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_100),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_165),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_15),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_109),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_11),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_21),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_28),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_164),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_42),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_175),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_168),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_123),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_31),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_99),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_160),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_191),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_145),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_1),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_146),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_94),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_65),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_166),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_135),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_89),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_180),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_199),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_125),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_138),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_131),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_187),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_182),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_115),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_13),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_140),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_188),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_61),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_50),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_105),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_51),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_33),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_183),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_67),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_60),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_93),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_211),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_172),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_154),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_56),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_217),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_119),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_159),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_63),
.Y(n_286)
);

INVxp33_ASAP7_75t_SL g287 ( 
.A(n_130),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_13),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_53),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_5),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_82),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_21),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_48),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_85),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_77),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_83),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_127),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_137),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_114),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_12),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_210),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_171),
.B(n_129),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_190),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_113),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_19),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_184),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_95),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_14),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_202),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_151),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_169),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_204),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_97),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_68),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_118),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_73),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_155),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_64),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_25),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_79),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_126),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_78),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_71),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_173),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_186),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_212),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_147),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_91),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_45),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_81),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_185),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_193),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_108),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_86),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_200),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_122),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_216),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_75),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_106),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_30),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_152),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_58),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_128),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_121),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_116),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_88),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_149),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_32),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_134),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_196),
.Y(n_350)
);

INVxp33_ASAP7_75t_L g351 ( 
.A(n_162),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_2),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_111),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_215),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_167),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_76),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_198),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_84),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_34),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_141),
.Y(n_360)
);

BUFx5_ASAP7_75t_L g361 ( 
.A(n_133),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_36),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_20),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_26),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_102),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_104),
.Y(n_366)
);

INVx5_ASAP7_75t_L g367 ( 
.A(n_234),
.Y(n_367)
);

BUFx12f_ASAP7_75t_L g368 ( 
.A(n_270),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_234),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_288),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_288),
.Y(n_371)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_234),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_234),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_218),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_245),
.Y(n_375)
);

OA21x2_ASAP7_75t_L g376 ( 
.A1(n_280),
.A2(n_0),
.B(n_1),
.Y(n_376)
);

OAI22x1_ASAP7_75t_SL g377 ( 
.A1(n_228),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_245),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_288),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_245),
.Y(n_380)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_245),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_327),
.Y(n_382)
);

BUFx8_ASAP7_75t_L g383 ( 
.A(n_289),
.Y(n_383)
);

CKINVDCx6p67_ASAP7_75t_R g384 ( 
.A(n_237),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_225),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_239),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_327),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_3),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_221),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_313),
.B(n_4),
.Y(n_390)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_327),
.Y(n_391)
);

BUFx12f_ASAP7_75t_L g392 ( 
.A(n_240),
.Y(n_392)
);

AND2x2_ASAP7_75t_SL g393 ( 
.A(n_227),
.B(n_6),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_327),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_243),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_280),
.B(n_6),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_223),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_364),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_224),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_306),
.B(n_7),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_254),
.B(n_8),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_361),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_274),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_260),
.B(n_8),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_268),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_290),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_311),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_361),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_311),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_316),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_292),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_318),
.B(n_9),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_226),
.Y(n_414)
);

BUFx8_ASAP7_75t_SL g415 ( 
.A(n_252),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_241),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_348),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_352),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_339),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_339),
.B(n_10),
.Y(n_420)
);

BUFx12f_ASAP7_75t_L g421 ( 
.A(n_247),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_219),
.Y(n_422)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_267),
.Y(n_423)
);

BUFx12f_ASAP7_75t_L g424 ( 
.A(n_300),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_231),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_359),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_364),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_222),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_230),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_305),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_308),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_319),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_250),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g434 ( 
.A(n_329),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_256),
.B(n_15),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_253),
.Y(n_436)
);

OAI22x1_ASAP7_75t_L g437 ( 
.A1(n_340),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_259),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_261),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_362),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_330),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_302),
.B(n_52),
.Y(n_442)
);

INVx5_ASAP7_75t_L g443 ( 
.A(n_244),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_269),
.Y(n_444)
);

BUFx12f_ASAP7_75t_L g445 ( 
.A(n_232),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_271),
.Y(n_446)
);

OA21x2_ASAP7_75t_L g447 ( 
.A1(n_272),
.A2(n_18),
.B(n_19),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_220),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_276),
.Y(n_449)
);

OAI22x1_ASAP7_75t_L g450 ( 
.A1(n_278),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_357),
.B(n_24),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_351),
.B(n_24),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_282),
.B(n_26),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_286),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_291),
.B(n_27),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_299),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_287),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_301),
.Y(n_458)
);

NOR2x1_ASAP7_75t_L g459 ( 
.A(n_303),
.B(n_54),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_304),
.B(n_29),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_235),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_310),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_263),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_229),
.B(n_34),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_314),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_233),
.B(n_35),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_320),
.Y(n_467)
);

OAI21x1_ASAP7_75t_L g468 ( 
.A1(n_366),
.A2(n_57),
.B(n_55),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_236),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_325),
.Y(n_470)
);

AOI22x1_ASAP7_75t_SL g471 ( 
.A1(n_279),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_238),
.Y(n_472)
);

INVx5_ASAP7_75t_L g473 ( 
.A(n_242),
.Y(n_473)
);

CKINVDCx6p67_ASAP7_75t_R g474 ( 
.A(n_281),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_328),
.B(n_37),
.Y(n_475)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_331),
.B(n_59),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_332),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_277),
.B(n_38),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_389),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_397),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_399),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_371),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_474),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_425),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_374),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_415),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_472),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_370),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_473),
.B(n_336),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_371),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_448),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_445),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_368),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_369),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_385),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_R g496 ( 
.A(n_430),
.B(n_298),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_379),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_463),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_369),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_414),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_369),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_R g502 ( 
.A(n_430),
.B(n_246),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_435),
.B(n_295),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_R g504 ( 
.A(n_432),
.B(n_326),
.Y(n_504)
);

NOR2xp67_ASAP7_75t_L g505 ( 
.A(n_443),
.B(n_337),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_386),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_461),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_392),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_407),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_407),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_469),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_421),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_383),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_383),
.Y(n_515)
);

NOR2x1p5_ASAP7_75t_L g516 ( 
.A(n_384),
.B(n_248),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_416),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_409),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_373),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_452),
.B(n_401),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_431),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_473),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_373),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_434),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_375),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_413),
.B(n_342),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_432),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_440),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_375),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_375),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_441),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_R g532 ( 
.A(n_447),
.B(n_376),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_444),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_393),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_378),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_404),
.B(n_322),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_451),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_423),
.B(n_249),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_409),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_378),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_380),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_380),
.Y(n_542)
);

AND3x2_ASAP7_75t_L g543 ( 
.A(n_464),
.B(n_346),
.C(n_345),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_503),
.B(n_388),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_503),
.B(n_478),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_536),
.B(n_466),
.Y(n_546)
);

BUFx5_ASAP7_75t_L g547 ( 
.A(n_488),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_509),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_529),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_510),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_536),
.B(n_390),
.Y(n_551)
);

INVx4_ASAP7_75t_SL g552 ( 
.A(n_529),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_527),
.B(n_423),
.Y(n_553)
);

AO221x1_ASAP7_75t_L g554 ( 
.A1(n_532),
.A2(n_450),
.B1(n_437),
.B2(n_353),
.C(n_354),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_494),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_520),
.B(n_367),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_526),
.B(n_391),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_529),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_533),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_529),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_491),
.Y(n_561)
);

NOR3xp33_ASAP7_75t_L g562 ( 
.A(n_485),
.B(n_475),
.C(n_405),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_526),
.B(n_391),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_538),
.B(n_391),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_528),
.B(n_453),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_499),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_480),
.B(n_455),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_518),
.B(n_372),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_539),
.B(n_381),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_537),
.B(n_396),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_519),
.B(n_381),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_501),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_523),
.B(n_442),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_SL g574 ( 
.A(n_496),
.B(n_350),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_531),
.B(n_400),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_540),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_504),
.B(n_420),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_530),
.Y(n_578)
);

BUFx8_ASAP7_75t_L g579 ( 
.A(n_513),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_525),
.B(n_535),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_541),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_542),
.B(n_460),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_540),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_540),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_495),
.B(n_429),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_490),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_479),
.B(n_420),
.Y(n_587)
);

CKINVDCx11_ASAP7_75t_R g588 ( 
.A(n_486),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_540),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_506),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_482),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_497),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_489),
.B(n_410),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_543),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_481),
.Y(n_595)
);

AO221x1_ASAP7_75t_L g596 ( 
.A1(n_543),
.A2(n_355),
.B1(n_356),
.B2(n_349),
.C(n_347),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_500),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_507),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_522),
.B(n_419),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_511),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_592),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_545),
.B(n_484),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_546),
.B(n_487),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_586),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_555),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_591),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_544),
.A2(n_476),
.B1(n_447),
.B2(n_376),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_556),
.B(n_476),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_567),
.B(n_516),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_595),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_554),
.A2(n_551),
.B1(n_562),
.B2(n_596),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_566),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_565),
.A2(n_502),
.B1(n_534),
.B2(n_521),
.Y(n_613)
);

AND2x4_ASAP7_75t_SL g614 ( 
.A(n_597),
.B(n_498),
.Y(n_614)
);

BUFx4f_ASAP7_75t_SL g615 ( 
.A(n_561),
.Y(n_615)
);

OR2x6_ASAP7_75t_L g616 ( 
.A(n_597),
.B(n_493),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_567),
.B(n_395),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_578),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_585),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_588),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_590),
.B(n_517),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_582),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_591),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_583),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_577),
.B(n_508),
.Y(n_625)
);

INVx5_ASAP7_75t_L g626 ( 
.A(n_594),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_580),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_570),
.A2(n_360),
.B1(n_457),
.B2(n_524),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_573),
.A2(n_468),
.B(n_459),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_547),
.B(n_505),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_547),
.B(n_358),
.Y(n_631)
);

INVxp67_ASAP7_75t_SL g632 ( 
.A(n_549),
.Y(n_632)
);

NAND3xp33_ASAP7_75t_L g633 ( 
.A(n_575),
.B(n_458),
.C(n_446),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_593),
.B(n_365),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_581),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_598),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_587),
.B(n_514),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_572),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_549),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_553),
.B(n_438),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_574),
.A2(n_255),
.B1(n_257),
.B2(n_251),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_548),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_584),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_600),
.B(n_515),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_599),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_589),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_550),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_564),
.B(n_456),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_559),
.B(n_492),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_571),
.Y(n_650)
);

AND2x6_ASAP7_75t_L g651 ( 
.A(n_557),
.B(n_402),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_563),
.B(n_512),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_568),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_569),
.B(n_549),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_558),
.B(n_560),
.Y(n_655)
);

NAND2xp33_ASAP7_75t_L g656 ( 
.A(n_558),
.B(n_258),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_607),
.A2(n_576),
.B(n_560),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_622),
.B(n_576),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_603),
.B(n_483),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_602),
.A2(n_264),
.B1(n_265),
.B2(n_262),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_653),
.B(n_462),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_621),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_627),
.B(n_467),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_601),
.Y(n_664)
);

A2O1A1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_611),
.A2(n_439),
.B(n_433),
.C(n_470),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_654),
.A2(n_387),
.B(n_382),
.Y(n_666)
);

AND2x6_ASAP7_75t_L g667 ( 
.A(n_608),
.B(n_408),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_630),
.A2(n_655),
.B(n_629),
.Y(n_668)
);

O2A1O1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_634),
.A2(n_433),
.B(n_439),
.C(n_477),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_650),
.B(n_266),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_624),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_639),
.Y(n_672)
);

BUFx12f_ASAP7_75t_L g673 ( 
.A(n_610),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_639),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_642),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_647),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_619),
.A2(n_477),
.B(n_411),
.C(n_273),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_645),
.A2(n_394),
.B(n_275),
.Y(n_678)
);

O2A1O1Ixp5_ASAP7_75t_SL g679 ( 
.A1(n_635),
.A2(n_403),
.B(n_412),
.C(n_406),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_631),
.A2(n_284),
.B(n_285),
.C(n_283),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_626),
.B(n_636),
.Y(n_681)
);

AND3x1_ASAP7_75t_SL g682 ( 
.A(n_628),
.B(n_377),
.C(n_471),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_613),
.A2(n_294),
.B1(n_296),
.B2(n_293),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_626),
.B(n_297),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_604),
.B(n_552),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_605),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_SL g687 ( 
.A(n_615),
.B(n_579),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_620),
.Y(n_688)
);

A2O1A1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_617),
.A2(n_338),
.B(n_307),
.C(n_309),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_643),
.Y(n_690)
);

A2O1A1Ixp33_ASAP7_75t_SL g691 ( 
.A1(n_606),
.A2(n_417),
.B(n_418),
.C(n_426),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_612),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_617),
.B(n_312),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_R g694 ( 
.A(n_652),
.B(n_315),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_640),
.B(n_604),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_632),
.A2(n_344),
.B1(n_317),
.B2(n_321),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g697 ( 
.A1(n_648),
.A2(n_324),
.B(n_323),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_614),
.B(n_398),
.Y(n_698)
);

OAI21x1_ASAP7_75t_L g699 ( 
.A1(n_668),
.A2(n_646),
.B(n_623),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_672),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_673),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_662),
.B(n_625),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_698),
.Y(n_703)
);

BUFx2_ASAP7_75t_R g704 ( 
.A(n_688),
.Y(n_704)
);

OAI21xp5_ASAP7_75t_L g705 ( 
.A1(n_679),
.A2(n_633),
.B(n_651),
.Y(n_705)
);

INVx5_ASAP7_75t_L g706 ( 
.A(n_672),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_672),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_674),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_657),
.A2(n_638),
.B(n_618),
.Y(n_709)
);

INVx8_ASAP7_75t_L g710 ( 
.A(n_674),
.Y(n_710)
);

INVx5_ASAP7_75t_L g711 ( 
.A(n_674),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_685),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_664),
.Y(n_713)
);

BUFx6f_ASAP7_75t_SL g714 ( 
.A(n_685),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_659),
.B(n_644),
.Y(n_715)
);

CKINVDCx16_ASAP7_75t_R g716 ( 
.A(n_687),
.Y(n_716)
);

AO21x2_ASAP7_75t_L g717 ( 
.A1(n_665),
.A2(n_641),
.B(n_656),
.Y(n_717)
);

OAI21x1_ASAP7_75t_L g718 ( 
.A1(n_666),
.A2(n_427),
.B(n_398),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_671),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_675),
.Y(n_720)
);

INVxp67_ASAP7_75t_SL g721 ( 
.A(n_671),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_676),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_695),
.A2(n_609),
.B(n_649),
.Y(n_723)
);

INVx5_ASAP7_75t_L g724 ( 
.A(n_667),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_681),
.B(n_609),
.Y(n_725)
);

OAI21x1_ASAP7_75t_L g726 ( 
.A1(n_658),
.A2(n_651),
.B(n_637),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_682),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_686),
.Y(n_728)
);

BUFx4f_ASAP7_75t_SL g729 ( 
.A(n_684),
.Y(n_729)
);

AO21x2_ASAP7_75t_L g730 ( 
.A1(n_677),
.A2(n_680),
.B(n_661),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_690),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_663),
.A2(n_616),
.B(n_334),
.Y(n_732)
);

BUFx4f_ASAP7_75t_SL g733 ( 
.A(n_693),
.Y(n_733)
);

CKINVDCx14_ASAP7_75t_R g734 ( 
.A(n_694),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_692),
.Y(n_735)
);

INVx5_ASAP7_75t_L g736 ( 
.A(n_667),
.Y(n_736)
);

BUFx2_ASAP7_75t_SL g737 ( 
.A(n_683),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_697),
.B(n_670),
.C(n_660),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_719),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_700),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_737),
.A2(n_715),
.B1(n_738),
.B2(n_733),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_722),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_702),
.A2(n_696),
.B1(n_689),
.B2(n_333),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_703),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_713),
.Y(n_745)
);

OAI21x1_ASAP7_75t_L g746 ( 
.A1(n_699),
.A2(n_669),
.B(n_678),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_SL g747 ( 
.A1(n_725),
.A2(n_428),
.B(n_422),
.Y(n_747)
);

OAI22xp33_ASAP7_75t_L g748 ( 
.A1(n_716),
.A2(n_335),
.B1(n_341),
.B2(n_343),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_719),
.Y(n_749)
);

OAI21x1_ASAP7_75t_L g750 ( 
.A1(n_709),
.A2(n_691),
.B(n_62),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_720),
.B(n_422),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_735),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_704),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_721),
.B(n_428),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_710),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_731),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_712),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_721),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_700),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_728),
.Y(n_760)
);

NOR2x1_ASAP7_75t_R g761 ( 
.A(n_701),
.B(n_436),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_710),
.Y(n_762)
);

NAND2x1p5_ASAP7_75t_L g763 ( 
.A(n_706),
.B(n_436),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_725),
.B(n_66),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_700),
.Y(n_765)
);

NAND2x1p5_ASAP7_75t_L g766 ( 
.A(n_706),
.B(n_436),
.Y(n_766)
);

AOI21x1_ASAP7_75t_L g767 ( 
.A1(n_723),
.A2(n_465),
.B(n_454),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_706),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_729),
.A2(n_454),
.B1(n_449),
.B2(n_42),
.Y(n_769)
);

OA21x2_ASAP7_75t_L g770 ( 
.A1(n_726),
.A2(n_449),
.B(n_150),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_711),
.B(n_69),
.Y(n_771)
);

AOI222xp33_ASAP7_75t_L g772 ( 
.A1(n_727),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.C1(n_44),
.C2(n_45),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_734),
.B(n_41),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_741),
.B(n_732),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_764),
.B(n_711),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_753),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_751),
.B(n_707),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_764),
.B(n_711),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_742),
.Y(n_779)
);

NOR3xp33_ASAP7_75t_SL g780 ( 
.A(n_748),
.B(n_705),
.C(n_714),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_755),
.B(n_762),
.Y(n_781)
);

OR2x6_ASAP7_75t_L g782 ( 
.A(n_771),
.B(n_708),
.Y(n_782)
);

CKINVDCx16_ASAP7_75t_R g783 ( 
.A(n_773),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_745),
.B(n_708),
.Y(n_784)
);

OR2x6_ASAP7_75t_L g785 ( 
.A(n_757),
.B(n_718),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_772),
.A2(n_717),
.B1(n_730),
.B2(n_724),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_760),
.B(n_724),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_756),
.Y(n_788)
);

NAND2xp33_ASAP7_75t_R g789 ( 
.A(n_739),
.B(n_70),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_740),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_758),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_744),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_SL g793 ( 
.A(n_747),
.B(n_736),
.C(n_724),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_R g794 ( 
.A(n_749),
.B(n_770),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_769),
.B(n_724),
.Y(n_795)
);

OR2x6_ASAP7_75t_L g796 ( 
.A(n_759),
.B(n_736),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_759),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_743),
.A2(n_736),
.B1(n_46),
.B2(n_47),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_R g799 ( 
.A(n_765),
.B(n_72),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_752),
.B(n_754),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_754),
.Y(n_801)
);

OR2x2_ASAP7_75t_SL g802 ( 
.A(n_761),
.B(n_87),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_791),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_800),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_801),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_779),
.B(n_768),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_788),
.B(n_750),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_785),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_SL g809 ( 
.A1(n_798),
.A2(n_763),
.B1(n_766),
.B2(n_746),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_785),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_792),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_784),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_786),
.B(n_767),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_774),
.B(n_766),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_780),
.B(n_777),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_787),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_781),
.B(n_775),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_796),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_796),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_797),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_775),
.B(n_90),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_782),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_776),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_778),
.B(n_92),
.Y(n_824)
);

NOR4xp25_ASAP7_75t_SL g825 ( 
.A(n_789),
.B(n_761),
.C(n_96),
.D(n_98),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_790),
.Y(n_826)
);

OR2x2_ASAP7_75t_L g827 ( 
.A(n_795),
.B(n_101),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_782),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_793),
.B(n_103),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_783),
.B(n_214),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_799),
.B(n_213),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_810),
.B(n_808),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_804),
.B(n_812),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_808),
.B(n_794),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_805),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_811),
.B(n_802),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_808),
.B(n_107),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_803),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_805),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_815),
.B(n_110),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_815),
.B(n_112),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_814),
.B(n_117),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_806),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_814),
.B(n_120),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_807),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_813),
.B(n_124),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_833),
.B(n_816),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_838),
.Y(n_848)
);

INVx6_ASAP7_75t_L g849 ( 
.A(n_837),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_845),
.B(n_816),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_839),
.B(n_827),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_832),
.B(n_828),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_847),
.B(n_843),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_848),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_851),
.A2(n_831),
.B(n_836),
.C(n_830),
.Y(n_855)
);

OR2x6_ASAP7_75t_L g856 ( 
.A(n_849),
.B(n_834),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_855),
.A2(n_831),
.B(n_841),
.C(n_840),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_854),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_856),
.A2(n_846),
.B1(n_829),
.B2(n_837),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_853),
.A2(n_852),
.B1(n_844),
.B2(n_842),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_857),
.A2(n_809),
.B1(n_825),
.B2(n_828),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_858),
.Y(n_862)
);

OAI221xp5_ASAP7_75t_L g863 ( 
.A1(n_859),
.A2(n_850),
.B1(n_822),
.B2(n_820),
.C(n_826),
.Y(n_863)
);

OAI22xp33_ASAP7_75t_L g864 ( 
.A1(n_860),
.A2(n_819),
.B1(n_818),
.B2(n_835),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_862),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_861),
.A2(n_823),
.B(n_817),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_866),
.A2(n_863),
.B(n_864),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_865),
.Y(n_868)
);

NOR3xp33_ASAP7_75t_L g869 ( 
.A(n_868),
.B(n_824),
.C(n_821),
.Y(n_869)
);

AOI211xp5_ASAP7_75t_L g870 ( 
.A1(n_867),
.A2(n_819),
.B(n_818),
.C(n_817),
.Y(n_870)
);

OAI211xp5_ASAP7_75t_L g871 ( 
.A1(n_870),
.A2(n_132),
.B(n_142),
.C(n_143),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_869),
.Y(n_872)
);

OAI22x1_ASAP7_75t_L g873 ( 
.A1(n_872),
.A2(n_148),
.B1(n_153),
.B2(n_156),
.Y(n_873)
);

NOR2x1p5_ASAP7_75t_L g874 ( 
.A(n_871),
.B(n_158),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_873),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_875),
.Y(n_876)
);

AO22x2_ASAP7_75t_L g877 ( 
.A1(n_876),
.A2(n_874),
.B1(n_161),
.B2(n_163),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_877),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_878),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_879),
.A2(n_179),
.B(n_181),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_880),
.A2(n_189),
.B1(n_192),
.B2(n_194),
.Y(n_881)
);

OR2x6_ASAP7_75t_L g882 ( 
.A(n_881),
.B(n_203),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_882),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_883)
);


endmodule