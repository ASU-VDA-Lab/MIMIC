module fake_netlist_5_1884_n_1684 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1684);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1684;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_150;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_851;
wire n_615;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_149;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_148;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx2_ASAP7_75t_L g148 ( 
.A(n_14),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_53),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_64),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_52),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_95),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_69),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_30),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_75),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_13),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_76),
.Y(n_163)
);

BUFx10_ASAP7_75t_L g164 ( 
.A(n_113),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_79),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_82),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_83),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_43),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_40),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_93),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_20),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_46),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_12),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_90),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_88),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_121),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_115),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_41),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_126),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_122),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_46),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_65),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_21),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_141),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_35),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_11),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_129),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_57),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_85),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_29),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_71),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_30),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_78),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_128),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_89),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_34),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_74),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_19),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_25),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_26),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_22),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_51),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_66),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_124),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_97),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_137),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_86),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_32),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_12),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_80),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_103),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_92),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_140),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_112),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_108),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_91),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_22),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_25),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_14),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_26),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_98),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_36),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_32),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_110),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_145),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_120),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_67),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_144),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_96),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_45),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_44),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_60),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_44),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_77),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_63),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_23),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_135),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_21),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_117),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_45),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_6),
.Y(n_245)
);

BUFx8_ASAP7_75t_SL g246 ( 
.A(n_58),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_116),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_47),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_42),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_50),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_55),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_107),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_125),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_42),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_40),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_34),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_2),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_38),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_4),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_31),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_27),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_100),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_72),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_132),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_19),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_2),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_119),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_102),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_18),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_106),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_131),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_105),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g273 ( 
.A(n_7),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_37),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_29),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_15),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_59),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_114),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_136),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_56),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_15),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_36),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_139),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_6),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_3),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_17),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_134),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_84),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_99),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_17),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g291 ( 
.A(n_101),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_133),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_54),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_87),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_104),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_184),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_246),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_149),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_184),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_151),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_152),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_273),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_273),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_157),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_150),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_158),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_214),
.Y(n_311)
);

BUFx6f_ASAP7_75t_SL g312 ( 
.A(n_164),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_161),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_162),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_150),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_273),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_254),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_258),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_163),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_254),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_153),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_254),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_254),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_174),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_169),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_153),
.Y(n_326)
);

BUFx2_ASAP7_75t_SL g327 ( 
.A(n_177),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_254),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_148),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_148),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_223),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_156),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_264),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_181),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_156),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_177),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_172),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_172),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_204),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_204),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_226),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_285),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_175),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_226),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_281),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_185),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_281),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_176),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_276),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_276),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_185),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_193),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_211),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_245),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_212),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_239),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_264),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_164),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_222),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_234),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_237),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_164),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_198),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_242),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_287),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_248),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_198),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_249),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_256),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_205),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_285),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_321),
.B(n_277),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_356),
.B(n_154),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_321),
.B(n_277),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_299),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_331),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_354),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_317),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_320),
.B(n_154),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_326),
.B(n_259),
.Y(n_380)
);

INVxp33_ASAP7_75t_SL g381 ( 
.A(n_297),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_309),
.A2(n_235),
.B1(n_257),
.B2(n_261),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_356),
.B(n_206),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_317),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_322),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_322),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_320),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_323),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_323),
.Y(n_389)
);

AND3x1_ASAP7_75t_L g390 ( 
.A(n_349),
.B(n_266),
.C(n_260),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_307),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_328),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_328),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_298),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_315),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_298),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_301),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_296),
.B(n_206),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_296),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_R g400 ( 
.A(n_302),
.B(n_205),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_301),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_296),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_296),
.B(n_267),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_300),
.B(n_267),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_358),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_300),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_304),
.Y(n_407)
);

NAND2xp33_ASAP7_75t_L g408 ( 
.A(n_303),
.B(n_168),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_304),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_300),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_305),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_300),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_305),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_307),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_308),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_326),
.B(n_272),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_316),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_306),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_306),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_326),
.B(n_272),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_316),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_352),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_310),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_352),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_365),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_314),
.B(n_225),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_319),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_353),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_333),
.B(n_155),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_353),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_324),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_343),
.B(n_160),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_365),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_313),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_348),
.Y(n_435)
);

AND2x6_ASAP7_75t_L g436 ( 
.A(n_333),
.B(n_184),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_329),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_318),
.A2(n_240),
.B1(n_168),
.B2(n_171),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_342),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_329),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_426),
.B(n_358),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_391),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_391),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_394),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_394),
.Y(n_445)
);

INVxp67_ASAP7_75t_SL g446 ( 
.A(n_414),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_396),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_396),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_391),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_397),
.B(n_333),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_391),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_397),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_380),
.B(n_357),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_401),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_417),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_401),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_400),
.B(n_362),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_417),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_407),
.Y(n_459)
);

AO21x2_ASAP7_75t_L g460 ( 
.A1(n_432),
.A2(n_187),
.B(n_179),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_387),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_429),
.A2(n_311),
.B1(n_357),
.B2(n_275),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_425),
.Y(n_463)
);

AO21x2_ASAP7_75t_L g464 ( 
.A1(n_407),
.A2(n_191),
.B(n_189),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_409),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_406),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_425),
.Y(n_467)
);

OAI22xp33_ASAP7_75t_L g468 ( 
.A1(n_434),
.A2(n_362),
.B1(n_195),
.B2(n_183),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_387),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_372),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_409),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_411),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_392),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_411),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_425),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_392),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_425),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_375),
.B(n_371),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_414),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_414),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_413),
.B(n_357),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_414),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_413),
.B(n_418),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_406),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_418),
.B(n_180),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_415),
.B(n_371),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_419),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_414),
.Y(n_488)
);

OAI21xp33_ASAP7_75t_SL g489 ( 
.A1(n_373),
.A2(n_383),
.B(n_380),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_414),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_423),
.B(n_312),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_425),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_419),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_421),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_378),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_378),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_384),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_372),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_384),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_398),
.B(n_287),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_421),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_406),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_427),
.B(n_216),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_374),
.B(n_349),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_406),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_429),
.B(n_182),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_429),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_425),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_421),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_421),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_431),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_385),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_433),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_433),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_421),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_433),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_433),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_429),
.B(n_192),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_421),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_433),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_374),
.B(n_350),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_433),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_399),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_399),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_377),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_406),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_377),
.B(n_216),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_379),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_416),
.B(n_350),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_406),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_416),
.B(n_330),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_398),
.B(n_184),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_435),
.B(n_312),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_385),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_416),
.A2(n_286),
.B1(n_274),
.B2(n_269),
.Y(n_535)
);

INVxp67_ASAP7_75t_SL g536 ( 
.A(n_410),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_386),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_398),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_408),
.B(n_312),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_416),
.B(n_330),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_405),
.B(n_231),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_398),
.B(n_287),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_402),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_410),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_412),
.Y(n_545)
);

OAI22xp33_ASAP7_75t_L g546 ( 
.A1(n_439),
.A2(n_282),
.B1(n_284),
.B2(n_186),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_386),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_405),
.B(n_231),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_376),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_420),
.B(n_190),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_388),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_393),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_388),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_393),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_376),
.B(n_312),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_420),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_389),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_410),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_410),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_381),
.B(n_327),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_438),
.B(n_327),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_403),
.B(n_287),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_379),
.B(n_207),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_389),
.Y(n_564)
);

INVxp33_ASAP7_75t_L g565 ( 
.A(n_382),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_410),
.Y(n_566)
);

AO21x2_ASAP7_75t_L g567 ( 
.A1(n_403),
.A2(n_217),
.B(n_213),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_410),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_403),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_395),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_403),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_382),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_440),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_390),
.B(n_268),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_422),
.B(n_325),
.Y(n_575)
);

OR2x6_ASAP7_75t_L g576 ( 
.A(n_420),
.B(n_219),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_422),
.B(n_334),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_436),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_404),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_404),
.B(n_420),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_440),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_379),
.B(n_268),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_379),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_404),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_424),
.B(n_336),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_424),
.B(n_346),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_SL g587 ( 
.A(n_428),
.B(n_278),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_428),
.B(n_332),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_525),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_441),
.B(n_278),
.Y(n_590)
);

NAND3xp33_ASAP7_75t_L g591 ( 
.A(n_462),
.B(n_173),
.C(n_159),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_470),
.B(n_279),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_538),
.B(n_556),
.Y(n_593)
);

NOR3xp33_ASAP7_75t_L g594 ( 
.A(n_503),
.B(n_430),
.C(n_359),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_504),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_578),
.B(n_184),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_538),
.B(n_404),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_556),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_583),
.B(n_436),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_583),
.B(n_436),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_578),
.B(n_209),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_442),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_444),
.B(n_436),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_575),
.B(n_351),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_577),
.B(n_363),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_569),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_444),
.B(n_436),
.Y(n_607)
);

OAI221xp5_ASAP7_75t_L g608 ( 
.A1(n_535),
.A2(n_430),
.B1(n_238),
.B2(n_236),
.C(n_251),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_464),
.A2(n_460),
.B1(n_567),
.B2(n_447),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_445),
.B(n_436),
.Y(n_610)
);

O2A1O1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_489),
.A2(n_359),
.B(n_355),
.C(n_360),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_578),
.B(n_209),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_549),
.B(n_367),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_445),
.B(n_436),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_578),
.B(n_209),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_489),
.A2(n_279),
.B1(n_370),
.B2(n_208),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_SL g617 ( 
.A(n_511),
.B(n_235),
.Y(n_617)
);

OAI22x1_ASAP7_75t_SL g618 ( 
.A1(n_572),
.A2(n_261),
.B1(n_257),
.B2(n_171),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_549),
.B(n_355),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_470),
.B(n_165),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_498),
.B(n_165),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_SL g622 ( 
.A1(n_527),
.A2(n_289),
.B1(n_250),
.B2(n_243),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_498),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_507),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_570),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_582),
.B(n_166),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_584),
.B(n_209),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_485),
.B(n_561),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_442),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_574),
.B(n_166),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_569),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_541),
.B(n_360),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_SL g633 ( 
.A1(n_565),
.A2(n_227),
.B1(n_224),
.B2(n_265),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_447),
.B(n_440),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_448),
.B(n_437),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_507),
.A2(n_210),
.B1(n_194),
.B2(n_196),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_448),
.B(n_452),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_584),
.B(n_209),
.Y(n_638)
);

NAND3xp33_ASAP7_75t_L g639 ( 
.A(n_587),
.B(n_255),
.C(n_221),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_571),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_464),
.A2(n_287),
.B1(n_291),
.B2(n_285),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_464),
.A2(n_287),
.B1(n_291),
.B2(n_368),
.Y(n_642)
);

OAI221xp5_ASAP7_75t_L g643 ( 
.A1(n_450),
.A2(n_361),
.B1(n_369),
.B2(n_368),
.C(n_366),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_452),
.B(n_437),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_454),
.B(n_167),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_454),
.B(n_456),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_456),
.B(n_197),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_459),
.B(n_200),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_459),
.B(n_215),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_465),
.B(n_218),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_571),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_443),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_443),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_504),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_453),
.B(n_361),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_465),
.B(n_220),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_471),
.B(n_472),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_471),
.B(n_472),
.Y(n_658)
);

BUFx5_ASAP7_75t_L g659 ( 
.A(n_532),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_474),
.B(n_228),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_487),
.B(n_229),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_443),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_521),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_487),
.B(n_230),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_449),
.Y(n_665)
);

BUFx5_ASAP7_75t_L g666 ( 
.A(n_532),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_579),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_521),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_464),
.A2(n_291),
.B1(n_366),
.B2(n_364),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_493),
.B(n_232),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_449),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_528),
.Y(n_672)
);

NOR2x1_ASAP7_75t_L g673 ( 
.A(n_491),
.B(n_364),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_580),
.B(n_291),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_483),
.B(n_233),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_580),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_449),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_518),
.B(n_291),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_531),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_468),
.B(n_167),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_518),
.B(n_291),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_460),
.A2(n_291),
.B1(n_369),
.B2(n_290),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_450),
.B(n_241),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_529),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_451),
.Y(n_685)
);

BUFx8_ASAP7_75t_L g686 ( 
.A(n_588),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_481),
.B(n_247),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_481),
.B(n_252),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_531),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_495),
.B(n_253),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_451),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_496),
.B(n_262),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_528),
.Y(n_693)
);

OAI22xp5_ASAP7_75t_L g694 ( 
.A1(n_528),
.A2(n_170),
.B1(n_271),
.B2(n_294),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_518),
.B(n_500),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_455),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_496),
.B(n_263),
.Y(n_697)
);

NAND2x1p5_ASAP7_75t_L g698 ( 
.A(n_529),
.B(n_332),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_585),
.B(n_586),
.Y(n_699)
);

NOR3xp33_ASAP7_75t_L g700 ( 
.A(n_548),
.B(n_203),
.C(n_178),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_497),
.B(n_270),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_550),
.B(n_170),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_540),
.Y(n_703)
);

INVx8_ASAP7_75t_L g704 ( 
.A(n_576),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_457),
.B(n_188),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_540),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_455),
.Y(n_707)
);

BUFx12f_ASAP7_75t_SL g708 ( 
.A(n_576),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_497),
.B(n_288),
.Y(n_709)
);

NAND2xp33_ASAP7_75t_L g710 ( 
.A(n_532),
.B(n_280),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_560),
.B(n_347),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_588),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_499),
.B(n_295),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_518),
.B(n_283),
.Y(n_714)
);

INVx8_ASAP7_75t_L g715 ( 
.A(n_576),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_L g716 ( 
.A(n_532),
.B(n_292),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_499),
.B(n_293),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_L g718 ( 
.A1(n_576),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_512),
.B(n_271),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_512),
.B(n_294),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_534),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_539),
.A2(n_295),
.B1(n_244),
.B2(n_344),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_506),
.A2(n_347),
.B1(n_345),
.B2(n_344),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_534),
.B(n_345),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_537),
.B(n_0),
.Y(n_725)
);

O2A1O1Ixp5_ASAP7_75t_L g726 ( 
.A1(n_500),
.A2(n_341),
.B(n_340),
.C(n_339),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_511),
.B(n_341),
.Y(n_727)
);

NOR2xp67_ASAP7_75t_L g728 ( 
.A(n_533),
.B(n_111),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_511),
.Y(n_729)
);

O2A1O1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_542),
.A2(n_562),
.B(n_564),
.C(n_547),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_542),
.B(n_339),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_537),
.B(n_338),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_563),
.B(n_338),
.Y(n_733)
);

O2A1O1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_562),
.A2(n_337),
.B(n_335),
.C(n_3),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_547),
.Y(n_735)
);

OR2x6_ASAP7_75t_L g736 ( 
.A(n_478),
.B(n_337),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_563),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_551),
.B(n_335),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_551),
.B(n_0),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_563),
.B(n_147),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_553),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_553),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_563),
.B(n_146),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_557),
.B(n_123),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_SL g745 ( 
.A1(n_511),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_557),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_564),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_458),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_676),
.B(n_460),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_613),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_699),
.B(n_486),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_628),
.B(n_460),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_625),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_628),
.B(n_573),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_658),
.B(n_637),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_606),
.Y(n_756)
);

BUFx8_ASAP7_75t_L g757 ( 
.A(n_589),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_658),
.B(n_573),
.Y(n_758)
);

INVx5_ASAP7_75t_L g759 ( 
.A(n_672),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_631),
.Y(n_760)
);

NOR3xp33_ASAP7_75t_SL g761 ( 
.A(n_590),
.B(n_546),
.C(n_680),
.Y(n_761)
);

INVx4_ASAP7_75t_L g762 ( 
.A(n_624),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_624),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_646),
.B(n_573),
.Y(n_764)
);

NOR3xp33_ASAP7_75t_SL g765 ( 
.A(n_590),
.B(n_555),
.C(n_5),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_699),
.B(n_514),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_729),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_640),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_693),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_651),
.Y(n_770)
);

OR2x6_ASAP7_75t_L g771 ( 
.A(n_704),
.B(n_566),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_729),
.Y(n_772)
);

AND2x2_ASAP7_75t_SL g773 ( 
.A(n_617),
.B(n_566),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_657),
.B(n_581),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_667),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_727),
.B(n_479),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_696),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_684),
.A2(n_567),
.B1(n_446),
.B2(n_536),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_686),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_679),
.A2(n_567),
.B1(n_544),
.B2(n_532),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_595),
.B(n_566),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_689),
.A2(n_706),
.B1(n_703),
.B2(n_702),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_721),
.Y(n_783)
);

CKINVDCx16_ASAP7_75t_R g784 ( 
.A(n_604),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_735),
.B(n_581),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_654),
.B(n_567),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_702),
.A2(n_532),
.B1(n_475),
.B2(n_513),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_592),
.B(n_479),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_741),
.B(n_581),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_742),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_707),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_686),
.Y(n_792)
);

NAND2x1_ASAP7_75t_SL g793 ( 
.A(n_680),
.B(n_526),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_672),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_695),
.A2(n_593),
.B(n_597),
.Y(n_795)
);

OAI22xp33_ASAP7_75t_L g796 ( 
.A1(n_616),
.A2(n_479),
.B1(n_480),
.B2(n_482),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_736),
.Y(n_797)
);

BUFx2_ASAP7_75t_SL g798 ( 
.A(n_623),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_746),
.Y(n_799)
);

NOR2xp67_ASAP7_75t_L g800 ( 
.A(n_639),
.B(n_526),
.Y(n_800)
);

INVx6_ASAP7_75t_L g801 ( 
.A(n_704),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_748),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_704),
.B(n_530),
.Y(n_803)
);

BUFx12f_ASAP7_75t_L g804 ( 
.A(n_619),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_598),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_605),
.B(n_514),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_737),
.A2(n_532),
.B1(n_517),
.B2(n_477),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_693),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_R g809 ( 
.A(n_708),
.B(n_526),
.Y(n_809)
);

INVx5_ASAP7_75t_L g810 ( 
.A(n_715),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_682),
.A2(n_552),
.B1(n_554),
.B2(n_501),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_623),
.B(n_514),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_632),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_715),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_711),
.B(n_480),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_663),
.B(n_480),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_602),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_695),
.A2(n_482),
.B(n_488),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_635),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_668),
.B(n_482),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_712),
.B(n_488),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_736),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_644),
.Y(n_823)
);

AND2x6_ASAP7_75t_SL g824 ( 
.A(n_630),
.B(n_8),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_747),
.B(n_488),
.Y(n_825)
);

NOR3xp33_ASAP7_75t_L g826 ( 
.A(n_626),
.B(n_568),
.C(n_558),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_736),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_655),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_698),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_682),
.A2(n_552),
.B1(n_554),
.B2(n_523),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_730),
.B(n_490),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_731),
.B(n_490),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_705),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_629),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_698),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_630),
.A2(n_475),
.B1(n_467),
.B2(n_477),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_634),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_718),
.B(n_490),
.Y(n_838)
);

NAND3xp33_ASAP7_75t_SL g839 ( 
.A(n_700),
.B(n_722),
.C(n_745),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_652),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_718),
.B(n_494),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_641),
.A2(n_669),
.B1(n_642),
.B2(n_609),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_724),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_731),
.B(n_494),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_732),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_653),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_611),
.B(n_494),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_719),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_725),
.B(n_501),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_662),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_725),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_665),
.Y(n_852)
);

NAND2xp33_ASAP7_75t_L g853 ( 
.A(n_659),
.B(n_466),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_671),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_738),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_673),
.Y(n_856)
);

NOR3xp33_ASAP7_75t_SL g857 ( 
.A(n_633),
.B(n_8),
.C(n_9),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_739),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_739),
.B(n_520),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_677),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_594),
.B(n_733),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_733),
.B(n_568),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_685),
.Y(n_863)
);

OAI21xp33_ASAP7_75t_L g864 ( 
.A1(n_620),
.A2(n_552),
.B(n_554),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_720),
.Y(n_865)
);

NAND2xp33_ASAP7_75t_SL g866 ( 
.A(n_740),
.B(n_466),
.Y(n_866)
);

AO22x1_ASAP7_75t_L g867 ( 
.A1(n_621),
.A2(n_520),
.B1(n_510),
.B2(n_515),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_691),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_715),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_645),
.A2(n_713),
.B(n_621),
.C(n_609),
.Y(n_870)
);

INVx5_ASAP7_75t_L g871 ( 
.A(n_659),
.Y(n_871)
);

OR2x6_ASAP7_75t_L g872 ( 
.A(n_740),
.B(n_530),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_674),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_674),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_714),
.B(n_568),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_683),
.B(n_510),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_687),
.A2(n_467),
.B1(n_477),
.B2(n_492),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_726),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_688),
.B(n_669),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_622),
.B(n_515),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_675),
.B(n_645),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_647),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_659),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_618),
.Y(n_884)
);

INVx4_ASAP7_75t_L g885 ( 
.A(n_659),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_723),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_678),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_694),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_648),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_713),
.B(n_509),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_636),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_603),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_607),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_743),
.B(n_568),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_649),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_650),
.Y(n_896)
);

NAND2x2_ASAP7_75t_L g897 ( 
.A(n_656),
.B(n_9),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_610),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_678),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_681),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_591),
.B(n_516),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_744),
.B(n_519),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_681),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_660),
.Y(n_904)
);

BUFx2_ASAP7_75t_L g905 ( 
.A(n_661),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_614),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_599),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_627),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_642),
.B(n_519),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_664),
.B(n_522),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_670),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_627),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_600),
.Y(n_913)
);

INVx4_ASAP7_75t_L g914 ( 
.A(n_659),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_638),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_638),
.Y(n_916)
);

NOR3xp33_ASAP7_75t_SL g917 ( 
.A(n_643),
.B(n_10),
.C(n_13),
.Y(n_917)
);

OR2x6_ASAP7_75t_L g918 ( 
.A(n_734),
.B(n_530),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_666),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_690),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_870),
.A2(n_751),
.B(n_858),
.C(n_851),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_810),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_882),
.B(n_692),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_760),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_882),
.B(n_709),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_813),
.B(n_717),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_756),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_768),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_SL g929 ( 
.A(n_842),
.B(n_728),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_755),
.B(n_697),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_755),
.B(n_701),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_881),
.A2(n_608),
.B(n_615),
.C(n_612),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_881),
.B(n_601),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_871),
.A2(n_516),
.B(n_596),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_761),
.A2(n_920),
.B(n_842),
.C(n_895),
.Y(n_935)
);

CKINVDCx6p67_ASAP7_75t_R g936 ( 
.A(n_753),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_895),
.A2(n_615),
.B(n_612),
.C(n_601),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_848),
.B(n_596),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_871),
.A2(n_716),
.B(n_710),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_752),
.A2(n_463),
.B1(n_477),
.B2(n_492),
.Y(n_940)
);

INVx6_ASAP7_75t_L g941 ( 
.A(n_757),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_871),
.A2(n_914),
.B(n_885),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_848),
.B(n_508),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_752),
.A2(n_754),
.B1(n_758),
.B2(n_879),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_879),
.A2(n_513),
.B(n_492),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_853),
.A2(n_502),
.B(n_559),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_813),
.B(n_524),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_766),
.B(n_526),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_843),
.B(n_558),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_814),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_770),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_759),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_819),
.B(n_558),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_775),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_845),
.B(n_508),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_783),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_833),
.A2(n_896),
.B(n_904),
.C(n_865),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_823),
.B(n_508),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_833),
.B(n_513),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_866),
.A2(n_517),
.B(n_524),
.C(n_545),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_861),
.A2(n_782),
.B(n_795),
.C(n_874),
.Y(n_961)
);

AND2x2_ASAP7_75t_SL g962 ( 
.A(n_773),
.B(n_523),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_861),
.A2(n_517),
.B(n_543),
.C(n_469),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_795),
.A2(n_484),
.B(n_559),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_814),
.B(n_517),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_790),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_905),
.B(n_559),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_R g968 ( 
.A(n_767),
.B(n_772),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_840),
.Y(n_969)
);

INVxp67_ASAP7_75t_SL g970 ( 
.A(n_808),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_784),
.B(n_476),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_750),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_804),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_889),
.B(n_505),
.Y(n_974)
);

INVx6_ASAP7_75t_L g975 ( 
.A(n_757),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_799),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_797),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_SL g978 ( 
.A1(n_891),
.A2(n_888),
.B1(n_798),
.B2(n_911),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_855),
.B(n_476),
.Y(n_979)
);

OA22x2_ASAP7_75t_L g980 ( 
.A1(n_827),
.A2(n_10),
.B1(n_16),
.B2(n_18),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_759),
.Y(n_981)
);

CKINVDCx6p67_ASAP7_75t_R g982 ( 
.A(n_779),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_837),
.B(n_473),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_822),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_828),
.B(n_473),
.Y(n_985)
);

NAND2xp33_ASAP7_75t_SL g986 ( 
.A(n_814),
.B(n_505),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_846),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_792),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_869),
.Y(n_989)
);

NAND2x1p5_ASAP7_75t_L g990 ( 
.A(n_810),
.B(n_505),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_763),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_856),
.B(n_505),
.Y(n_992)
);

BUFx4_ASAP7_75t_SL g993 ( 
.A(n_824),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_846),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_806),
.B(n_461),
.Y(n_995)
);

NOR3xp33_ASAP7_75t_SL g996 ( 
.A(n_884),
.B(n_16),
.C(n_20),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_869),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_758),
.A2(n_461),
.B1(n_505),
.B2(n_484),
.Y(n_998)
);

INVx1_ASAP7_75t_SL g999 ( 
.A(n_793),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_821),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_838),
.A2(n_23),
.B(n_24),
.C(n_27),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_794),
.Y(n_1002)
);

CKINVDCx11_ASAP7_75t_R g1003 ( 
.A(n_897),
.Y(n_1003)
);

INVx1_ASAP7_75t_SL g1004 ( 
.A(n_786),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_869),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_805),
.B(n_812),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_763),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_909),
.A2(n_666),
.B(n_484),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_781),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_810),
.Y(n_1010)
);

BUFx12f_ASAP7_75t_L g1011 ( 
.A(n_801),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_873),
.A2(n_484),
.B(n_466),
.C(n_33),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_809),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_SL g1014 ( 
.A(n_765),
.B(n_28),
.C(n_31),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_883),
.A2(n_484),
.B(n_466),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_749),
.A2(n_28),
.B1(n_33),
.B2(n_37),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_764),
.B(n_61),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_786),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_887),
.A2(n_39),
.B(n_47),
.C(n_48),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_841),
.A2(n_48),
.B(n_49),
.C(n_62),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_835),
.B(n_49),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_919),
.A2(n_70),
.B(n_81),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_777),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_794),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_762),
.B(n_769),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_899),
.A2(n_900),
.B(n_903),
.C(n_886),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_808),
.B(n_764),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_875),
.A2(n_862),
.B1(n_829),
.B2(n_880),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_769),
.B(n_816),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_749),
.A2(n_901),
.B(n_908),
.C(n_916),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_857),
.B(n_875),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_801),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_788),
.A2(n_815),
.B(n_776),
.C(n_820),
.Y(n_1033)
);

NOR3xp33_ASAP7_75t_L g1034 ( 
.A(n_910),
.B(n_796),
.C(n_876),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_801),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_917),
.B(n_862),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_810),
.B(n_894),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_785),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_894),
.A2(n_800),
.B1(n_826),
.B2(n_872),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_913),
.B(n_825),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_771),
.B(n_803),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_791),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_876),
.A2(n_909),
.B(n_774),
.Y(n_1043)
);

NAND3xp33_ASAP7_75t_SL g1044 ( 
.A(n_826),
.B(n_780),
.C(n_890),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_774),
.A2(n_872),
.B(n_902),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_872),
.A2(n_912),
.B1(n_913),
.B2(n_907),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_830),
.A2(n_849),
.B1(n_859),
.B2(n_890),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_913),
.B(n_825),
.Y(n_1048)
);

AOI21xp33_ASAP7_75t_L g1049 ( 
.A1(n_921),
.A2(n_847),
.B(n_864),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_1045),
.A2(n_902),
.B(n_831),
.Y(n_1050)
);

AO31x2_ASAP7_75t_L g1051 ( 
.A1(n_944),
.A2(n_811),
.A3(n_831),
.B(n_878),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_929),
.A2(n_1043),
.B(n_942),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_SL g1053 ( 
.A1(n_1020),
.A2(n_818),
.B(n_785),
.Y(n_1053)
);

NAND3xp33_ASAP7_75t_L g1054 ( 
.A(n_923),
.B(n_778),
.C(n_836),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_944),
.A2(n_811),
.B(n_906),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_924),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_971),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_968),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_928),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_935),
.A2(n_844),
.B(n_832),
.Y(n_1060)
);

OA22x2_ASAP7_75t_L g1061 ( 
.A1(n_972),
.A2(n_918),
.B1(n_771),
.B2(n_807),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_925),
.B(n_850),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_1041),
.B(n_771),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1044),
.A2(n_832),
.B(n_844),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_964),
.A2(n_789),
.B(n_877),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_995),
.A2(n_789),
.B(n_867),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_978),
.A2(n_898),
.B1(n_893),
.B2(n_892),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_926),
.B(n_834),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_957),
.B(n_860),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1000),
.B(n_863),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_951),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1038),
.B(n_915),
.Y(n_1072)
);

OAI22x1_ASAP7_75t_L g1073 ( 
.A1(n_1031),
.A2(n_787),
.B1(n_868),
.B2(n_817),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1047),
.A2(n_803),
.B(n_918),
.Y(n_1074)
);

NOR2x1_ASAP7_75t_SL g1075 ( 
.A(n_922),
.B(n_852),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_1041),
.B(n_854),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_1015),
.A2(n_802),
.B(n_946),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_933),
.B(n_1040),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_938),
.B(n_1006),
.Y(n_1079)
);

OA21x2_ASAP7_75t_L g1080 ( 
.A1(n_945),
.A2(n_1030),
.B(n_1008),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_936),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_954),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_962),
.B(n_1004),
.Y(n_1083)
);

AND2x6_ASAP7_75t_SL g1084 ( 
.A(n_1021),
.B(n_993),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1004),
.B(n_1009),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_933),
.A2(n_961),
.B1(n_1018),
.B2(n_1028),
.Y(n_1086)
);

OAI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_956),
.A2(n_976),
.B(n_966),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1036),
.B(n_947),
.Y(n_1088)
);

NOR2xp67_ASAP7_75t_L g1089 ( 
.A(n_1011),
.B(n_927),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1048),
.B(n_1027),
.Y(n_1090)
);

NAND2x1p5_ASAP7_75t_L g1091 ( 
.A(n_922),
.B(n_1010),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_SL g1092 ( 
.A1(n_937),
.A2(n_932),
.B(n_1017),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1026),
.B(n_979),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_998),
.A2(n_940),
.B(n_934),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_943),
.B(n_983),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_SL g1096 ( 
.A1(n_1001),
.A2(n_1033),
.B(n_1046),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_967),
.B(n_959),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_1010),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1023),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1013),
.B(n_991),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1034),
.A2(n_1017),
.B(n_963),
.Y(n_1101)
);

AOI211x1_ASAP7_75t_L g1102 ( 
.A1(n_1014),
.A2(n_1016),
.B(n_985),
.C(n_1037),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_SL g1103 ( 
.A1(n_1039),
.A2(n_948),
.B(n_1012),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_958),
.A2(n_953),
.B(n_990),
.Y(n_1104)
);

NOR2xp67_ASAP7_75t_L g1105 ( 
.A(n_973),
.B(n_1032),
.Y(n_1105)
);

NAND3xp33_ASAP7_75t_L g1106 ( 
.A(n_1019),
.B(n_1016),
.C(n_996),
.Y(n_1106)
);

AO31x2_ASAP7_75t_L g1107 ( 
.A1(n_960),
.A2(n_953),
.A3(n_955),
.B(n_949),
.Y(n_1107)
);

OAI21xp33_ASAP7_75t_L g1108 ( 
.A1(n_980),
.A2(n_1029),
.B(n_988),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1002),
.B(n_1024),
.Y(n_1109)
);

AO31x2_ASAP7_75t_L g1110 ( 
.A1(n_974),
.A2(n_992),
.A3(n_1022),
.B(n_994),
.Y(n_1110)
);

AO21x1_ASAP7_75t_L g1111 ( 
.A1(n_986),
.A2(n_970),
.B(n_1025),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_977),
.Y(n_1112)
);

OAI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_980),
.A2(n_1042),
.B(n_999),
.Y(n_1113)
);

NOR2xp67_ASAP7_75t_L g1114 ( 
.A(n_969),
.B(n_987),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_952),
.A2(n_981),
.B(n_1024),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_981),
.A2(n_965),
.B(n_1007),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_R g1117 ( 
.A(n_1035),
.B(n_1005),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_965),
.A2(n_989),
.B(n_950),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_950),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_950),
.B(n_989),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_989),
.Y(n_1121)
);

AO31x2_ASAP7_75t_L g1122 ( 
.A1(n_984),
.A2(n_1003),
.A3(n_997),
.B(n_1005),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_997),
.B(n_1005),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1035),
.B(n_982),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_1035),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_941),
.A2(n_842),
.B1(n_870),
.B2(n_755),
.Y(n_1126)
);

AO21x1_ASAP7_75t_L g1127 ( 
.A1(n_941),
.A2(n_929),
.B(n_842),
.Y(n_1127)
);

AO22x2_ASAP7_75t_L g1128 ( 
.A1(n_975),
.A2(n_1016),
.B1(n_842),
.B2(n_839),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_975),
.A2(n_751),
.B(n_699),
.C(n_628),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_964),
.A2(n_818),
.B(n_939),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_964),
.A2(n_818),
.B(n_939),
.Y(n_1131)
);

BUFx12f_ASAP7_75t_L g1132 ( 
.A(n_1003),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_924),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1045),
.A2(n_871),
.B(n_929),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_968),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_923),
.B(n_699),
.Y(n_1136)
);

AO21x1_ASAP7_75t_L g1137 ( 
.A1(n_929),
.A2(n_842),
.B(n_866),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1045),
.A2(n_871),
.B(n_929),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_944),
.A2(n_870),
.A3(n_1047),
.B(n_1030),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_924),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_964),
.A2(n_818),
.B(n_939),
.Y(n_1141)
);

AOI21xp33_ASAP7_75t_L g1142 ( 
.A1(n_921),
.A2(n_699),
.B(n_751),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_964),
.A2(n_818),
.B(n_939),
.Y(n_1143)
);

NOR3xp33_ASAP7_75t_SL g1144 ( 
.A(n_1014),
.B(n_884),
.C(n_572),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1045),
.A2(n_871),
.B(n_929),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_964),
.A2(n_818),
.B(n_939),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1045),
.A2(n_870),
.B(n_944),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_930),
.B(n_931),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_924),
.Y(n_1149)
);

NAND2x1p5_ASAP7_75t_L g1150 ( 
.A(n_922),
.B(n_810),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_924),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_923),
.B(n_604),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1045),
.A2(n_870),
.B(n_944),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_935),
.A2(n_751),
.B(n_699),
.C(n_628),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_SL g1155 ( 
.A(n_988),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_930),
.B(n_931),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_930),
.B(n_931),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1045),
.A2(n_870),
.B(n_944),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_930),
.B(n_931),
.Y(n_1159)
);

NAND3x1_ASAP7_75t_L g1160 ( 
.A(n_1021),
.B(n_751),
.C(n_699),
.Y(n_1160)
);

OA21x2_ASAP7_75t_L g1161 ( 
.A1(n_1045),
.A2(n_945),
.B(n_1043),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_1011),
.Y(n_1162)
);

OAI21xp33_ASAP7_75t_SL g1163 ( 
.A1(n_930),
.A2(n_842),
.B(n_755),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1045),
.A2(n_871),
.B(n_929),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_924),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_SL g1166 ( 
.A1(n_1020),
.A2(n_1001),
.B(n_1033),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_930),
.B(n_931),
.Y(n_1167)
);

BUFx4_ASAP7_75t_SL g1168 ( 
.A(n_988),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_924),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1045),
.A2(n_871),
.B(n_929),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1045),
.A2(n_870),
.B(n_944),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1045),
.A2(n_870),
.B(n_944),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_924),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_922),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_930),
.B(n_931),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1045),
.A2(n_871),
.B(n_929),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1136),
.A2(n_1154),
.B(n_1142),
.C(n_1148),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1138),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1164),
.A2(n_1176),
.B(n_1170),
.Y(n_1179)
);

XNOR2xp5_ASAP7_75t_L g1180 ( 
.A(n_1160),
.B(n_1058),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1082),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1077),
.A2(n_1131),
.B(n_1130),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1133),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1141),
.A2(n_1146),
.B(n_1143),
.Y(n_1184)
);

AO21x2_ASAP7_75t_L g1185 ( 
.A1(n_1052),
.A2(n_1074),
.B(n_1147),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1168),
.Y(n_1186)
);

OAI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1157),
.A2(n_1175),
.B1(n_1159),
.B2(n_1156),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1156),
.B(n_1167),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1149),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1167),
.B(n_1152),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1088),
.B(n_1068),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1165),
.Y(n_1192)
);

OAI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1106),
.A2(n_1079),
.B1(n_1142),
.B2(n_1126),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1065),
.A2(n_1094),
.B(n_1104),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_SL g1195 ( 
.A1(n_1127),
.A2(n_1096),
.B(n_1166),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1062),
.B(n_1057),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1129),
.B(n_1078),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1073),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1169),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1097),
.A2(n_1067),
.B1(n_1069),
.B2(n_1061),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1085),
.Y(n_1201)
);

CKINVDCx16_ASAP7_75t_R g1202 ( 
.A(n_1155),
.Y(n_1202)
);

AO21x2_ASAP7_75t_L g1203 ( 
.A1(n_1147),
.A2(n_1171),
.B(n_1153),
.Y(n_1203)
);

AO32x2_ASAP7_75t_L g1204 ( 
.A1(n_1126),
.A2(n_1086),
.A3(n_1139),
.B1(n_1172),
.B2(n_1171),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1078),
.B(n_1090),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1128),
.A2(n_1108),
.B1(n_1086),
.B2(n_1137),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1053),
.A2(n_1101),
.B(n_1115),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1056),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1092),
.A2(n_1153),
.B(n_1172),
.Y(n_1209)
);

INVx4_ASAP7_75t_SL g1210 ( 
.A(n_1122),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1059),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1071),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1140),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1128),
.A2(n_1113),
.B1(n_1054),
.B2(n_1158),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1101),
.A2(n_1158),
.B(n_1055),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1151),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1055),
.A2(n_1066),
.B(n_1060),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1144),
.A2(n_1063),
.B1(n_1155),
.B2(n_1100),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1163),
.A2(n_1049),
.B1(n_1061),
.B2(n_1087),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1049),
.A2(n_1064),
.B1(n_1060),
.B2(n_1090),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1173),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1063),
.A2(n_1076),
.B1(n_1135),
.B2(n_1089),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1116),
.B(n_1076),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1093),
.A2(n_1111),
.A3(n_1075),
.B(n_1095),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1064),
.A2(n_1161),
.B(n_1093),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1072),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1099),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1080),
.A2(n_1109),
.B(n_1070),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1150),
.A2(n_1080),
.B(n_1091),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1084),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_1112),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1098),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1174),
.A2(n_1118),
.B(n_1083),
.Y(n_1233)
);

AOI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1114),
.A2(n_1120),
.B(n_1123),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1139),
.A2(n_1105),
.B(n_1102),
.C(n_1174),
.Y(n_1235)
);

OA21x2_ASAP7_75t_L g1236 ( 
.A1(n_1051),
.A2(n_1107),
.B(n_1110),
.Y(n_1236)
);

AOI22x1_ASAP7_75t_L g1237 ( 
.A1(n_1119),
.A2(n_1125),
.B1(n_1121),
.B2(n_1162),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_1051),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1162),
.A2(n_1132),
.B1(n_1081),
.B2(n_1120),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1123),
.B(n_1124),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1162),
.A2(n_1124),
.B1(n_1121),
.B2(n_1122),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1122),
.B(n_1117),
.Y(n_1242)
);

O2A1O1Ixp33_ASAP7_75t_SL g1243 ( 
.A1(n_1107),
.A2(n_1154),
.B(n_870),
.C(n_842),
.Y(n_1243)
);

OR2x6_ASAP7_75t_L g1244 ( 
.A(n_1061),
.B(n_1103),
.Y(n_1244)
);

OR2x6_ASAP7_75t_L g1245 ( 
.A(n_1061),
.B(n_1103),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1057),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1136),
.A2(n_699),
.B1(n_1142),
.B2(n_751),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1136),
.B(n_1148),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1082),
.Y(n_1249)
);

OA21x2_ASAP7_75t_L g1250 ( 
.A1(n_1147),
.A2(n_1158),
.B(n_1153),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1082),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1136),
.B(n_699),
.Y(n_1252)
);

AOI221xp5_ASAP7_75t_L g1253 ( 
.A1(n_1136),
.A2(n_699),
.B1(n_751),
.B2(n_1142),
.C(n_1154),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1057),
.Y(n_1254)
);

OA21x2_ASAP7_75t_L g1255 ( 
.A1(n_1147),
.A2(n_1158),
.B(n_1153),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1082),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1082),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1168),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1136),
.A2(n_699),
.B1(n_1142),
.B2(n_751),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1063),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1130),
.A2(n_1141),
.B(n_1131),
.Y(n_1261)
);

AOI22x1_ASAP7_75t_L g1262 ( 
.A1(n_1128),
.A2(n_858),
.B1(n_851),
.B2(n_1073),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1063),
.B(n_1041),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1130),
.A2(n_1141),
.B(n_1131),
.Y(n_1264)
);

AO21x2_ASAP7_75t_L g1265 ( 
.A1(n_1052),
.A2(n_1074),
.B(n_1176),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1058),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_SL g1267 ( 
.A1(n_1127),
.A2(n_1096),
.B(n_1166),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1137),
.A2(n_1073),
.A3(n_1050),
.B(n_1074),
.Y(n_1268)
);

AO21x2_ASAP7_75t_L g1269 ( 
.A1(n_1052),
.A2(n_1074),
.B(n_1176),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1138),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_SL g1271 ( 
.A1(n_1127),
.A2(n_1096),
.B(n_1166),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1130),
.A2(n_1141),
.B(n_1131),
.Y(n_1272)
);

AOI22x1_ASAP7_75t_L g1273 ( 
.A1(n_1128),
.A2(n_858),
.B1(n_851),
.B2(n_1073),
.Y(n_1273)
);

INVx4_ASAP7_75t_L g1274 ( 
.A(n_1162),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1136),
.B(n_1148),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1136),
.B(n_1148),
.Y(n_1276)
);

AO21x2_ASAP7_75t_L g1277 ( 
.A1(n_1052),
.A2(n_1074),
.B(n_1176),
.Y(n_1277)
);

AO21x2_ASAP7_75t_L g1278 ( 
.A1(n_1052),
.A2(n_1074),
.B(n_1176),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1130),
.A2(n_1141),
.B(n_1131),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_SL g1280 ( 
.A1(n_1127),
.A2(n_1096),
.B(n_1166),
.Y(n_1280)
);

AND2x6_ASAP7_75t_L g1281 ( 
.A(n_1067),
.B(n_1041),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1082),
.Y(n_1282)
);

NAND2x1p5_ASAP7_75t_L g1283 ( 
.A(n_1098),
.B(n_810),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1136),
.A2(n_1160),
.B1(n_699),
.B2(n_1157),
.Y(n_1284)
);

INVx8_ASAP7_75t_L g1285 ( 
.A(n_1155),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_1147),
.A2(n_1158),
.B(n_1153),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1112),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1136),
.A2(n_1160),
.B1(n_699),
.B2(n_1157),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_1168),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1082),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1130),
.A2(n_1141),
.B(n_1131),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1082),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1077),
.A2(n_1131),
.B(n_1130),
.Y(n_1293)
);

AOI21xp33_ASAP7_75t_L g1294 ( 
.A1(n_1136),
.A2(n_699),
.B(n_751),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1112),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1063),
.B(n_1041),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1082),
.Y(n_1297)
);

OA21x2_ASAP7_75t_L g1298 ( 
.A1(n_1147),
.A2(n_1158),
.B(n_1153),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1191),
.B(n_1190),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_SL g1300 ( 
.A1(n_1209),
.A2(n_1187),
.B(n_1253),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1246),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_SL g1302 ( 
.A1(n_1187),
.A2(n_1177),
.B(n_1284),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1178),
.A2(n_1270),
.B(n_1179),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1205),
.B(n_1188),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1254),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1252),
.A2(n_1247),
.B1(n_1259),
.B2(n_1275),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1287),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1201),
.B(n_1254),
.Y(n_1308)
);

NAND2xp33_ASAP7_75t_SL g1309 ( 
.A(n_1266),
.B(n_1248),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1201),
.B(n_1196),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1263),
.B(n_1296),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1213),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1193),
.B(n_1177),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1252),
.A2(n_1247),
.B1(n_1259),
.B2(n_1276),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1240),
.B(n_1214),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1203),
.A2(n_1298),
.B(n_1250),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1223),
.B(n_1260),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1208),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1193),
.B(n_1226),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1294),
.A2(n_1244),
.B1(n_1245),
.B2(n_1206),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1203),
.A2(n_1298),
.B(n_1250),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1288),
.A2(n_1200),
.B(n_1235),
.C(n_1197),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1244),
.A2(n_1245),
.B1(n_1206),
.B2(n_1214),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1199),
.B(n_1251),
.Y(n_1324)
);

O2A1O1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1235),
.A2(n_1271),
.B(n_1267),
.C(n_1195),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1251),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1223),
.B(n_1260),
.Y(n_1327)
);

INVx4_ASAP7_75t_L g1328 ( 
.A(n_1186),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1226),
.B(n_1220),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1211),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1256),
.B(n_1257),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1255),
.A2(n_1286),
.B(n_1185),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1256),
.Y(n_1333)
);

INVx4_ASAP7_75t_L g1334 ( 
.A(n_1186),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1232),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_SL g1336 ( 
.A1(n_1255),
.A2(n_1286),
.B(n_1180),
.Y(n_1336)
);

NOR2xp67_ASAP7_75t_L g1337 ( 
.A(n_1218),
.B(n_1222),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1231),
.B(n_1266),
.Y(n_1338)
);

AOI21x1_ASAP7_75t_SL g1339 ( 
.A1(n_1242),
.A2(n_1198),
.B(n_1238),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1286),
.A2(n_1185),
.B(n_1277),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1212),
.Y(n_1341)
);

OA21x2_ASAP7_75t_L g1342 ( 
.A1(n_1225),
.A2(n_1217),
.B(n_1194),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1257),
.B(n_1290),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1258),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1292),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1220),
.B(n_1219),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1280),
.A2(n_1243),
.B(n_1221),
.C(n_1216),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1219),
.A2(n_1239),
.B1(n_1241),
.B2(n_1183),
.Y(n_1348)
);

OA21x2_ASAP7_75t_L g1349 ( 
.A1(n_1217),
.A2(n_1194),
.B(n_1182),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1227),
.Y(n_1350)
);

BUFx5_ASAP7_75t_L g1351 ( 
.A(n_1281),
.Y(n_1351)
);

AOI21x1_ASAP7_75t_SL g1352 ( 
.A1(n_1210),
.A2(n_1273),
.B(n_1262),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_SL g1353 ( 
.A1(n_1274),
.A2(n_1283),
.B(n_1265),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1297),
.B(n_1181),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1297),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1293),
.A2(n_1207),
.B(n_1215),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1215),
.A2(n_1184),
.B(n_1261),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1189),
.Y(n_1358)
);

CKINVDCx6p67_ASAP7_75t_R g1359 ( 
.A(n_1202),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1192),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1249),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1232),
.B(n_1234),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_SL g1363 ( 
.A1(n_1274),
.A2(n_1283),
.B(n_1265),
.Y(n_1363)
);

AOI21x1_ASAP7_75t_SL g1364 ( 
.A1(n_1285),
.A2(n_1230),
.B(n_1224),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1282),
.B(n_1295),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1281),
.B(n_1233),
.Y(n_1366)
);

O2A1O1Ixp33_ASAP7_75t_L g1367 ( 
.A1(n_1269),
.A2(n_1278),
.B(n_1239),
.C(n_1289),
.Y(n_1367)
);

NOR2xp67_ASAP7_75t_L g1368 ( 
.A(n_1258),
.B(n_1230),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1285),
.A2(n_1237),
.B1(n_1204),
.B2(n_1236),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1224),
.B(n_1281),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1228),
.B(n_1224),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1281),
.A2(n_1236),
.B(n_1204),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1281),
.B(n_1229),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1184),
.A2(n_1272),
.B(n_1291),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1228),
.B(n_1268),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1268),
.B(n_1236),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1261),
.A2(n_1279),
.B(n_1264),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1191),
.B(n_1190),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_SL g1379 ( 
.A1(n_1209),
.A2(n_1154),
.B(n_842),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1187),
.B(n_1205),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1187),
.B(n_1205),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1191),
.B(n_1190),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_SL g1383 ( 
.A1(n_1197),
.A2(n_1242),
.B(n_1031),
.Y(n_1383)
);

O2A1O1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1294),
.A2(n_699),
.B(n_1154),
.C(n_1129),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1209),
.A2(n_1154),
.B(n_842),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1191),
.B(n_1190),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1223),
.B(n_1260),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1263),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1187),
.B(n_1205),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1191),
.B(n_1190),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1191),
.B(n_1190),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1308),
.B(n_1376),
.Y(n_1392)
);

OAI221xp5_ASAP7_75t_L g1393 ( 
.A1(n_1384),
.A2(n_1300),
.B1(n_1302),
.B2(n_1313),
.C(n_1306),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_L g1394 ( 
.A(n_1306),
.B(n_1314),
.C(n_1313),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1380),
.B(n_1381),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1318),
.B(n_1330),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1341),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1340),
.A2(n_1303),
.B(n_1374),
.Y(n_1398)
);

OR2x6_ASAP7_75t_L g1399 ( 
.A(n_1372),
.B(n_1303),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1323),
.A2(n_1314),
.B1(n_1320),
.B2(n_1337),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1373),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1350),
.Y(n_1402)
);

AO21x2_ASAP7_75t_L g1403 ( 
.A1(n_1332),
.A2(n_1316),
.B(n_1321),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1351),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1357),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1338),
.B(n_1299),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1317),
.B(n_1327),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1301),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1380),
.B(n_1381),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1370),
.B(n_1305),
.Y(n_1410)
);

INVxp67_ASAP7_75t_SL g1411 ( 
.A(n_1347),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1389),
.B(n_1329),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1375),
.B(n_1371),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1387),
.B(n_1370),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1389),
.B(n_1329),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1373),
.B(n_1342),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1342),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1369),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1319),
.B(n_1304),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1387),
.B(n_1336),
.Y(n_1420)
);

INVx4_ASAP7_75t_L g1421 ( 
.A(n_1362),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1319),
.B(n_1304),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1312),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1310),
.B(n_1315),
.Y(n_1424)
);

AO21x2_ASAP7_75t_L g1425 ( 
.A1(n_1379),
.A2(n_1385),
.B(n_1346),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1358),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1378),
.B(n_1391),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1346),
.B(n_1333),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1360),
.Y(n_1429)
);

OAI22x1_ASAP7_75t_L g1430 ( 
.A1(n_1366),
.A2(n_1362),
.B1(n_1361),
.B2(n_1356),
.Y(n_1430)
);

AO21x2_ASAP7_75t_L g1431 ( 
.A1(n_1367),
.A2(n_1320),
.B(n_1322),
.Y(n_1431)
);

AO21x2_ASAP7_75t_L g1432 ( 
.A1(n_1325),
.A2(n_1363),
.B(n_1353),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1345),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1349),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1355),
.B(n_1356),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_SL g1436 ( 
.A1(n_1348),
.A2(n_1307),
.B(n_1365),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1377),
.Y(n_1437)
);

NAND2xp33_ASAP7_75t_SL g1438 ( 
.A(n_1328),
.B(n_1334),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_1354),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1382),
.B(n_1386),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1351),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1390),
.B(n_1351),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_SL g1443 ( 
.A1(n_1326),
.A2(n_1343),
.B(n_1324),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1437),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1393),
.A2(n_1309),
.B(n_1383),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1412),
.B(n_1415),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1404),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1395),
.B(n_1388),
.Y(n_1448)
);

NAND3xp33_ASAP7_75t_L g1449 ( 
.A(n_1394),
.B(n_1331),
.C(n_1335),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1416),
.B(n_1351),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1393),
.A2(n_1351),
.B1(n_1359),
.B2(n_1388),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1392),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1441),
.B(n_1335),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1399),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1416),
.B(n_1311),
.Y(n_1455)
);

INVx3_ASAP7_75t_SL g1456 ( 
.A(n_1399),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1397),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1392),
.B(n_1339),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1402),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1435),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1410),
.B(n_1328),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1405),
.B(n_1368),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1405),
.B(n_1352),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1410),
.B(n_1418),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1405),
.B(n_1364),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1424),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1417),
.B(n_1344),
.Y(n_1467)
);

OAI322xp33_ASAP7_75t_L g1468 ( 
.A1(n_1446),
.A2(n_1395),
.A3(n_1409),
.B1(n_1394),
.B2(n_1415),
.C1(n_1412),
.C2(n_1422),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1447),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1457),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1445),
.A2(n_1425),
.B1(n_1431),
.B2(n_1411),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1457),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1450),
.B(n_1447),
.Y(n_1473)
);

AOI211xp5_ASAP7_75t_L g1474 ( 
.A1(n_1445),
.A2(n_1436),
.B(n_1409),
.C(n_1418),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1446),
.B(n_1466),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1452),
.Y(n_1476)
);

NAND2xp33_ASAP7_75t_R g1477 ( 
.A(n_1467),
.B(n_1420),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1452),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1451),
.A2(n_1400),
.B1(n_1425),
.B2(n_1431),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1451),
.A2(n_1425),
.B1(n_1431),
.B2(n_1399),
.Y(n_1480)
);

NAND3xp33_ASAP7_75t_L g1481 ( 
.A(n_1449),
.B(n_1436),
.C(n_1399),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1455),
.B(n_1450),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1448),
.B(n_1424),
.Y(n_1483)
);

OAI221xp5_ASAP7_75t_L g1484 ( 
.A1(n_1449),
.A2(n_1419),
.B1(n_1422),
.B2(n_1399),
.C(n_1411),
.Y(n_1484)
);

OAI222xp33_ASAP7_75t_L g1485 ( 
.A1(n_1461),
.A2(n_1399),
.B1(n_1420),
.B2(n_1419),
.C1(n_1442),
.C2(n_1428),
.Y(n_1485)
);

AOI222xp33_ASAP7_75t_L g1486 ( 
.A1(n_1448),
.A2(n_1406),
.B1(n_1428),
.B2(n_1439),
.C1(n_1440),
.C2(n_1427),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1455),
.B(n_1413),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_R g1488 ( 
.A(n_1467),
.B(n_1438),
.Y(n_1488)
);

NAND2xp33_ASAP7_75t_SL g1489 ( 
.A(n_1456),
.B(n_1432),
.Y(n_1489)
);

INVx4_ASAP7_75t_L g1490 ( 
.A(n_1453),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1450),
.B(n_1401),
.Y(n_1491)
);

AOI221xp5_ASAP7_75t_L g1492 ( 
.A1(n_1458),
.A2(n_1430),
.B1(n_1427),
.B2(n_1443),
.C(n_1408),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1459),
.Y(n_1493)
);

AOI33xp33_ASAP7_75t_L g1494 ( 
.A1(n_1462),
.A2(n_1426),
.A3(n_1429),
.B1(n_1396),
.B2(n_1433),
.B3(n_1423),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1461),
.B(n_1407),
.Y(n_1495)
);

OA21x2_ASAP7_75t_L g1496 ( 
.A1(n_1444),
.A2(n_1417),
.B(n_1434),
.Y(n_1496)
);

AO21x1_ASAP7_75t_SL g1497 ( 
.A1(n_1458),
.A2(n_1435),
.B(n_1408),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1455),
.B(n_1414),
.Y(n_1498)
);

AND2x4_ASAP7_75t_SL g1499 ( 
.A(n_1462),
.B(n_1421),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1493),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1469),
.Y(n_1501)
);

NAND2x1_ASAP7_75t_L g1502 ( 
.A(n_1490),
.B(n_1454),
.Y(n_1502)
);

OAI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1471),
.A2(n_1465),
.B(n_1463),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1493),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1496),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1496),
.Y(n_1506)
);

BUFx4f_ASAP7_75t_L g1507 ( 
.A(n_1474),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1470),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1472),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1476),
.Y(n_1510)
);

INVx4_ASAP7_75t_SL g1511 ( 
.A(n_1473),
.Y(n_1511)
);

INVx2_ASAP7_75t_SL g1512 ( 
.A(n_1499),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1478),
.Y(n_1513)
);

AO21x2_ASAP7_75t_L g1514 ( 
.A1(n_1481),
.A2(n_1403),
.B(n_1398),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1494),
.B(n_1460),
.Y(n_1515)
);

INVx5_ASAP7_75t_L g1516 ( 
.A(n_1469),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1494),
.B(n_1454),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1482),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1497),
.B(n_1487),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1489),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1519),
.B(n_1497),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1515),
.B(n_1464),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1506),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1515),
.B(n_1486),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1519),
.B(n_1516),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1519),
.B(n_1473),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1502),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1502),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1506),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1519),
.B(n_1473),
.Y(n_1530)
);

INVx1_ASAP7_75t_SL g1531 ( 
.A(n_1501),
.Y(n_1531)
);

AND2x2_ASAP7_75t_SL g1532 ( 
.A(n_1507),
.B(n_1520),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1515),
.B(n_1464),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1504),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1506),
.Y(n_1535)
);

AOI211xp5_ASAP7_75t_L g1536 ( 
.A1(n_1503),
.A2(n_1484),
.B(n_1468),
.C(n_1485),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1507),
.A2(n_1479),
.B1(n_1454),
.B2(n_1480),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1517),
.B(n_1464),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1516),
.B(n_1491),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1506),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1510),
.B(n_1475),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1506),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1517),
.B(n_1510),
.Y(n_1543)
);

NAND3xp33_ASAP7_75t_L g1544 ( 
.A(n_1503),
.B(n_1492),
.C(n_1489),
.Y(n_1544)
);

INVxp67_ASAP7_75t_SL g1545 ( 
.A(n_1513),
.Y(n_1545)
);

AOI21xp33_ASAP7_75t_L g1546 ( 
.A1(n_1507),
.A2(n_1461),
.B(n_1477),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1508),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1508),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1513),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1505),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1501),
.Y(n_1551)
);

INVx3_ASAP7_75t_SL g1552 ( 
.A(n_1516),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1509),
.B(n_1483),
.Y(n_1553)
);

CKINVDCx16_ASAP7_75t_R g1554 ( 
.A(n_1503),
.Y(n_1554)
);

NAND2xp33_ASAP7_75t_L g1555 ( 
.A(n_1507),
.B(n_1488),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1524),
.B(n_1507),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1536),
.B(n_1507),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1536),
.B(n_1498),
.Y(n_1558)
);

NOR4xp25_ASAP7_75t_L g1559 ( 
.A(n_1544),
.B(n_1518),
.C(n_1512),
.D(n_1500),
.Y(n_1559)
);

AOI21xp33_ASAP7_75t_L g1560 ( 
.A1(n_1544),
.A2(n_1514),
.B(n_1520),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1549),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1521),
.B(n_1511),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1524),
.B(n_1495),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_1551),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1554),
.B(n_1498),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1521),
.B(n_1511),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1549),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1554),
.B(n_1487),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1555),
.A2(n_1454),
.B1(n_1512),
.B2(n_1456),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1526),
.B(n_1511),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1547),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1521),
.B(n_1526),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1547),
.Y(n_1573)
);

NAND2x1p5_ASAP7_75t_L g1574 ( 
.A(n_1532),
.B(n_1516),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1526),
.B(n_1511),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1530),
.B(n_1511),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1530),
.B(n_1511),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1532),
.B(n_1501),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1545),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1551),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1548),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1537),
.A2(n_1512),
.B1(n_1516),
.B2(n_1454),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1525),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1530),
.B(n_1511),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1532),
.A2(n_1454),
.B1(n_1512),
.B2(n_1456),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1525),
.B(n_1511),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1525),
.B(n_1501),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1548),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1572),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1579),
.B(n_1545),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1564),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1572),
.B(n_1552),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1562),
.B(n_1552),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1567),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1557),
.A2(n_1546),
.B1(n_1514),
.B2(n_1539),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1556),
.B(n_1553),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1588),
.Y(n_1597)
);

AND3x1_ASAP7_75t_L g1598 ( 
.A(n_1559),
.B(n_1528),
.C(n_1527),
.Y(n_1598)
);

NAND2x1p5_ASAP7_75t_L g1599 ( 
.A(n_1564),
.B(n_1531),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1563),
.B(n_1553),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1558),
.B(n_1531),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1562),
.B(n_1552),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1561),
.B(n_1522),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1566),
.B(n_1539),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1574),
.B(n_1546),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1578),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1588),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1580),
.B(n_1566),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1569),
.A2(n_1543),
.B1(n_1538),
.B2(n_1516),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1565),
.B(n_1568),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1585),
.B(n_1541),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1571),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1580),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1611),
.A2(n_1560),
.B1(n_1582),
.B2(n_1584),
.Y(n_1614)
);

NOR2x1p5_ASAP7_75t_L g1615 ( 
.A(n_1601),
.B(n_1570),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1604),
.B(n_1587),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1590),
.B(n_1533),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1606),
.B(n_1574),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1604),
.B(n_1587),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1613),
.Y(n_1620)
);

NAND2x1_ASAP7_75t_SL g1621 ( 
.A(n_1608),
.B(n_1527),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1597),
.Y(n_1622)
);

INVxp67_ASAP7_75t_L g1623 ( 
.A(n_1608),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1591),
.B(n_1583),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1597),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1598),
.A2(n_1570),
.B1(n_1584),
.B2(n_1576),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1599),
.Y(n_1627)
);

OAI31xp33_ASAP7_75t_SL g1628 ( 
.A1(n_1605),
.A2(n_1570),
.A3(n_1586),
.B(n_1577),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1594),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1599),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1607),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1608),
.B(n_1575),
.Y(n_1632)
);

INVx2_ASAP7_75t_SL g1633 ( 
.A(n_1621),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1623),
.B(n_1600),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1620),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1620),
.B(n_1591),
.Y(n_1636)
);

NOR2x1_ASAP7_75t_L g1637 ( 
.A(n_1627),
.B(n_1594),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1616),
.B(n_1589),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1621),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1616),
.B(n_1589),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1632),
.B(n_1593),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1632),
.Y(n_1642)
);

OAI221xp5_ASAP7_75t_SL g1643 ( 
.A1(n_1639),
.A2(n_1614),
.B1(n_1628),
.B2(n_1626),
.C(n_1595),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1633),
.B(n_1574),
.Y(n_1644)
);

OAI311xp33_ASAP7_75t_L g1645 ( 
.A1(n_1638),
.A2(n_1624),
.A3(n_1617),
.B1(n_1590),
.C1(n_1596),
.Y(n_1645)
);

OAI211xp5_ASAP7_75t_SL g1646 ( 
.A1(n_1636),
.A2(n_1629),
.B(n_1618),
.C(n_1630),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1634),
.B(n_1629),
.Y(n_1647)
);

AOI221xp5_ASAP7_75t_L g1648 ( 
.A1(n_1635),
.A2(n_1630),
.B1(n_1627),
.B2(n_1610),
.C(n_1609),
.Y(n_1648)
);

AOI211xp5_ASAP7_75t_SL g1649 ( 
.A1(n_1640),
.A2(n_1617),
.B(n_1625),
.C(n_1622),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1637),
.A2(n_1599),
.B(n_1619),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1639),
.Y(n_1651)
);

OAI21xp33_ASAP7_75t_L g1652 ( 
.A1(n_1643),
.A2(n_1641),
.B(n_1619),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1646),
.A2(n_1642),
.B1(n_1615),
.B2(n_1592),
.Y(n_1653)
);

OAI211xp5_ASAP7_75t_L g1654 ( 
.A1(n_1650),
.A2(n_1631),
.B(n_1612),
.C(n_1593),
.Y(n_1654)
);

AOI21xp33_ASAP7_75t_SL g1655 ( 
.A1(n_1647),
.A2(n_1603),
.B(n_1543),
.Y(n_1655)
);

AOI221xp5_ASAP7_75t_SL g1656 ( 
.A1(n_1648),
.A2(n_1602),
.B1(n_1592),
.B2(n_1607),
.C(n_1603),
.Y(n_1656)
);

NOR3x1_ASAP7_75t_L g1657 ( 
.A(n_1654),
.B(n_1644),
.C(n_1645),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1653),
.B(n_1651),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1656),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1652),
.B(n_1649),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1655),
.Y(n_1661)
);

NAND3xp33_ASAP7_75t_L g1662 ( 
.A(n_1652),
.B(n_1602),
.C(n_1583),
.Y(n_1662)
);

NOR4xp25_ASAP7_75t_L g1663 ( 
.A(n_1660),
.B(n_1581),
.C(n_1573),
.D(n_1550),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1661),
.Y(n_1664)
);

CKINVDCx20_ASAP7_75t_R g1665 ( 
.A(n_1659),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1662),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1659),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1666),
.B(n_1658),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1664),
.Y(n_1669)
);

NAND3xp33_ASAP7_75t_L g1670 ( 
.A(n_1667),
.B(n_1657),
.C(n_1586),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1668),
.B(n_1665),
.Y(n_1671)
);

OAI211xp5_ASAP7_75t_L g1672 ( 
.A1(n_1671),
.A2(n_1667),
.B(n_1670),
.C(n_1669),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1672),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1672),
.Y(n_1674)
);

INVx2_ASAP7_75t_SL g1675 ( 
.A(n_1674),
.Y(n_1675)
);

INVx1_ASAP7_75t_SL g1676 ( 
.A(n_1673),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_SL g1677 ( 
.A1(n_1676),
.A2(n_1663),
.B1(n_1527),
.B2(n_1528),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_SL g1678 ( 
.A1(n_1675),
.A2(n_1528),
.B1(n_1527),
.B2(n_1534),
.Y(n_1678)
);

XNOR2xp5_ASAP7_75t_L g1679 ( 
.A(n_1677),
.B(n_1678),
.Y(n_1679)
);

AO221x1_ASAP7_75t_L g1680 ( 
.A1(n_1679),
.A2(n_1528),
.B1(n_1540),
.B2(n_1535),
.C(n_1542),
.Y(n_1680)
);

NAND2x1_ASAP7_75t_L g1681 ( 
.A(n_1680),
.B(n_1575),
.Y(n_1681)
);

AOI22x1_ASAP7_75t_L g1682 ( 
.A1(n_1681),
.A2(n_1523),
.B1(n_1542),
.B2(n_1540),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1682),
.A2(n_1576),
.B1(n_1577),
.B2(n_1529),
.Y(n_1683)
);

AOI211xp5_ASAP7_75t_L g1684 ( 
.A1(n_1683),
.A2(n_1535),
.B(n_1523),
.C(n_1529),
.Y(n_1684)
);


endmodule