module fake_jpeg_2904_n_414 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_414);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_414;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_292;
wire n_213;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_44),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_13),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_45),
.B(n_53),
.Y(n_111)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_46),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_49),
.Y(n_127)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_75),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_51),
.Y(n_144)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_25),
.B(n_33),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_58),
.B(n_65),
.Y(n_128)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_59),
.Y(n_149)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_40),
.B(n_1),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g159 ( 
.A(n_66),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_14),
.Y(n_67)
);

NOR3xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_80),
.C(n_91),
.Y(n_103)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_68),
.Y(n_160)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_73),
.Y(n_134)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_38),
.B(n_14),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_76),
.Y(n_158)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_77),
.Y(n_136)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_79),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_82),
.Y(n_107)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_84),
.Y(n_108)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_37),
.B(n_1),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_88),
.Y(n_110)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_37),
.B(n_1),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_90),
.Y(n_129)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_93),
.Y(n_133)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_95),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_17),
.B(n_2),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_98),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_30),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_10),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_100),
.B(n_125),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_22),
.B1(n_27),
.B2(n_18),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_106),
.A2(n_149),
.B1(n_118),
.B2(n_105),
.Y(n_193)
);

OR2x4_ASAP7_75t_L g112 ( 
.A(n_53),
.B(n_27),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_112),
.A2(n_107),
.B(n_156),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_24),
.B1(n_22),
.B2(n_21),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_114),
.A2(n_118),
.B1(n_127),
.B2(n_115),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_45),
.A2(n_31),
.B(n_26),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_117),
.A2(n_136),
.B(n_135),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_74),
.A2(n_31),
.B1(n_24),
.B2(n_21),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_120),
.A2(n_138),
.B1(n_145),
.B2(n_148),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_75),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_141),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_54),
.B(n_18),
.C(n_17),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_47),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_131),
.A2(n_132),
.B1(n_147),
.B2(n_79),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_49),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_68),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_58),
.B(n_11),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_96),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_57),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_66),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_62),
.B(n_8),
.C(n_9),
.Y(n_151)
);

NAND2x1_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_156),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_71),
.B(n_10),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_155),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_48),
.B(n_10),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_63),
.B(n_11),
.C(n_76),
.Y(n_156)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_109),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_165),
.B(n_172),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_110),
.A2(n_112),
.B1(n_111),
.B2(n_140),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_174),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_167),
.A2(n_178),
.B1(n_190),
.B2(n_191),
.Y(n_211)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_100),
.A2(n_91),
.B1(n_97),
.B2(n_82),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_171),
.A2(n_194),
.B1(n_115),
.B2(n_137),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_133),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_159),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_173),
.B(n_188),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_122),
.A2(n_114),
.B1(n_129),
.B2(n_131),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_132),
.A2(n_147),
.B1(n_125),
.B2(n_134),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_L g237 ( 
.A1(n_175),
.A2(n_207),
.B1(n_161),
.B2(n_185),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_141),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_189),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_117),
.A2(n_134),
.B1(n_157),
.B2(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_101),
.A2(n_103),
.B(n_151),
.C(n_108),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_184),
.A2(n_198),
.B(n_201),
.C(n_200),
.Y(n_227)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_186),
.Y(n_214)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_126),
.B(n_142),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_158),
.B1(n_130),
.B2(n_142),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_126),
.A2(n_124),
.B1(n_149),
.B2(n_105),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_193),
.B(n_199),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_113),
.Y(n_195)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_203),
.B(n_139),
.Y(n_220)
);

A2O1A1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_135),
.A2(n_136),
.B(n_119),
.C(n_102),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_150),
.B(n_119),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_102),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_200),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_150),
.A2(n_123),
.B(n_143),
.C(n_146),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_123),
.B(n_146),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_202),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_L g203 ( 
.A1(n_143),
.A2(n_127),
.B(n_104),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_104),
.B(n_139),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_204),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_104),
.Y(n_205)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_115),
.B(n_137),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_205),
.C(n_201),
.Y(n_232)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_222),
.A2(n_226),
.B1(n_227),
.B2(n_237),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_137),
.B(n_198),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_223),
.A2(n_227),
.B(n_232),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_167),
.A2(n_137),
.B1(n_174),
.B2(n_182),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_194),
.A2(n_171),
.B1(n_182),
.B2(n_184),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_230),
.A2(n_240),
.B1(n_190),
.B2(n_195),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_202),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_166),
.A2(n_182),
.B(n_172),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_233),
.A2(n_170),
.B(n_177),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_180),
.A2(n_189),
.B1(n_165),
.B2(n_192),
.Y(n_240)
);

AOI32xp33_ASAP7_75t_L g241 ( 
.A1(n_170),
.A2(n_176),
.A3(n_180),
.B1(n_177),
.B2(n_186),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_204),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_242),
.A2(n_262),
.B(n_265),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_177),
.C(n_179),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_248),
.C(n_216),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g244 ( 
.A(n_208),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_244),
.B(n_241),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_212),
.B(n_215),
.Y(n_269)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_223),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_250),
.Y(n_275)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_238),
.Y(n_249)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_220),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_183),
.Y(n_251)
);

INVxp33_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_163),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_256),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_187),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_195),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_259),
.Y(n_288)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_169),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_261),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_230),
.A2(n_168),
.B1(n_196),
.B2(n_181),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_214),
.B(n_209),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_228),
.Y(n_281)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_239),
.A2(n_162),
.B1(n_164),
.B2(n_207),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_226),
.A2(n_211),
.B1(n_221),
.B2(n_239),
.Y(n_267)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_269),
.B(n_283),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_251),
.Y(n_279)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_282),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_240),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_257),
.B(n_212),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_242),
.B(n_212),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_285),
.B(n_291),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_286),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_243),
.C(n_285),
.Y(n_294)
);

AND2x6_ASAP7_75t_L g289 ( 
.A(n_245),
.B(n_211),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g309 ( 
.A1(n_289),
.A2(n_259),
.B(n_248),
.C(n_222),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_229),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_290),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_256),
.B(n_238),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_294),
.B(n_296),
.C(n_311),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_267),
.B1(n_260),
.B2(n_266),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_295),
.A2(n_312),
.B1(n_289),
.B2(n_252),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_243),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_266),
.B1(n_262),
.B2(n_255),
.Y(n_298)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_275),
.A2(n_247),
.B(n_250),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_303),
.A2(n_274),
.B(n_288),
.Y(n_317)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_270),
.Y(n_304)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_304),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_275),
.A2(n_265),
.B(n_261),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_305),
.A2(n_277),
.B(n_228),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_306),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_282),
.A2(n_272),
.B1(n_280),
.B2(n_288),
.Y(n_307)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_307),
.Y(n_325)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_308),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_309),
.B(n_289),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_269),
.B(n_264),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_272),
.A2(n_276),
.B1(n_283),
.B2(n_280),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_273),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_273),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_274),
.B(n_253),
.C(n_246),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_278),
.C(n_271),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_317),
.A2(n_314),
.B(n_301),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_303),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_318),
.B(n_322),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_320),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_291),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_324),
.A2(n_299),
.B(n_292),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_297),
.B(n_278),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_326),
.B(n_213),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_329),
.B(n_331),
.C(n_300),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_330),
.A2(n_336),
.B1(n_316),
.B2(n_335),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_294),
.C(n_300),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_271),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_332),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_333),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_277),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_334),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_249),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_293),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_295),
.A2(n_301),
.B1(n_309),
.B2(n_305),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_340),
.C(n_323),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_354),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_311),
.C(n_299),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_342),
.A2(n_352),
.B1(n_323),
.B2(n_326),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_292),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_349),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_327),
.B(n_302),
.Y(n_345)
);

MAJx2_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_351),
.C(n_353),
.Y(n_367)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_346),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_329),
.Y(n_349)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_350),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_327),
.B(n_229),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_219),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_219),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_348),
.A2(n_325),
.B1(n_316),
.B2(n_318),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_319),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_357),
.B(n_358),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_317),
.C(n_333),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_337),
.Y(n_360)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

FAx1_ASAP7_75t_L g362 ( 
.A(n_342),
.B(n_324),
.CI(n_317),
.CON(n_362),
.SN(n_362)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_362),
.B(n_341),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_322),
.Y(n_363)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_363),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_340),
.B(n_330),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_368),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_345),
.B(n_336),
.C(n_334),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_365),
.B(n_344),
.C(n_353),
.Y(n_370)
);

AOI221xp5_ASAP7_75t_L g369 ( 
.A1(n_355),
.A2(n_343),
.B1(n_341),
.B2(n_332),
.C(n_320),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_369),
.A2(n_362),
.B1(n_328),
.B2(n_315),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_379),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_372),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_354),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_373),
.B(n_377),
.Y(n_383)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_356),
.Y(n_376)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_376),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_361),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_378),
.B(n_319),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_366),
.B(n_338),
.C(n_351),
.Y(n_379)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_381),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_378),
.A2(n_362),
.B1(n_358),
.B2(n_365),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_384),
.B(n_386),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_367),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_387),
.B(n_389),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_366),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_375),
.B(n_357),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_390),
.B(n_370),
.Y(n_393)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_393),
.A2(n_394),
.B(n_388),
.Y(n_400)
);

O2A1O1Ixp33_ASAP7_75t_SL g394 ( 
.A1(n_385),
.A2(n_372),
.B(n_380),
.C(n_364),
.Y(n_394)
);

MAJx2_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_379),
.C(n_374),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_396),
.B(n_397),
.Y(n_399)
);

AOI322xp5_ASAP7_75t_L g397 ( 
.A1(n_381),
.A2(n_372),
.A3(n_315),
.B1(n_321),
.B2(n_367),
.C1(n_258),
.C2(n_231),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_321),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_398),
.B(n_395),
.Y(n_403)
);

AO21x1_ASAP7_75t_L g407 ( 
.A1(n_400),
.A2(n_403),
.B(n_404),
.Y(n_407)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_392),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_401),
.B(n_402),
.Y(n_405)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_391),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_391),
.A2(n_382),
.B(n_387),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_399),
.B(n_382),
.C(n_235),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_406),
.A2(n_408),
.B(n_225),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_404),
.B(n_258),
.Y(n_408)
);

BUFx5_ASAP7_75t_L g409 ( 
.A(n_407),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_409),
.A2(n_410),
.B(n_405),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_411),
.A2(n_412),
.B(n_218),
.Y(n_413)
);

AOI322xp5_ASAP7_75t_L g412 ( 
.A1(n_409),
.A2(n_231),
.A3(n_213),
.B1(n_216),
.B2(n_210),
.C1(n_235),
.C2(n_218),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_413),
.B(n_225),
.Y(n_414)
);


endmodule