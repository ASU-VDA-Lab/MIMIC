module real_jpeg_14642_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g91 ( 
.A(n_3),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_4),
.A2(n_35),
.B(n_36),
.C(n_42),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_4),
.B(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_4),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_4),
.A2(n_38),
.B1(n_68),
.B2(n_70),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_4),
.A2(n_50),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_4),
.B(n_83),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_5),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_62),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_5),
.A2(n_62),
.B1(n_68),
.B2(n_70),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_62),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_10),
.A2(n_68),
.B1(n_70),
.B2(n_74),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_74),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_12),
.A2(n_54),
.B1(n_68),
.B2(n_70),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_13),
.A2(n_68),
.B1(n_70),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_13),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_94),
.Y(n_113)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_15),
.A2(n_39),
.B1(n_40),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_15),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_15),
.A2(n_68),
.B1(n_70),
.B2(n_85),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_85),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_117),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_115),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_97),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_19),
.B(n_97),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_75),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_48),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_34),
.B1(n_46),
.B2(n_47),
.Y(n_21)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_23),
.B(n_52),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_23),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_23),
.A2(n_28),
.B1(n_139),
.B2(n_141),
.Y(n_138)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_23),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_24),
.A2(n_25),
.B1(n_89),
.B2(n_90),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_24),
.B(n_38),
.C(n_90),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_24),
.B(n_146),
.Y(n_145)
);

CKINVDCx6p67_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_28),
.B(n_113),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_50),
.B(n_51),
.Y(n_49)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_35),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B(n_39),
.Y(n_36)
);

HAxp5_ASAP7_75t_SL g110 ( 
.A(n_38),
.B(n_40),
.CON(n_110),
.SN(n_110)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_38),
.B(n_50),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_38),
.B(n_92),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_39),
.A2(n_40),
.B1(n_66),
.B2(n_67),
.Y(n_71)
);

NOR3xp33_ASAP7_75t_L g111 ( 
.A(n_39),
.B(n_67),
.C(n_68),
.Y(n_111)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.C(n_59),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_49),
.A2(n_55),
.B1(n_56),
.B2(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_50),
.B(n_53),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_50),
.A2(n_140),
.B1(n_148),
.B2(n_149),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_76)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_59),
.B(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_65),
.B2(n_72),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_61),
.A2(n_64),
.B1(n_83),
.B2(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_73),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_71),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

OA22x2_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_SL g108 ( 
.A1(n_66),
.A2(n_70),
.B(n_109),
.C(n_111),
.Y(n_108)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_68),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_70),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_70),
.B(n_132),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_81),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_93),
.B(n_95),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_87),
.A2(n_104),
.B1(n_106),
.B2(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_87),
.A2(n_106),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_87),
.A2(n_106),
.B1(n_125),
.B2(n_135),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.C(n_107),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_107),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B(n_105),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_112),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_126),
.B(n_171),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_121),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.C(n_124),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_124),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_166),
.B(n_170),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_155),
.B(n_165),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_143),
.B(n_154),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_138),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_138),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_136),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_149),
.B(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_150),
.B(n_153),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_152),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_157),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_161),
.C(n_164),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_169),
.Y(n_170)
);


endmodule