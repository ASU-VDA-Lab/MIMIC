module fake_jpeg_1996_n_262 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_107;
wire n_39;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx10_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_41),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_57),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_28),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_58),
.Y(n_86)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_28),
.B(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_60),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_15),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_61),
.Y(n_105)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_20),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_74),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_73),
.Y(n_92)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_36),
.B(n_0),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_15),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_44),
.A2(n_18),
.B1(n_36),
.B2(n_35),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_79),
.A2(n_95),
.B1(n_114),
.B2(n_9),
.Y(n_148)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_25),
.B1(n_35),
.B2(n_34),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_89),
.A2(n_117),
.B1(n_9),
.B2(n_11),
.Y(n_151)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_40),
.A2(n_24),
.B1(n_34),
.B2(n_30),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_104),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_46),
.B(n_20),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_41),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_24),
.B1(n_30),
.B2(n_25),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_21),
.B1(n_9),
.B2(n_11),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_51),
.B(n_3),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_115),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_42),
.A2(n_39),
.B1(n_29),
.B2(n_23),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_L g115 ( 
.A(n_60),
.B(n_15),
.C(n_29),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_42),
.A2(n_39),
.B1(n_23),
.B2(n_22),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_59),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_3),
.B(n_4),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_130),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_65),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_138),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_91),
.B(n_3),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_125),
.B(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_50),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_127),
.B(n_139),
.Y(n_168)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_55),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_77),
.A2(n_63),
.B1(n_41),
.B2(n_21),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_141),
.B1(n_83),
.B2(n_137),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_55),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_6),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_78),
.B(n_21),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_137),
.A2(n_87),
.B(n_106),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_6),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_7),
.Y(n_139)
);

OA21x2_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_104),
.B(n_79),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_78),
.B(n_7),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_149),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_89),
.A2(n_95),
.B(n_114),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_147),
.Y(n_174)
);

HAxp5_ASAP7_75t_SL g145 ( 
.A(n_81),
.B(n_12),
.CON(n_145),
.SN(n_145)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_145),
.Y(n_171)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_148),
.A2(n_150),
.B1(n_151),
.B2(n_88),
.Y(n_170)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_140),
.A2(n_117),
.B1(n_113),
.B2(n_99),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_152),
.A2(n_165),
.B1(n_170),
.B2(n_175),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_103),
.B(n_106),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_153),
.A2(n_177),
.B(n_147),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_119),
.A2(n_113),
.B1(n_99),
.B2(n_98),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_159),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_121),
.A2(n_98),
.B1(n_84),
.B2(n_82),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_SL g162 ( 
.A(n_138),
.B(n_12),
.C(n_94),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_118),
.C(n_141),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_129),
.A2(n_103),
.B1(n_84),
.B2(n_116),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_88),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_173),
.B(n_176),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_83),
.B1(n_129),
.B2(n_135),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_140),
.A2(n_129),
.B(n_124),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_168),
.B(n_125),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_185),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_163),
.B(n_132),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_158),
.Y(n_204)
);

NAND3xp33_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_132),
.C(n_142),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_153),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_187),
.B(n_189),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_150),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_192),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_120),
.C(n_131),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_199),
.C(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_SL g207 ( 
.A1(n_193),
.A2(n_197),
.B(n_198),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_146),
.B1(n_160),
.B2(n_167),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_128),
.Y(n_197)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_149),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_202),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_193),
.A2(n_157),
.B(n_173),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_211),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_156),
.B(n_174),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_215),
.B(n_166),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_172),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_195),
.A2(n_156),
.B1(n_174),
.B2(n_175),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_213),
.A2(n_214),
.B1(n_186),
.B2(n_179),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_152),
.B1(n_158),
.B2(n_177),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_166),
.C(n_159),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_220),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_204),
.B(n_191),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_180),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_201),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_223),
.B(n_224),
.Y(n_235)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_212),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_225),
.A2(n_226),
.B1(n_228),
.B2(n_215),
.Y(n_229)
);

OAI22x1_ASAP7_75t_L g226 ( 
.A1(n_214),
.A2(n_198),
.B1(n_196),
.B2(n_179),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_183),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_227),
.A2(n_200),
.B(n_203),
.C(n_211),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_213),
.A2(n_182),
.B1(n_192),
.B2(n_181),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_237),
.B1(n_216),
.B2(n_206),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_231),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_222),
.B(n_171),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_227),
.C(n_223),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_220),
.B(n_219),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_236),
.Y(n_238)
);

A2O1A1O1Ixp25_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_201),
.B(n_162),
.C(n_171),
.D(n_154),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_226),
.B1(n_217),
.B2(n_228),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_239),
.A2(n_235),
.B1(n_216),
.B2(n_237),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_143),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_224),
.C(n_221),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_232),
.C(n_206),
.Y(n_246)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_244),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_245),
.B(n_246),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_249),
.C(n_245),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_190),
.B(n_123),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_241),
.C(n_239),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_188),
.C(n_194),
.Y(n_256)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_246),
.B(n_240),
.CI(n_241),
.CON(n_251),
.SN(n_251)
);

NOR2x1_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_248),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_238),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_254),
.A2(n_253),
.B(n_250),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_255),
.B(n_256),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_255),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_259),
.B(n_260),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_257),
.A2(n_251),
.B1(n_123),
.B2(n_143),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_143),
.Y(n_262)
);


endmodule