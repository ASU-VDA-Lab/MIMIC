module real_jpeg_6722_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_487;
wire n_242;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g168 ( 
.A(n_0),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_0),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_0),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_0),
.Y(n_283)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_0),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_0),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_1),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_1),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_1),
.A2(n_54),
.B1(n_204),
.B2(n_274),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_1),
.A2(n_204),
.B1(n_285),
.B2(n_390),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g450 ( 
.A1(n_1),
.A2(n_204),
.B1(n_451),
.B2(n_453),
.Y(n_450)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_2),
.Y(n_190)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_2),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_2),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_3),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_3),
.A2(n_49),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_3),
.A2(n_49),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_3),
.A2(n_49),
.B1(n_285),
.B2(n_287),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_4),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_5),
.A2(n_42),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_5),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_5),
.A2(n_189),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g401 ( 
.A1(n_5),
.A2(n_189),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_5),
.A2(n_189),
.B1(n_424),
.B2(n_427),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_8),
.Y(n_118)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_8),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_8),
.Y(n_384)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_9),
.Y(n_94)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_10),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_10),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_10),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_11),
.A2(n_217),
.B1(n_219),
.B2(n_222),
.Y(n_216)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_11),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_11),
.A2(n_222),
.B1(n_260),
.B2(n_271),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_11),
.A2(n_181),
.B1(n_222),
.B2(n_305),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_L g364 ( 
.A1(n_11),
.A2(n_222),
.B1(n_365),
.B2(n_366),
.Y(n_364)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_12),
.Y(n_83)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_13),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_13),
.A2(n_162),
.B1(n_219),
.B2(n_378),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_13),
.B(n_384),
.C(n_385),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_13),
.B(n_90),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_13),
.B(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_13),
.B(n_132),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_13),
.B(n_212),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_14),
.A2(n_58),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_14),
.A2(n_75),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_14),
.A2(n_75),
.B1(n_218),
.B2(n_226),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_14),
.A2(n_75),
.B1(n_348),
.B2(n_349),
.Y(n_347)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_16),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_16),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_16),
.A2(n_72),
.B1(n_169),
.B2(n_174),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_16),
.A2(n_72),
.B1(n_225),
.B2(n_230),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_16),
.A2(n_72),
.B1(n_209),
.B2(n_322),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_17),
.A2(n_53),
.B1(n_57),
.B2(n_60),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_17),
.A2(n_60),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_17),
.A2(n_60),
.B1(n_169),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_17),
.A2(n_60),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_18),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_18),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_18),
.A2(n_193),
.B1(n_209),
.B2(n_211),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_18),
.A2(n_193),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_18),
.A2(n_193),
.B1(n_306),
.B2(n_397),
.Y(n_396)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_62),
.B(n_528),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_50),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_26),
.B(n_50),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_37),
.B(n_44),
.Y(n_26)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_27),
.B(n_192),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_27),
.B(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_28),
.A2(n_51),
.B1(n_188),
.B2(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_28),
.B(n_162),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_33),
.Y(n_152)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_33),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_35),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_35),
.Y(n_206)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_35),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_35),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_37),
.B(n_192),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_37),
.A2(n_250),
.B(n_254),
.Y(n_249)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_41),
.Y(n_156)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_42),
.Y(n_194)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_43),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_43),
.B(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_51),
.B1(n_52),
.B2(n_61),
.Y(n_50)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_50),
.B(n_64),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_61),
.B1(n_68),
.B2(n_73),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_51),
.A2(n_52),
.B1(n_61),
.B2(n_73),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_51),
.A2(n_255),
.B(n_273),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_51),
.A2(n_61),
.B1(n_68),
.B2(n_500),
.Y(n_499)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_56),
.Y(n_253)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_61),
.A2(n_188),
.B(n_191),
.Y(n_187)
);

AO21x1_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_141),
.B(n_527),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_137),
.C(n_138),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_65),
.A2(n_66),
.B1(n_523),
.B2(n_524),
.Y(n_522)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_76),
.C(n_108),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_67),
.B(n_515),
.Y(n_514)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_76),
.A2(n_108),
.B1(n_109),
.B2(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_76),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_99),
.B1(n_104),
.B2(n_105),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g139 ( 
.A(n_77),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_77),
.A2(n_104),
.B1(n_201),
.B2(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_77),
.A2(n_104),
.B1(n_270),
.B2(n_321),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_77),
.A2(n_99),
.B1(n_104),
.B2(n_504),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_90),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_82),
.Y(n_464)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_84),
.Y(n_212)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_85),
.Y(n_352)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_88),
.Y(n_348)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_89),
.Y(n_203)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_89),
.Y(n_259)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_90),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

AOI22x1_ASAP7_75t_L g267 ( 
.A1(n_90),
.A2(n_139),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_90),
.A2(n_139),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

AO22x2_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_93),
.B1(n_95),
.B2(n_97),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_93),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_94),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_94),
.Y(n_246)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_94),
.Y(n_404)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_94),
.Y(n_467)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_113),
.B1(n_116),
.B2(n_119),
.Y(n_112)
);

INVx11_ASAP7_75t_L g402 ( 
.A(n_95),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_96),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_96),
.Y(n_233)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_97),
.Y(n_468)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_100),
.Y(n_260)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_104),
.B(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_104),
.A2(n_257),
.B(n_302),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_108),
.A2(n_109),
.B1(n_502),
.B2(n_503),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_108),
.B(n_499),
.C(n_502),
.Y(n_510)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_131),
.B(n_133),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_110),
.A2(n_131),
.B1(n_216),
.B2(n_223),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_110),
.A2(n_377),
.B(n_379),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_110),
.A2(n_131),
.B1(n_401),
.B2(n_450),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_110),
.A2(n_379),
.B(n_450),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_111),
.B(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_111),
.A2(n_132),
.B1(n_224),
.B2(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_111),
.A2(n_132),
.B1(n_279),
.B2(n_329),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_111),
.A2(n_132),
.B1(n_329),
.B2(n_355),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_122),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_122),
.A2(n_243),
.B(n_401),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_128),
.B2(n_130),
.Y(n_122)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_126),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_127),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_129),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g428 ( 
.A(n_129),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_131),
.A2(n_216),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_132),
.B(n_244),
.Y(n_379)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_133),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_135),
.Y(n_332)
);

INVx5_ASAP7_75t_L g452 ( 
.A(n_135),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_137),
.B(n_138),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_139),
.A2(n_200),
.B(n_207),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_139),
.B(n_268),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_139),
.A2(n_207),
.B(n_456),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_521),
.B(n_526),
.Y(n_141)
);

AOI21x1_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_493),
.B(n_518),
.Y(n_142)
);

OAI311xp33_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_314),
.A3(n_370),
.B1(n_487),
.C1(n_492),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_292),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_146),
.A2(n_489),
.B(n_490),
.Y(n_488)
);

NOR2x1_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_261),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_147),
.B(n_261),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_213),
.C(n_241),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_148),
.B(n_312),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_185),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_149),
.B(n_186),
.C(n_199),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_163),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_150),
.A2(n_163),
.B1(n_164),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_150),
.Y(n_299)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_153),
.A3(n_154),
.B1(n_157),
.B2(n_161),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_158),
.Y(n_157)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_SL g250 ( 
.A1(n_161),
.A2(n_162),
.B(n_251),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_162),
.A2(n_165),
.B(n_393),
.Y(n_420)
);

OAI21xp33_ASAP7_75t_SL g456 ( 
.A1(n_162),
.A2(n_322),
.B(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_172),
.B1(n_175),
.B2(n_178),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_165),
.A2(n_236),
.B1(n_281),
.B2(n_284),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_165),
.A2(n_284),
.B(n_334),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_165),
.A2(n_389),
.B(n_393),
.Y(n_388)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_166),
.A2(n_179),
.B1(n_235),
.B2(n_239),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_166),
.A2(n_173),
.B1(n_304),
.B2(n_309),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_166),
.B(n_396),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_166),
.A2(n_437),
.B1(n_438),
.B2(n_439),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_168),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_168),
.Y(n_419)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_168),
.Y(n_431)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

BUFx8_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g289 ( 
.A(n_171),
.Y(n_289)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_171),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_171),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_184),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_198),
.B2(n_199),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_190),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_191),
.B(n_363),
.Y(n_362)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_208),
.Y(n_268)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_213),
.A2(n_214),
.B1(n_241),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_234),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_215),
.B(n_234),
.Y(n_265)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_229),
.Y(n_382)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_233),
.Y(n_378)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_237),
.Y(n_397)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_238),
.Y(n_386)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_241),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_248),
.C(n_256),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_242),
.B(n_256),
.Y(n_295)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AOI32xp33_ASAP7_75t_L g462 ( 
.A1(n_246),
.A2(n_260),
.A3(n_458),
.B1(n_463),
.B2(n_465),
.Y(n_462)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_247),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_248),
.A2(n_249),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_262),
.B(n_277),
.C(n_290),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_277),
.B1(n_290),
.B2(n_291),
.Y(n_263)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_265),
.B(n_267),
.C(n_276),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_272),
.B1(n_275),
.B2(n_276),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_267),
.Y(n_275)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_272),
.Y(n_276)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_278),
.B(n_280),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_311),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_293),
.B(n_311),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_297),
.C(n_300),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_294),
.B(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_297),
.A2(n_298),
.B1(n_300),
.B2(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_300),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.C(n_310),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_301),
.B(n_478),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_303),
.B(n_310),
.Y(n_478)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_304),
.Y(n_461)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_SL g306 ( 
.A(n_307),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp33_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_367),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_SL g487 ( 
.A1(n_315),
.A2(n_367),
.B(n_488),
.C(n_491),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_339),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_316),
.B(n_339),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_326),
.C(n_338),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g369 ( 
.A(n_317),
.B(n_326),
.CI(n_338),
.CON(n_369),
.SN(n_369)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_318),
.B(n_320),
.C(n_325),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_325),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_321),
.Y(n_346)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_333),
.B2(n_337),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_333),
.Y(n_359)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_333),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_333),
.A2(n_337),
.B1(n_361),
.B2(n_362),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_333),
.A2(n_359),
.B(n_362),
.Y(n_496)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_340),
.B(n_343),
.C(n_357),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_343),
.B1(n_357),
.B2(n_358),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_353),
.B(n_356),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_345),
.B(n_354),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_347),
.Y(n_504)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

FAx1_ASAP7_75t_SL g495 ( 
.A(n_356),
.B(n_496),
.CI(n_497),
.CON(n_495),
.SN(n_495)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_356),
.B(n_496),
.C(n_497),
.Y(n_517)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_364),
.Y(n_500)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_365),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_368),
.B(n_369),
.Y(n_491)
);

BUFx24_ASAP7_75t_SL g531 ( 
.A(n_369),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_481),
.B(n_486),
.Y(n_370)
);

AO21x1_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_470),
.B(n_480),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_373),
.A2(n_444),
.B(n_469),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_407),
.B(n_443),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_387),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_375),
.B(n_387),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_380),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_376),
.A2(n_380),
.B1(n_381),
.B2(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_376),
.Y(n_441)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_398),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_388),
.B(n_399),
.C(n_406),
.Y(n_445)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_389),
.Y(n_438)
);

INVx6_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_396),
.Y(n_393)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_399),
.A2(n_400),
.B1(n_405),
.B2(n_406),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_402),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_435),
.B(n_442),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_421),
.B(n_434),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_420),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_417),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_418),
.Y(n_439)
);

INVx8_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_422),
.B(n_433),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_433),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_429),
.B(n_432),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_423),
.Y(n_437)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_431),
.A2(n_432),
.B(n_461),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_440),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_436),
.B(n_440),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_445),
.B(n_446),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_459),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_449),
.B1(n_454),
.B2(n_455),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_454),
.C(n_459),
.Y(n_471)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVxp33_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_462),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_462),
.Y(n_476)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_468),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_472),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_471),
.B(n_472),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_473),
.A2(n_474),
.B1(n_477),
.B2(n_479),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_475),
.B(n_476),
.C(n_479),
.Y(n_482)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_477),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_483),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_482),
.B(n_483),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_507),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_495),
.B(n_506),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_495),
.B(n_506),
.Y(n_519)
);

BUFx24_ASAP7_75t_SL g530 ( 
.A(n_495),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_498),
.A2(n_499),
.B1(n_501),
.B2(n_505),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_498),
.A2(n_499),
.B1(n_513),
.B2(n_514),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_498),
.B(n_509),
.C(n_513),
.Y(n_525)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_501),
.Y(n_505)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_507),
.A2(n_519),
.B(n_520),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_508),
.B(n_517),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_517),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_509),
.A2(n_510),
.B1(n_511),
.B2(n_512),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_525),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_522),
.B(n_525),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_524),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_529),
.Y(n_528)
);


endmodule