module fake_jpeg_4613_n_321 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_16),
.B(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_25),
.Y(n_67)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx2_ASAP7_75t_SL g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_49),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_12),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_45),
.B(n_12),
.Y(n_76)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

AND2x4_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_32),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_50),
.A2(n_22),
.B(n_1),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_19),
.B1(n_20),
.B2(n_34),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_53),
.A2(n_69),
.B1(n_89),
.B2(n_95),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_19),
.B(n_32),
.C(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_54),
.B(n_55),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_26),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_19),
.B1(n_20),
.B2(n_34),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_56),
.A2(n_77),
.B(n_10),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_58),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_15),
.Y(n_59)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_32),
.B1(n_29),
.B2(n_23),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_60),
.B(n_66),
.C(n_3),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_15),
.Y(n_61)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_39),
.A2(n_31),
.B1(n_28),
.B2(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_70),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_28),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_68),
.B(n_78),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_17),
.B1(n_33),
.B2(n_16),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_31),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_79),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_35),
.B1(n_18),
.B2(n_14),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_73),
.A2(n_98),
.B1(n_0),
.B2(n_1),
.Y(n_117)
);

CKINVDCx6p67_ASAP7_75t_R g74 ( 
.A(n_41),
.Y(n_74)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_41),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_75),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_80),
.Y(n_109)
);

HAxp5_ASAP7_75t_SL g77 ( 
.A(n_41),
.B(n_25),
.CON(n_77),
.SN(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_27),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_82),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_25),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_27),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_83),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_22),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_0),
.Y(n_114)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_86),
.Y(n_116)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_91),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_40),
.A2(n_22),
.B1(n_35),
.B2(n_18),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_36),
.A2(n_27),
.B1(n_24),
.B2(n_18),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_90),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_37),
.B(n_24),
.Y(n_91)
);

CKINVDCx6p67_ASAP7_75t_R g92 ( 
.A(n_46),
.Y(n_92)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_94),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_22),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_36),
.A2(n_24),
.B1(n_35),
.B2(n_18),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_40),
.A2(n_22),
.B1(n_35),
.B2(n_11),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_101),
.A2(n_115),
.B(n_77),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_0),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_60),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_114),
.B(n_126),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_127),
.B1(n_128),
.B2(n_50),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_87),
.B(n_92),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_55),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_50),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_129),
.B(n_130),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_101),
.A2(n_94),
.B1(n_54),
.B2(n_63),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_131),
.A2(n_142),
.B(n_104),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_66),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_132),
.B(n_135),
.Y(n_200)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_133),
.B(n_134),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_127),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_51),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_136),
.A2(n_110),
.B(n_122),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_84),
.C(n_67),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_139),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_87),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_140),
.B(n_141),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_82),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_105),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_144),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_113),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_92),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_108),
.B(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_146),
.B(n_151),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

INVxp33_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_52),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_65),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_156),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_56),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_103),
.B(n_86),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_152),
.B(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_95),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_154),
.B(n_157),
.Y(n_190)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_92),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_105),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_70),
.Y(n_158)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_117),
.B1(n_112),
.B2(n_126),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_159),
.A2(n_164),
.B1(n_64),
.B2(n_97),
.Y(n_189)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_124),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_104),
.B(n_70),
.Y(n_162)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_93),
.B1(n_85),
.B2(n_72),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_159),
.A2(n_110),
.B1(n_128),
.B2(n_125),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_171),
.A2(n_188),
.B1(n_189),
.B2(n_193),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_111),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_173),
.A2(n_186),
.B(n_136),
.Y(n_214)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_114),
.Y(n_180)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_182),
.B(n_201),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_114),
.Y(n_184)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_124),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_185),
.B(n_194),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_141),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_130),
.A2(n_72),
.B1(n_97),
.B2(n_81),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_140),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_151),
.A2(n_64),
.B1(n_120),
.B2(n_106),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_106),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_134),
.A2(n_120),
.B1(n_58),
.B2(n_74),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_145),
.B1(n_100),
.B2(n_158),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_74),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_202),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_143),
.A2(n_120),
.B1(n_74),
.B2(n_107),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_199),
.B1(n_164),
.B2(n_129),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_143),
.A2(n_107),
.B1(n_57),
.B2(n_100),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_149),
.B(n_62),
.Y(n_201)
);

NOR3xp33_ASAP7_75t_L g202 ( 
.A(n_132),
.B(n_6),
.C(n_8),
.Y(n_202)
);

NAND2xp33_ASAP7_75t_SL g205 ( 
.A(n_178),
.B(n_142),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_205),
.B(n_223),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_215),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_183),
.A2(n_186),
.B1(n_192),
.B2(n_131),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_226),
.B1(n_188),
.B2(n_169),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_137),
.C(n_146),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_166),
.C(n_194),
.Y(n_233)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_214),
.A2(n_200),
.B(n_185),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_181),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_147),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_216),
.B(n_219),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_168),
.A2(n_160),
.B1(n_139),
.B2(n_133),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_227),
.B1(n_167),
.B2(n_175),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_191),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_218),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_190),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_197),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_220),
.B(n_221),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_173),
.Y(n_221)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_179),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_177),
.B(n_135),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_176),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_170),
.B(n_147),
.Y(n_229)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_229),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_189),
.A2(n_138),
.B1(n_154),
.B2(n_139),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_230),
.A2(n_168),
.B1(n_170),
.B2(n_182),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_232),
.A2(n_244),
.B1(n_249),
.B2(n_209),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_236),
.C(n_237),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_241),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_235),
.B(n_250),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_165),
.C(n_201),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_165),
.C(n_187),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_204),
.Y(n_238)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_221),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_184),
.C(n_180),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_251),
.C(n_207),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_169),
.B1(n_171),
.B2(n_196),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_248),
.A2(n_203),
.B(n_220),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_169),
.B1(n_200),
.B2(n_195),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_173),
.B1(n_198),
.B2(n_167),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_199),
.C(n_193),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_206),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_253),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_248),
.A2(n_203),
.B(n_213),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_254),
.A2(n_265),
.B(n_237),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_256),
.A2(n_259),
.B1(n_268),
.B2(n_208),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_258),
.A2(n_241),
.B(n_238),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_209),
.B1(n_232),
.B2(n_249),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_261),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_214),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_263),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_251),
.A2(n_218),
.B(n_207),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_219),
.B1(n_228),
.B2(n_227),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_240),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_234),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_205),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_284),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_258),
.A2(n_243),
.B(n_252),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_275),
.A2(n_285),
.B1(n_264),
.B2(n_262),
.Y(n_292)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_266),
.B(n_247),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_278),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_269),
.B(n_215),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_266),
.B(n_239),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_162),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_263),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_267),
.A2(n_236),
.B1(n_242),
.B2(n_233),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_174),
.B1(n_225),
.B2(n_163),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_271),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_255),
.C(n_260),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_290),
.C(n_293),
.Y(n_299)
);

O2A1O1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_262),
.B(n_254),
.C(n_270),
.Y(n_287)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_265),
.Y(n_290)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_255),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_294),
.B(n_283),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_264),
.C(n_263),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_297),
.B(n_272),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_280),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_283),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_302),
.B(n_305),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_303),
.Y(n_308)
);

OAI21xp33_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_276),
.B(n_285),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_274),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_281),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_310),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_304),
.B(n_291),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_210),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_287),
.B1(n_295),
.B2(n_174),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_302),
.B(n_281),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_300),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_316),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_314),
.A2(n_307),
.B(n_282),
.C(n_308),
.Y(n_317)
);

NAND3xp33_ASAP7_75t_SL g316 ( 
.A(n_312),
.B(n_288),
.C(n_290),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_315),
.C(n_299),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_318),
.C(n_299),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_303),
.Y(n_321)
);


endmodule