module fake_jpeg_6826_n_317 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_16),
.Y(n_35)
);

INVx5_ASAP7_75t_SL g95 ( 
.A(n_35),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_22),
.B(n_12),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_22),
.B(n_12),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_14),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_41),
.B(n_14),
.Y(n_64)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx5_ASAP7_75t_SL g123 ( 
.A(n_48),
.Y(n_123)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_50),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_23),
.B1(n_18),
.B2(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_51),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_106)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_57),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_18),
.B1(n_23),
.B2(n_34),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_56),
.A2(n_74),
.B1(n_77),
.B2(n_81),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_58),
.B(n_72),
.Y(n_100)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_64),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_25),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_61),
.A2(n_67),
.B(n_69),
.C(n_76),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_66),
.B(n_71),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_23),
.B1(n_24),
.B2(n_19),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_27),
.B(n_29),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_28),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g112 ( 
.A(n_73),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_40),
.A2(n_17),
.B1(n_26),
.B2(n_21),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_36),
.B(n_17),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_75),
.B(n_78),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_15),
.B1(n_21),
.B2(n_26),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_43),
.A2(n_15),
.B1(n_47),
.B2(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_20),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_20),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_79),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_44),
.B(n_27),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_80),
.B(n_85),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_33),
.B1(n_27),
.B2(n_29),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_20),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_44),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_37),
.B(n_33),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_90),
.Y(n_107)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_41),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_39),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_42),
.A2(n_29),
.B1(n_32),
.B2(n_31),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_37),
.B(n_1),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_2),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_110),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_32),
.B1(n_31),
.B2(n_4),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_120),
.B1(n_77),
.B2(n_76),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_61),
.A2(n_32),
.B(n_31),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_116),
.A2(n_97),
.B(n_96),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_48),
.A2(n_32),
.B1(n_31),
.B2(n_4),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_90),
.A2(n_32),
.B1(n_3),
.B2(n_4),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_133),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_138),
.B1(n_140),
.B2(n_143),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_101),
.A2(n_94),
.B1(n_95),
.B2(n_93),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

NOR2x1_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_67),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_132),
.A2(n_8),
.B(n_9),
.Y(n_199)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_117),
.B(n_49),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_145),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_80),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_136),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_107),
.B(n_56),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_85),
.B1(n_68),
.B2(n_73),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_114),
.B1(n_119),
.B2(n_121),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_127),
.A2(n_88),
.B1(n_87),
.B2(n_53),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_64),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_139),
.B(n_141),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_127),
.A2(n_84),
.B1(n_83),
.B2(n_71),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_49),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_63),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_142),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_127),
.A2(n_52),
.B1(n_66),
.B2(n_68),
.Y(n_143)
);

AO21x1_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_60),
.B(n_58),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_144),
.A2(n_160),
.B(n_8),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_148),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_117),
.B(n_52),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_50),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_50),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_152),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_99),
.B(n_2),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_63),
.Y(n_153)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_118),
.A2(n_59),
.B1(n_106),
.B2(n_121),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_54),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_115),
.B(n_2),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_3),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_113),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_100),
.C(n_111),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_136),
.C(n_143),
.Y(n_166)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_3),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_5),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_186),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_149),
.C(n_147),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_145),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_169),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_171),
.A2(n_11),
.B(n_175),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_156),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_173),
.B(n_174),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_109),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_182),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_162),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_178),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_132),
.A2(n_103),
.B1(n_119),
.B2(n_122),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_100),
.B1(n_120),
.B2(n_108),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_185),
.B1(n_187),
.B2(n_192),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_110),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_137),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_183),
.B(n_191),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_138),
.A2(n_108),
.B1(n_103),
.B2(n_55),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_132),
.A2(n_105),
.B1(n_102),
.B2(n_7),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_159),
.A2(n_55),
.B1(n_97),
.B2(n_96),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_137),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_160),
.A2(n_62),
.B1(n_105),
.B2(n_102),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_133),
.B(n_3),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_152),
.Y(n_205)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_194),
.Y(n_200)
);

A2O1A1O1Ixp25_ASAP7_75t_L g196 ( 
.A1(n_158),
.A2(n_105),
.B(n_102),
.C(n_62),
.D(n_10),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_199),
.C(n_137),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_130),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_197),
.A2(n_198),
.B1(n_128),
.B2(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_227),
.C(n_198),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_212),
.Y(n_247)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_134),
.A3(n_144),
.B1(n_139),
.B2(n_141),
.C1(n_153),
.C2(n_137),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_176),
.A3(n_196),
.B1(n_181),
.B2(n_189),
.C1(n_184),
.C2(n_173),
.Y(n_237)
);

NAND3xp33_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_196),
.C(n_177),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_216),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_151),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_128),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_214),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_148),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_R g217 ( 
.A(n_199),
.B(n_144),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_190),
.B(n_181),
.Y(n_231)
);

OAI32xp33_ASAP7_75t_L g219 ( 
.A1(n_164),
.A2(n_146),
.A3(n_157),
.B1(n_155),
.B2(n_161),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_219),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_164),
.A2(n_150),
.B1(n_10),
.B2(n_11),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_183),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_191),
.A2(n_10),
.B1(n_11),
.B2(n_180),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_225),
.Y(n_244)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_165),
.B(n_170),
.C(n_187),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_234),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_218),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_230),
.B(n_184),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_231),
.A2(n_245),
.B(n_205),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_176),
.C(n_172),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_215),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_236),
.Y(n_260)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_237),
.Y(n_267)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_239),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_220),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_212),
.B(n_172),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_241),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_203),
.B(n_182),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_174),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_243),
.Y(n_253)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_185),
.C(n_189),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_201),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_213),
.B(n_193),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_201),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_224),
.B(n_215),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_251),
.A2(n_265),
.B(n_266),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_206),
.B1(n_222),
.B2(n_208),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_254),
.A2(n_255),
.B1(n_262),
.B2(n_186),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_206),
.B1(n_211),
.B2(n_171),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_256),
.B(n_259),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_234),
.C(n_240),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_248),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_233),
.A2(n_179),
.B1(n_210),
.B2(n_167),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_247),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_236),
.A2(n_221),
.B(n_219),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_247),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_249),
.B(n_242),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_281),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_274),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_243),
.B1(n_238),
.B2(n_231),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_272),
.A2(n_261),
.B1(n_254),
.B2(n_262),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_229),
.B(n_242),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_273),
.A2(n_269),
.B(n_279),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_263),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_255),
.A2(n_249),
.B1(n_246),
.B2(n_228),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_275),
.B(n_277),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_278),
.C(n_264),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_241),
.C(n_250),
.Y(n_278)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_251),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_280),
.A2(n_229),
.B1(n_232),
.B2(n_216),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_271),
.B1(n_270),
.B2(n_280),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_289),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_258),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_290),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_293),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_226),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_258),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_292),
.C(n_275),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_266),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_302),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_295),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_223),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_299),
.C(n_301),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_273),
.B1(n_272),
.B2(n_265),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_223),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_296),
.A2(n_279),
.B(n_282),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_307),
.B(n_308),
.Y(n_310)
);

OAI21x1_ASAP7_75t_SL g307 ( 
.A1(n_294),
.A2(n_292),
.B(n_225),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_286),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_306),
.A2(n_300),
.B(n_301),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_312),
.C(n_306),
.Y(n_313)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_305),
.B(n_297),
.CI(n_291),
.CON(n_311),
.SN(n_311)
);

NAND3xp33_ASAP7_75t_SL g314 ( 
.A(n_311),
.B(n_267),
.C(n_200),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_232),
.B1(n_197),
.B2(n_290),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g315 ( 
.A(n_313),
.B(n_314),
.CI(n_310),
.CON(n_315),
.SN(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_225),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_194),
.Y(n_317)
);


endmodule