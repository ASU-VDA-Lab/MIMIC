module real_jpeg_12148_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_2),
.Y(n_78)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_4),
.A2(n_19),
.B1(n_27),
.B2(n_31),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_4),
.A2(n_31),
.B1(n_45),
.B2(n_46),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_4),
.A2(n_6),
.B(n_27),
.C(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_4),
.B(n_19),
.C(n_38),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_4),
.A2(n_31),
.B1(n_76),
.B2(n_77),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_4),
.B(n_46),
.C(n_60),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_4),
.B(n_23),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

AO22x1_ASAP7_75t_L g23 ( 
.A1(n_6),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_8),
.A2(n_19),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_8),
.A2(n_28),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_8),
.A2(n_28),
.B1(n_76),
.B2(n_77),
.Y(n_85)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_102),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_100),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_70),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_13),
.B(n_70),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_56),
.C(n_64),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_14),
.A2(n_15),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_33),
.B1(n_54),
.B2(n_55),
.Y(n_15)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_16),
.B(n_34),
.C(n_41),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_26),
.B1(n_29),
.B2(n_32),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_18),
.B(n_30),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_21),
.Y(n_22)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_19),
.A2(n_27),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_SL g67 ( 
.A1(n_21),
.A2(n_24),
.B(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_24),
.A2(n_25),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_25),
.B(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_26),
.A2(n_32),
.B(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_31),
.B(n_42),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_31),
.B(n_97),
.Y(n_135)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OA21x2_ASAP7_75t_L g84 ( 
.A1(n_37),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_37),
.B(n_89),
.Y(n_88)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_38),
.A2(n_39),
.B1(n_76),
.B2(n_77),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_40),
.B(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_40),
.B(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_41),
.B(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B(n_49),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_46),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_42),
.A2(n_44),
.B1(n_51),
.B2(n_53),
.Y(n_81)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_50),
.Y(n_69)
);

AO22x1_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_46),
.B1(n_59),
.B2(n_60),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_45),
.B(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_56),
.A2(n_64),
.B1(n_65),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_56),
.A2(n_113),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_56),
.B(n_81),
.C(n_123),
.Y(n_140)
);

AO22x1_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_56)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_63),
.Y(n_107)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_68),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_82),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_80),
.B2(n_81),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_80),
.A2(n_81),
.B1(n_121),
.B2(n_124),
.Y(n_120)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_81),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_81),
.B(n_135),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_90),
.B2(n_91),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_94),
.B1(n_95),
.B2(n_99),
.Y(n_91)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_92),
.A2(n_99),
.B1(n_105),
.B2(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B(n_98),
.Y(n_95)
);

OA21x2_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_106),
.B(n_107),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_105),
.C(n_108),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_114),
.B(n_145),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_110),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_104),
.B(n_110),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_105),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_118),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_105),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_108),
.A2(n_109),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_139),
.B(n_144),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_125),
.B(n_138),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_120),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_118),
.Y(n_128)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_122),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_130),
.B(n_137),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_134),
.B(n_136),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_140),
.B(n_141),
.Y(n_144)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);


endmodule