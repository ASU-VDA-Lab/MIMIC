module fake_jpeg_31725_n_485 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_485);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_485;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_133;
wire n_419;
wire n_132;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_50),
.B(n_74),
.Y(n_118)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_28),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_55),
.B(n_67),
.Y(n_126)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_57),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_58),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_60),
.Y(n_152)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_75),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_20),
.B(n_15),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_79),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_81),
.B(n_83),
.Y(n_150)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_84),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_25),
.B(n_15),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_85),
.B(n_102),
.Y(n_141)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_31),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_90),
.B(n_93),
.Y(n_151)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_42),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_42),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_96),
.B(n_98),
.Y(n_153)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_18),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_17),
.Y(n_101)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_18),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_67),
.B(n_35),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_103),
.A2(n_39),
.B(n_46),
.Y(n_178)
);

INVx6_ASAP7_75t_SL g115 ( 
.A(n_72),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_115),
.Y(n_177)
);

INVx6_ASAP7_75t_SL g116 ( 
.A(n_72),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_116),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_88),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_120),
.B(n_135),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_52),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_95),
.Y(n_172)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_53),
.A2(n_17),
.B1(n_32),
.B2(n_44),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_100),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_80),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_145),
.B(n_147),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_69),
.A2(n_25),
.B(n_37),
.Y(n_146)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_32),
.B(n_44),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_71),
.Y(n_147)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_54),
.A2(n_36),
.B1(n_47),
.B2(n_29),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_35),
.B1(n_39),
.B2(n_47),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_95),
.A2(n_101),
.B1(n_43),
.B2(n_97),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_160),
.A2(n_32),
.B1(n_58),
.B2(n_102),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_99),
.B(n_20),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_29),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_119),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_162),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_152),
.A2(n_59),
.B1(n_68),
.B2(n_64),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_163),
.A2(n_114),
.B1(n_148),
.B2(n_121),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_164),
.Y(n_251)
);

AOI21xp33_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_71),
.B(n_101),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_167),
.A2(n_181),
.B(n_203),
.Y(n_257)
);

BUFx12_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_168),
.Y(n_219)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_169),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_170),
.B(n_175),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_171),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_127),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_178),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_37),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_179),
.B(n_185),
.Y(n_225)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_180),
.Y(n_231)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_183),
.A2(n_196),
.B1(n_208),
.B2(n_209),
.Y(n_224)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_49),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_119),
.A2(n_43),
.B1(n_86),
.B2(n_82),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_186),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_189),
.Y(n_229)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_104),
.Y(n_188)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_131),
.B(n_49),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_190),
.B(n_191),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_141),
.A2(n_94),
.B1(n_65),
.B2(n_76),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_118),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_192),
.B(n_198),
.Y(n_254)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_193),
.Y(n_241)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_194),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_141),
.A2(n_78),
.B1(n_63),
.B2(n_36),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_210),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_111),
.A2(n_43),
.B1(n_46),
.B2(n_36),
.Y(n_196)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_128),
.B(n_14),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_110),
.Y(n_199)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_138),
.B(n_18),
.Y(n_201)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_144),
.A2(n_32),
.B1(n_66),
.B2(n_18),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_202),
.A2(n_158),
.B(n_124),
.Y(n_240)
);

AOI21xp33_ASAP7_75t_L g203 ( 
.A1(n_144),
.A2(n_89),
.B(n_1),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_204),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_117),
.B(n_58),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_205),
.Y(n_227)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_108),
.Y(n_206)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_122),
.Y(n_207)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_106),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_114),
.A2(n_26),
.B1(n_1),
.B2(n_3),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_113),
.B(n_0),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_105),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_211),
.A2(n_214),
.B1(n_215),
.B2(n_105),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_130),
.B(n_84),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_212),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_139),
.B(n_0),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_125),
.Y(n_230)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_142),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_108),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_216),
.A2(n_240),
.B1(n_252),
.B2(n_162),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_136),
.C(n_125),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_236),
.C(n_253),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_213),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_190),
.A2(n_148),
.B1(n_133),
.B2(n_121),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_233),
.A2(n_137),
.B1(n_140),
.B2(n_211),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_180),
.B(n_112),
.C(n_134),
.Y(n_236)
);

OAI22x1_ASAP7_75t_R g242 ( 
.A1(n_202),
.A2(n_160),
.B1(n_130),
.B2(n_158),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_195),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_170),
.A2(n_175),
.B1(n_199),
.B2(n_191),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_182),
.B(n_112),
.C(n_134),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_130),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_206),
.C(n_169),
.Y(n_284)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_260),
.A2(n_240),
.B(n_266),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_284),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_222),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_267),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_220),
.B(n_173),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_264),
.B(n_271),
.Y(n_307)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_265),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_214),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_266),
.A2(n_270),
.B(n_281),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_165),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_176),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_268),
.B(n_274),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_166),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_269),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_248),
.A2(n_162),
.B1(n_177),
.B2(n_215),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_177),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_228),
.Y(n_272)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_272),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_273),
.A2(n_285),
.B1(n_222),
.B2(n_250),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_204),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_200),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_278),
.Y(n_314)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_237),
.Y(n_276)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_276),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_218),
.Y(n_277)
);

BUFx4f_ASAP7_75t_SL g294 ( 
.A(n_277),
.Y(n_294)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_231),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_235),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_279),
.A2(n_289),
.B1(n_292),
.B2(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_231),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_280),
.B(n_282),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_174),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_232),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_226),
.B(n_174),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_287),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_255),
.A2(n_133),
.B1(n_140),
.B2(n_137),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_248),
.A2(n_194),
.B1(n_188),
.B2(n_193),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_286),
.A2(n_270),
.B(n_273),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_226),
.B(n_217),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_232),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_291),
.Y(n_321)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_228),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_290),
.A2(n_171),
.B1(n_250),
.B2(n_234),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_226),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_242),
.A2(n_187),
.B1(n_159),
.B2(n_207),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_244),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_296),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_262),
.B(n_221),
.C(n_253),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_299),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_274),
.C(n_261),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_287),
.A2(n_257),
.B(n_242),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_301),
.A2(n_286),
.B(n_285),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_268),
.B(n_217),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_303),
.B(n_304),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_266),
.A2(n_224),
.B(n_236),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_254),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_323),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_308),
.A2(n_309),
.B1(n_319),
.B2(n_305),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_311),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_R g312 ( 
.A(n_291),
.B(n_238),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_312),
.A2(n_305),
.B(n_321),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_281),
.A2(n_238),
.B(n_223),
.Y(n_316)
);

A2O1A1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_316),
.A2(n_322),
.B(n_312),
.C(n_301),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_260),
.A2(n_227),
.B1(n_247),
.B2(n_234),
.Y(n_319)
);

A2O1A1O1Ixp25_ASAP7_75t_L g322 ( 
.A1(n_281),
.A2(n_249),
.B(n_219),
.C(n_187),
.D(n_168),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_265),
.B(n_249),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_276),
.B(n_244),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_288),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_326),
.A2(n_330),
.B1(n_350),
.B2(n_324),
.Y(n_368)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_328),
.Y(n_358)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_315),
.Y(n_329)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_329),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_308),
.A2(n_258),
.B1(n_290),
.B2(n_278),
.Y(n_330)
);

INVx13_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_342),
.Y(n_369)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_323),
.Y(n_332)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_332),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_334),
.B(n_339),
.Y(n_378)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_302),
.Y(n_335)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_335),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_337),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_325),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_338),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_264),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_314),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_343),
.A2(n_296),
.B(n_317),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_307),
.B(n_251),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_344),
.B(n_352),
.Y(n_373)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_345),
.Y(n_372)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_302),
.Y(n_346)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_346),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_321),
.B(n_282),
.Y(n_347)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_347),
.Y(n_382)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_320),
.Y(n_348)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_348),
.Y(n_367)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_320),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_351),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_309),
.A2(n_258),
.B1(n_280),
.B2(n_289),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_314),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_310),
.B(n_251),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_300),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_353),
.Y(n_364)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_297),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_355),
.Y(n_370)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_297),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_351),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_379),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_336),
.B(n_295),
.C(n_298),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_361),
.B(n_366),
.C(n_333),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_295),
.C(n_299),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_368),
.A2(n_331),
.B1(n_294),
.B2(n_243),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_371),
.A2(n_355),
.B(n_354),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_330),
.A2(n_258),
.B1(n_311),
.B2(n_317),
.Y(n_374)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_374),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_319),
.Y(n_376)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_327),
.A2(n_304),
.B1(n_322),
.B2(n_316),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_377),
.A2(n_380),
.B1(n_383),
.B2(n_349),
.Y(n_391)
);

AO22x2_ASAP7_75t_L g379 ( 
.A1(n_327),
.A2(n_318),
.B1(n_272),
.B2(n_294),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_328),
.A2(n_306),
.B1(n_303),
.B2(n_318),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_340),
.B(n_313),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_243),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_329),
.A2(n_313),
.B1(n_279),
.B2(n_259),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_368),
.A2(n_332),
.B1(n_338),
.B2(n_341),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_385),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_362),
.A2(n_341),
.B1(n_326),
.B2(n_350),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_386),
.B(n_387),
.C(n_389),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_333),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_366),
.B(n_334),
.C(n_345),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_380),
.B(n_343),
.C(n_337),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_390),
.B(n_395),
.C(n_400),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_391),
.B(n_398),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_378),
.A2(n_348),
.B1(n_346),
.B2(n_335),
.Y(n_392)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_392),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_393),
.A2(n_397),
.B(n_370),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_394),
.A2(n_375),
.B1(n_365),
.B2(n_367),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_277),
.Y(n_395)
);

INVx13_ASAP7_75t_L g396 ( 
.A(n_369),
.Y(n_396)
);

INVxp33_ASAP7_75t_L g420 ( 
.A(n_396),
.Y(n_420)
);

OA21x2_ASAP7_75t_L g397 ( 
.A1(n_376),
.A2(n_294),
.B(n_187),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_364),
.A2(n_293),
.B1(n_241),
.B2(n_218),
.Y(n_399)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_399),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_241),
.C(n_184),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_363),
.B(n_377),
.C(n_360),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_401),
.B(n_404),
.C(n_406),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_373),
.B(n_3),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_403),
.B(n_365),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_363),
.B(n_168),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_129),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_388),
.A2(n_359),
.B1(n_358),
.B2(n_356),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_407),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_405),
.A2(n_382),
.B1(n_356),
.B2(n_360),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_409),
.A2(n_412),
.B1(n_419),
.B2(n_385),
.Y(n_428)
);

XOR2x2_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_382),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_410),
.B(n_424),
.C(n_400),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_414),
.B(n_415),
.Y(n_432)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_384),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_417),
.A2(n_4),
.B(n_5),
.Y(n_440)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_402),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_418),
.B(n_397),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_406),
.A2(n_372),
.B1(n_379),
.B2(n_375),
.Y(n_419)
);

A2O1A1Ixp33_ASAP7_75t_L g421 ( 
.A1(n_390),
.A2(n_372),
.B(n_370),
.C(n_379),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_421),
.A2(n_419),
.B(n_397),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_386),
.B(n_367),
.C(n_379),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_428),
.Y(n_443)
);

INVx13_ASAP7_75t_L g427 ( 
.A(n_420),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_435),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_420),
.B(n_401),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_430),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_431),
.A2(n_439),
.B(n_440),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_412),
.A2(n_394),
.B1(n_389),
.B2(n_379),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_433),
.A2(n_425),
.B1(n_422),
.B2(n_410),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_404),
.Y(n_435)
);

FAx1_ASAP7_75t_SL g436 ( 
.A(n_425),
.B(n_395),
.CI(n_387),
.CON(n_436),
.SN(n_436)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_436),
.B(n_423),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_424),
.B(n_396),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_437),
.B(n_416),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_164),
.C(n_197),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_416),
.C(n_408),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_417),
.B(n_3),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g444 ( 
.A1(n_433),
.A2(n_411),
.B1(n_413),
.B2(n_421),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_444),
.A2(n_448),
.B1(n_132),
.B2(n_26),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_445),
.B(n_436),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_446),
.B(n_434),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_447),
.B(n_132),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_426),
.B(n_423),
.C(n_422),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_449),
.B(n_453),
.C(n_436),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_438),
.A2(n_129),
.B(n_123),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_450),
.A2(n_451),
.B(n_439),
.Y(n_458)
);

NOR2xp67_ASAP7_75t_SL g451 ( 
.A(n_429),
.B(n_159),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_123),
.Y(n_453)
);

OAI21x1_ASAP7_75t_L g468 ( 
.A1(n_454),
.A2(n_462),
.B(n_4),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_455),
.B(n_457),
.Y(n_469)
);

AO21x1_ASAP7_75t_L g456 ( 
.A1(n_441),
.A2(n_431),
.B(n_430),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_456),
.B(n_458),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_441),
.A2(n_432),
.B1(n_434),
.B2(n_439),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_459),
.A2(n_448),
.B1(n_452),
.B2(n_443),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_445),
.B(n_428),
.C(n_435),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_460),
.B(n_461),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_427),
.C(n_440),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_463),
.B(n_453),
.Y(n_466)
);

OA21x2_ASAP7_75t_SL g464 ( 
.A1(n_457),
.A2(n_442),
.B(n_449),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_464),
.B(n_460),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_465),
.B(n_468),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_466),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_471),
.A2(n_470),
.B(n_467),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_467),
.B(n_461),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_472),
.B(n_475),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_469),
.B(n_456),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_473),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_477),
.B(n_478),
.Y(n_479)
);

AOI322xp5_ASAP7_75t_L g480 ( 
.A1(n_476),
.A2(n_474),
.A3(n_466),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_5),
.Y(n_480)
);

AO221x1_ASAP7_75t_L g481 ( 
.A1(n_480),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_481),
.Y(n_482)
);

OAI321xp33_ASAP7_75t_L g483 ( 
.A1(n_482),
.A2(n_479),
.A3(n_10),
.B1(n_12),
.B2(n_13),
.C(n_9),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_483),
.B(n_9),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_484),
.A2(n_9),
.B(n_12),
.Y(n_485)
);


endmodule