module fake_jpeg_28688_n_403 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_403);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_403;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx2_ASAP7_75t_SL g112 ( 
.A(n_46),
.Y(n_112)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_51),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_22),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_23),
.B(n_7),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_54),
.Y(n_85)
);

BUFx2_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_64),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_7),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_63),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_27),
.B(n_41),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_67),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_27),
.B(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_69),
.B(n_70),
.Y(n_127)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_38),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_72),
.B(n_73),
.Y(n_129)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_33),
.B(n_8),
.C(n_12),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_18),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_80),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_16),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_35),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_40),
.B(n_42),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_88),
.B(n_115),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_45),
.A2(n_43),
.B1(n_18),
.B2(n_16),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_93),
.A2(n_31),
.B1(n_24),
.B2(n_0),
.Y(n_154)
);

AO22x2_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_43),
.B1(n_34),
.B2(n_28),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_42),
.B1(n_40),
.B2(n_36),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_30),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_99),
.B(n_103),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_46),
.B(n_30),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_46),
.B(n_41),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_105),
.B(n_128),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_83),
.A2(n_38),
.B1(n_25),
.B2(n_34),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_108),
.A2(n_114),
.B1(n_120),
.B2(n_125),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_49),
.A2(n_38),
.B1(n_25),
.B2(n_34),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_60),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_55),
.A2(n_25),
.B1(n_28),
.B2(n_43),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_37),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_37),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_31),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_75),
.A2(n_18),
.B1(n_28),
.B2(n_16),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_80),
.B(n_20),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_81),
.B1(n_68),
.B2(n_59),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_131),
.A2(n_143),
.B1(n_87),
.B2(n_86),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_132),
.B(n_145),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_133),
.B(n_147),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_24),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_134),
.B(n_165),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_79),
.B(n_62),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_135),
.A2(n_171),
.B(n_1),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_84),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_136),
.B(n_142),
.Y(n_192)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_137),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_95),
.A2(n_36),
.B1(n_65),
.B2(n_58),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_35),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_129),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_125),
.A2(n_57),
.B1(n_65),
.B2(n_58),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_80),
.C(n_31),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_152),
.C(n_156),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_100),
.A2(n_31),
.B1(n_24),
.B2(n_35),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_21),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_91),
.B(n_21),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_155),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_150),
.B(n_163),
.Y(n_208)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_112),
.B(n_109),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_154),
.A2(n_86),
.B1(n_110),
.B2(n_118),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_89),
.B(n_9),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_24),
.C(n_31),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_126),
.Y(n_159)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_98),
.A2(n_24),
.B1(n_9),
.B2(n_3),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_161),
.A2(n_167),
.B1(n_119),
.B2(n_102),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_89),
.B(n_6),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_96),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_89),
.B(n_90),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_114),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_109),
.A2(n_3),
.B1(n_4),
.B2(n_11),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_90),
.B(n_0),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_113),
.Y(n_207)
);

O2A1O1Ixp33_ASAP7_75t_SL g171 ( 
.A1(n_108),
.A2(n_0),
.B(n_1),
.C(n_4),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_97),
.B(n_11),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_175),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_120),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_178),
.Y(n_233)
);

BUFx12_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_193),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_102),
.B1(n_119),
.B2(n_87),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_185),
.A2(n_167),
.B1(n_141),
.B2(n_144),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_165),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_186),
.B(n_205),
.Y(n_225)
);

BUFx12_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_206),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_138),
.Y(n_198)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_137),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_201),
.A2(n_213),
.B1(n_217),
.B2(n_147),
.Y(n_243)
);

OA21x2_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_135),
.B(n_171),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_152),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_210),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_134),
.B(n_118),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_142),
.B(n_107),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_212),
.B(n_214),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_175),
.A2(n_161),
.B1(n_154),
.B2(n_132),
.Y(n_213)
);

AND2x6_ASAP7_75t_L g214 ( 
.A(n_157),
.B(n_107),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_152),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_172),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_172),
.A2(n_110),
.B1(n_97),
.B2(n_117),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_145),
.C(n_146),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_218),
.B(n_246),
.C(n_250),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_232),
.Y(n_255)
);

OAI32xp33_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_150),
.A3(n_168),
.B1(n_169),
.B2(n_132),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_222),
.B(n_196),
.Y(n_283)
);

AO21x2_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_171),
.B(n_164),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_223),
.A2(n_237),
.B(n_201),
.Y(n_267)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

AO21x1_ASAP7_75t_L g231 ( 
.A1(n_184),
.A2(n_145),
.B(n_132),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g282 ( 
.A1(n_231),
.A2(n_253),
.B(n_188),
.Y(n_282)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_181),
.B(n_136),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_235),
.B(n_239),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_170),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_244),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_143),
.B(n_159),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_191),
.Y(n_238)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_238),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_163),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_243),
.B1(n_195),
.B2(n_177),
.Y(n_254)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_242),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_156),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_184),
.B(n_207),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_247),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_179),
.B(n_184),
.C(n_189),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_160),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_151),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_211),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_189),
.B(n_176),
.C(n_117),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_211),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_190),
.B(n_12),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_254),
.A2(n_278),
.B1(n_228),
.B2(n_223),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_241),
.Y(n_256)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_221),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_257),
.B(n_281),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_237),
.A2(n_177),
.B(n_214),
.Y(n_261)
);

AO21x1_ASAP7_75t_L g292 ( 
.A1(n_261),
.A2(n_282),
.B(n_285),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_266),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_218),
.B(n_192),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_279),
.C(n_280),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_226),
.B(n_183),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_267),
.A2(n_219),
.B(n_223),
.Y(n_300)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_224),
.Y(n_269)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_226),
.B(n_183),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_275),
.Y(n_303)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_230),
.Y(n_272)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_272),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_236),
.B(n_209),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_228),
.A2(n_209),
.B1(n_194),
.B2(n_200),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_215),
.C(n_178),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_245),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_220),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_247),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g284 ( 
.A(n_241),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_180),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_227),
.A2(n_215),
.B(n_188),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_287),
.B(n_290),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_289),
.A2(n_297),
.B1(n_298),
.B2(n_304),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_273),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_250),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_299),
.C(n_301),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_260),
.B(n_222),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_296),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_262),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_263),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_254),
.A2(n_228),
.B1(n_240),
.B2(n_225),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_268),
.B(n_231),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_300),
.A2(n_267),
.B(n_255),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_249),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_302),
.A2(n_285),
.B1(n_282),
.B2(n_262),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_266),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_284),
.A2(n_223),
.B1(n_233),
.B2(n_230),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_305),
.A2(n_307),
.B1(n_278),
.B2(n_260),
.Y(n_325)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_306),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_271),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_264),
.B(n_223),
.C(n_219),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_261),
.C(n_255),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_253),
.Y(n_309)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_255),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_327),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_323),
.Y(n_339)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_288),
.Y(n_320)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_321),
.A2(n_303),
.B(n_294),
.Y(n_344)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_322),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_279),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_253),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_324),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_325),
.A2(n_302),
.B(n_308),
.Y(n_334)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_310),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_328),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_259),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_311),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_329),
.A2(n_297),
.B1(n_307),
.B2(n_304),
.Y(n_335)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_311),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_332),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_301),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_292),
.Y(n_342)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_293),
.Y(n_332)
);

XNOR2x2_ASAP7_75t_L g333 ( 
.A(n_292),
.B(n_259),
.Y(n_333)
);

AOI21xp33_ASAP7_75t_L g336 ( 
.A1(n_333),
.A2(n_295),
.B(n_309),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_334),
.A2(n_344),
.B(n_329),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_335),
.A2(n_312),
.B1(n_344),
.B2(n_317),
.Y(n_358)
);

OAI21xp33_ASAP7_75t_L g360 ( 
.A1(n_336),
.A2(n_318),
.B(n_316),
.Y(n_360)
);

NOR3xp33_ASAP7_75t_SL g338 ( 
.A(n_324),
.B(n_290),
.C(n_292),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_338),
.B(n_348),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_333),
.Y(n_340)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_340),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_346),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_293),
.Y(n_345)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_345),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_303),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_294),
.C(n_269),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_337),
.C(n_346),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_315),
.B(n_265),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_258),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_350),
.B(n_314),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_353),
.B(n_361),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_343),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_358),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_340),
.B(n_321),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_356),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_360),
.B(n_363),
.Y(n_367)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_352),
.Y(n_362)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_362),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_351),
.A2(n_327),
.B1(n_313),
.B2(n_277),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_355),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_341),
.A2(n_276),
.B(n_274),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_365),
.B(n_349),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_359),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_371),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_366),
.B(n_347),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_363),
.B(n_339),
.C(n_350),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_372),
.B(n_339),
.C(n_361),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_375),
.Y(n_387)
);

AOI21x1_ASAP7_75t_L g377 ( 
.A1(n_356),
.A2(n_334),
.B(n_338),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_377),
.A2(n_357),
.B(n_337),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_381),
.C(n_385),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_364),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_382),
.Y(n_394)
);

NAND2x1p5_ASAP7_75t_L g380 ( 
.A(n_377),
.B(n_342),
.Y(n_380)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_380),
.Y(n_388)
);

XNOR2x1_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_357),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_376),
.A2(n_354),
.B(n_360),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_270),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_383),
.Y(n_390)
);

AOI31xp33_ASAP7_75t_L g389 ( 
.A1(n_384),
.A2(n_376),
.A3(n_372),
.B(n_373),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_272),
.Y(n_385)
);

NAND3xp33_ASAP7_75t_L g395 ( 
.A(n_389),
.B(n_381),
.C(n_380),
.Y(n_395)
);

NAND3xp33_ASAP7_75t_L g391 ( 
.A(n_386),
.B(n_233),
.C(n_14),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_391),
.A2(n_193),
.B(n_394),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_378),
.B(n_198),
.C(n_180),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_393),
.B(n_390),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_395),
.B(n_396),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_392),
.B(n_387),
.C(n_193),
.Y(n_396)
);

AOI21x1_ASAP7_75t_L g400 ( 
.A1(n_397),
.A2(n_398),
.B(n_391),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_400),
.B(n_388),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_401),
.B(n_399),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_402),
.Y(n_403)
);


endmodule