module fake_jpeg_10483_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_35),
.Y(n_49)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_42),
.B(n_44),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_19),
.B1(n_28),
.B2(n_24),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_35),
.B1(n_28),
.B2(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_54),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_35),
.B1(n_22),
.B2(n_24),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_28),
.B1(n_24),
.B2(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_43),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_18),
.B1(n_34),
.B2(n_33),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_18),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_64),
.B(n_37),
.Y(n_90)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_70),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_26),
.B1(n_17),
.B2(n_32),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_31),
.B1(n_44),
.B2(n_42),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_30),
.C(n_20),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_26),
.B1(n_17),
.B2(n_21),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_38),
.A2(n_27),
.B1(n_21),
.B2(n_29),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_0),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_73),
.Y(n_110)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_78),
.B(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_79),
.B(n_81),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_44),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_44),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_87),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g132 ( 
.A(n_83),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_86),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_39),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_1),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_96),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_90),
.A2(n_45),
.B(n_30),
.Y(n_127)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_92),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_99),
.B1(n_107),
.B2(n_109),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_38),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_97),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_1),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_48),
.A2(n_40),
.B1(n_27),
.B2(n_21),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_57),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_101),
.Y(n_130)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_50),
.Y(n_104)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_65),
.B(n_12),
.Y(n_105)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

BUFx16f_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_45),
.C(n_40),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_136),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_45),
.Y(n_115)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_116),
.B(n_127),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_82),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_46),
.B1(n_40),
.B2(n_67),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_135),
.B1(n_92),
.B2(n_93),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_98),
.A2(n_40),
.B1(n_67),
.B2(n_62),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_107),
.B1(n_109),
.B2(n_47),
.Y(n_146)
);

OR2x2_ASAP7_75t_SL g131 ( 
.A(n_84),
.B(n_45),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_131),
.B(n_74),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_90),
.A2(n_47),
.B1(n_30),
.B2(n_29),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_72),
.A2(n_30),
.B(n_20),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_137),
.A2(n_108),
.B1(n_30),
.B2(n_95),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_139),
.B(n_143),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_76),
.Y(n_140)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_140),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_141),
.Y(n_184)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_78),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_80),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_145),
.B(n_147),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_154),
.B1(n_112),
.B2(n_123),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_71),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_85),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_148),
.B(n_149),
.Y(n_201)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_150),
.A2(n_160),
.B(n_164),
.Y(n_174)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_153),
.Y(n_177)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_74),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_157),
.Y(n_195)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_106),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_115),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_159),
.A2(n_161),
.B1(n_163),
.B2(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

NOR2x1_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_106),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_162),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_133),
.B(n_108),
.Y(n_165)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_134),
.Y(n_166)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_120),
.B(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_115),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_168),
.A2(n_170),
.B(n_171),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_113),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_135),
.Y(n_171)
);

AOI21x1_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_127),
.B(n_114),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_172),
.A2(n_178),
.B(n_202),
.Y(n_228)
);

OAI22x1_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_118),
.B1(n_119),
.B2(n_112),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_173),
.A2(n_181),
.B1(n_132),
.B2(n_95),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_116),
.B(n_117),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_120),
.C(n_116),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_196),
.C(n_199),
.Y(n_213)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_186),
.B(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_188),
.B(n_189),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_141),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_155),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_177),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_162),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_197),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_117),
.C(n_129),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_144),
.B(n_129),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_125),
.B(n_134),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_150),
.B(n_27),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_143),
.C(n_164),
.Y(n_223)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_211),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_201),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_205),
.B(n_218),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_156),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_207),
.C(n_223),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_156),
.Y(n_207)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_216),
.Y(n_232)
);

OAI321xp33_ASAP7_75t_L g215 ( 
.A1(n_173),
.A2(n_171),
.A3(n_139),
.B1(n_153),
.B2(n_157),
.C(n_152),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_217),
.A3(n_175),
.B1(n_188),
.B2(n_182),
.C1(n_180),
.C2(n_187),
.Y(n_234)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

NOR4xp25_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_163),
.C(n_149),
.D(n_151),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_202),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_222),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_176),
.B(n_186),
.Y(n_221)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_160),
.Y(n_224)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_226),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_169),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_185),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_227),
.A2(n_132),
.B1(n_30),
.B2(n_29),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_179),
.A2(n_125),
.B(n_123),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_175),
.B(n_192),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_181),
.B1(n_180),
.B2(n_194),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_191),
.C(n_196),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_235),
.C(n_240),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_234),
.B(n_9),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_179),
.C(n_199),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_178),
.C(n_203),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_242),
.A2(n_243),
.B1(n_246),
.B2(n_236),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_197),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_248),
.Y(n_253)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_228),
.A3(n_219),
.B1(n_211),
.B2(n_216),
.C1(n_212),
.C2(n_220),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_229),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_230),
.A2(n_128),
.B1(n_88),
.B2(n_104),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_246),
.A2(n_251),
.B1(n_214),
.B2(n_209),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_103),
.C(n_57),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_208),
.A2(n_89),
.B1(n_83),
.B2(n_57),
.Y(n_250)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_250),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_210),
.A2(n_25),
.B1(n_3),
.B2(n_4),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_204),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_269),
.Y(n_275)
);

O2A1O1Ixp33_ASAP7_75t_L g285 ( 
.A1(n_256),
.A2(n_257),
.B(n_264),
.C(n_265),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_243),
.A2(n_221),
.B1(n_226),
.B2(n_223),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_214),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_267),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_262),
.Y(n_284)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_263),
.B(n_270),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_238),
.A2(n_225),
.B1(n_3),
.B2(n_4),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_25),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_242),
.A2(n_10),
.B1(n_14),
.B2(n_7),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_268),
.A2(n_11),
.B1(n_14),
.B2(n_7),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_251),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_232),
.B(n_9),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_261),
.A2(n_238),
.B1(n_241),
.B2(n_235),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_272),
.A2(n_2),
.B1(n_4),
.B2(n_11),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_233),
.C(n_240),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_278),
.C(n_280),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_237),
.B1(n_248),
.B2(n_250),
.Y(n_277)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_244),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_9),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_257),
.B(n_8),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_286),
.B(n_12),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_276),
.A2(n_262),
.B(n_256),
.Y(n_287)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_264),
.Y(n_288)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

OAI211xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_255),
.B(n_258),
.C(n_267),
.Y(n_289)
);

AO21x1_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_297),
.B(n_285),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_253),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_290),
.B(n_295),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_284),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_253),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_290),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_281),
.Y(n_295)
);

AOI21xp33_ASAP7_75t_L g297 ( 
.A1(n_275),
.A2(n_280),
.B(n_285),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_8),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_298),
.B(n_2),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_299),
.A2(n_274),
.B1(n_279),
.B2(n_282),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_293),
.B(n_15),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_304),
.Y(n_311)
);

AOI21x1_ASAP7_75t_SL g315 ( 
.A1(n_303),
.A2(n_307),
.B(n_15),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_306),
.Y(n_313)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_299),
.B(n_12),
.CI(n_14),
.CON(n_307),
.SN(n_307)
);

AO21x1_ASAP7_75t_L g309 ( 
.A1(n_305),
.A2(n_291),
.B(n_296),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_314),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_308),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_310)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

NOR3xp33_ASAP7_75t_SL g318 ( 
.A(n_312),
.B(n_306),
.C(n_2),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_307),
.A2(n_15),
.B1(n_2),
.B2(n_4),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_301),
.Y(n_319)
);

AOI21x1_ASAP7_75t_SL g320 ( 
.A1(n_318),
.A2(n_319),
.B(n_313),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_320),
.Y(n_322)
);

OAI21x1_ASAP7_75t_SL g321 ( 
.A1(n_317),
.A2(n_309),
.B(n_311),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_322),
.B(n_316),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_321),
.C(n_300),
.Y(n_324)
);


endmodule