module real_jpeg_32517_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_561, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_561;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_0),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_0),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_0),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_0),
.Y(n_332)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_0),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_1),
.B(n_62),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_1),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_1),
.B(n_260),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_1),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_1),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_1),
.B(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_1),
.B(n_451),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_1),
.Y(n_474)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_2),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_2),
.B(n_281),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_2),
.B(n_467),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_SL g497 ( 
.A(n_2),
.B(n_498),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_3),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_3),
.Y(n_559)
);

INVx2_ASAP7_75t_R g100 ( 
.A(n_4),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_4),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_4),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_4),
.B(n_278),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_4),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_4),
.B(n_338),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_5),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_6),
.Y(n_99)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_7),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_8),
.B(n_60),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_8),
.Y(n_88)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_8),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_8),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_8),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_8),
.B(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_9),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_9),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_10),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_10),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_10),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_10),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_10),
.B(n_144),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_10),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_10),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_10),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_11),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_11),
.B(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_11),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_11),
.Y(n_314)
);

AND2x2_ASAP7_75t_SL g465 ( 
.A(n_11),
.B(n_218),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_11),
.B(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_11),
.B(n_509),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_12),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_12),
.Y(n_159)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_12),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_13),
.Y(n_321)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_14),
.Y(n_85)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_14),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_15),
.B(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_15),
.A2(n_140),
.B1(n_316),
.B2(n_318),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_15),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_15),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_15),
.B(n_377),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_15),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_15),
.B(n_501),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_15),
.B(n_514),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_16),
.Y(n_181)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_16),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_38),
.Y(n_37)
);

NAND2x1_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_17),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_17),
.B(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_17),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_17),
.B(n_171),
.Y(n_170)
);

OAI211xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_187),
.B(n_554),
.C(n_558),
.Y(n_18)
);

NAND3xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_118),
.C(n_182),
.Y(n_19)
);

AOI332xp33_ASAP7_75t_L g558 ( 
.A1(n_20),
.A2(n_21),
.A3(n_119),
.B1(n_182),
.B2(n_555),
.B3(n_556),
.C1(n_559),
.C2(n_561),
.Y(n_558)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND3xp33_ASAP7_75t_L g554 ( 
.A(n_21),
.B(n_187),
.C(n_555),
.Y(n_554)
);

AO21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_76),
.B(n_117),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_22),
.B(n_76),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_54),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_24)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_25),
.B(n_66),
.C(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_25),
.A2(n_40),
.B1(n_81),
.B2(n_82),
.Y(n_129)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_28),
.Y(n_134)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_42),
.C(n_48),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_31),
.A2(n_32),
.B1(n_50),
.B2(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_31),
.B(n_216),
.C(n_219),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_32),
.B(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_36),
.A2(n_37),
.B1(n_177),
.B2(n_178),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_36),
.A2(n_37),
.B1(n_202),
.B2(n_203),
.Y(n_262)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_37),
.B(n_169),
.C(n_177),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_37),
.B(n_199),
.C(n_202),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_39),
.Y(n_260)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_39),
.Y(n_287)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_44),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVxp67_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_44),
.B(n_139),
.C(n_143),
.Y(n_138)
);

XOR2x2_ASAP7_75t_L g160 ( 
.A(n_44),
.B(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_47),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_50),
.A2(n_58),
.B1(n_65),
.B2(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_50),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_50),
.A2(n_58),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_52),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_53),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.C(n_64),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_65),
.C(n_70),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_59),
.B(n_64),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_63),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_65),
.A2(n_66),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_65),
.A2(n_66),
.B1(n_280),
.B2(n_282),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_65),
.B(n_277),
.C(n_280),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_68),
.Y(n_258)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_70),
.B(n_135),
.C(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_72),
.B(n_156),
.Y(n_212)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_74),
.Y(n_345)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_114),
.C(n_115),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_101),
.C(n_112),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_86),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_87),
.C(n_92),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_131),
.C(n_135),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_81),
.A2(n_82),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_81),
.A2(n_82),
.B1(n_291),
.B2(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_82),
.B(n_291),
.C(n_294),
.Y(n_290)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_85),
.Y(n_175)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_85),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_88),
.B(n_103),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_88),
.B(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_91),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_100),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_99),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_100),
.B(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_112),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.C(n_109),
.Y(n_101)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_106),
.B(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_106),
.B(n_170),
.C(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_106),
.B(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_108),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_108),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_108),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_109),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_115),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_SL g557 ( 
.A(n_120),
.B(n_122),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.C(n_146),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_123),
.B(n_126),
.Y(n_224)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.C(n_138),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_127),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_130),
.B(n_138),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_135),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_135),
.B(n_250),
.Y(n_335)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_137),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_137),
.Y(n_449)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_137),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_143),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_143),
.A2(n_162),
.B1(n_235),
.B2(n_361),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_146),
.A2(n_147),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_164),
.C(n_168),
.Y(n_147)
);

XNOR2x1_ASAP7_75t_SL g194 ( 
.A(n_148),
.B(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.C(n_160),
.Y(n_148)
);

XOR2x2_ASAP7_75t_L g266 ( 
.A(n_149),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OA21x2_ASAP7_75t_L g453 ( 
.A1(n_152),
.A2(n_250),
.B(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_152),
.B(n_250),
.Y(n_454)
);

OAI21xp33_ASAP7_75t_L g485 ( 
.A1(n_152),
.A2(n_250),
.B(n_454),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_153),
.A2(n_154),
.B1(n_160),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_159),
.Y(n_384)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_160),
.Y(n_268)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_162),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_168),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.C(n_173),
.Y(n_169)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_172),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_170),
.B(n_200),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_170),
.B(n_446),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_170),
.B(n_447),
.Y(n_481)
);

INVx8_ASAP7_75t_L g523 ( 
.A(n_171),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_173),
.B(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_173),
.B(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_173),
.B(n_348),
.C(n_353),
.Y(n_362)
);

OR2x2_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_181),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_183),
.B(n_556),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21x1_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_269),
.B(n_551),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_225),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_190),
.A2(n_552),
.B(n_553),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_222),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_191),
.B(n_222),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_R g191 ( 
.A(n_192),
.B(n_194),
.C(n_196),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_194),
.Y(n_227)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_206),
.C(n_210),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_198),
.A2(n_207),
.B1(n_208),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_198),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_199),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_200),
.B(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_200),
.B(n_284),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_201),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_201),
.Y(n_516)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g263 ( 
.A(n_210),
.B(n_264),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.C(n_215),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_211),
.B(n_215),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_213),
.B(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_220),
.Y(n_246)
);

INVxp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_226),
.B(n_228),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_263),
.C(n_266),
.Y(n_228)
);

XNOR2x1_ASAP7_75t_L g418 ( 
.A(n_229),
.B(n_419),
.Y(n_418)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_247),
.C(n_261),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_230),
.B(n_410),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.C(n_244),
.Y(n_230)
);

XNOR2x1_ASAP7_75t_L g402 ( 
.A(n_231),
.B(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_233),
.A2(n_234),
.B1(n_244),
.B2(n_245),
.Y(n_403)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.C(n_240),
.Y(n_234)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_235),
.Y(n_361)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_240),
.Y(n_359)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_247),
.B(n_261),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_256),
.C(n_259),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_248),
.B(n_399),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.C(n_253),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_303)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_252),
.Y(n_511)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_255),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_259),
.Y(n_400)
);

XNOR2x1_ASAP7_75t_L g419 ( 
.A(n_263),
.B(n_266),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_431),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_405),
.B(n_427),
.Y(n_270)
);

OAI21x1_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_387),
.B(n_404),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_363),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_273),
.B(n_363),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_323),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_274),
.B(n_324),
.C(n_355),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_300),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g391 ( 
.A(n_275),
.B(n_301),
.C(n_304),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_283),
.C(n_289),
.Y(n_275)
);

XOR2x2_ASAP7_75t_L g385 ( 
.A(n_276),
.B(n_386),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_280),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_283),
.B(n_290),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NOR2x1_ASAP7_75t_L g353 ( 
.A(n_288),
.B(n_354),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_288),
.B(n_449),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_288),
.B(n_526),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_291),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_293),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_294),
.B(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_297),
.Y(n_463)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_299),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_304),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_315),
.B2(n_322),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_312),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_307),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_309),
.Y(n_502)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx6_ASAP7_75t_L g452 ( 
.A(n_310),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_311),
.Y(n_529)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_312),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_314),
.B(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_315),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g395 ( 
.A(n_315),
.B(n_396),
.C(n_397),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx5_ASAP7_75t_L g475 ( 
.A(n_317),
.Y(n_475)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

OA21x2_ASAP7_75t_SL g325 ( 
.A1(n_322),
.A2(n_326),
.B(n_330),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_355),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_333),
.C(n_346),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_325),
.B(n_346),
.Y(n_365)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx4f_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_333),
.B(n_365),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_336),
.C(n_341),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_334),
.A2(n_335),
.B1(n_442),
.B2(n_443),
.Y(n_441)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_336),
.A2(n_337),
.B1(n_341),
.B2(n_342),
.Y(n_443)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XNOR2x2_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_353),
.Y(n_346)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

XOR2x2_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_362),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

MAJx2_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_358),
.C(n_362),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

MAJx2_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.C(n_385),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_364),
.B(n_435),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_367),
.B(n_385),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_372),
.C(n_373),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_369),
.B(n_439),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_372),
.A2(n_373),
.B1(n_374),
.B2(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_372),
.Y(n_440)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_380),
.C(n_382),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_375),
.A2(n_376),
.B1(n_380),
.B2(n_381),
.Y(n_489)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_382),
.B(n_489),
.Y(n_488)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_388),
.B(n_550),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_390),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_391),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_402),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_393),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_401),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_398),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_395),
.B(n_413),
.C(n_414),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_398),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_401),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_425),
.C(n_426),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_SL g431 ( 
.A(n_405),
.B(n_432),
.C(n_549),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_417),
.B1(n_420),
.B2(n_423),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_407),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g428 ( 
.A(n_407),
.B(n_418),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_407),
.B(n_418),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_411),
.C(n_415),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_409),
.B(n_415),
.Y(n_422)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_412),
.B(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_421),
.B(n_424),
.Y(n_429)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_429),
.B(n_430),
.Y(n_427)
);

AO21x2_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_455),
.B(n_548),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_436),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_434),
.B(n_436),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_441),
.C(n_444),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_437),
.A2(n_438),
.B1(n_546),
.B2(n_547),
.Y(n_545)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_438),
.B(n_542),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_SL g542 ( 
.A(n_441),
.B(n_444),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_441),
.B(n_444),
.Y(n_547)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_450),
.C(n_453),
.Y(n_444)
);

XNOR2x1_ASAP7_75t_L g483 ( 
.A(n_445),
.B(n_484),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_450),
.A2(n_453),
.B1(n_485),
.B2(n_486),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_450),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_456),
.A2(n_540),
.B(n_544),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_457),
.A2(n_491),
.B(n_539),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_482),
.Y(n_457)
);

NOR2x1_ASAP7_75t_L g539 ( 
.A(n_458),
.B(n_482),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_471),
.C(n_481),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_460),
.B(n_536),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_464),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_465),
.C(n_470),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_462),
.B(n_521),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_465),
.A2(n_466),
.B1(n_469),
.B2(n_470),
.Y(n_464)
);

CKINVDCx14_ASAP7_75t_R g469 ( 
.A(n_465),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_466),
.Y(n_470)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

AO22x1_ASAP7_75t_L g536 ( 
.A1(n_471),
.A2(n_472),
.B1(n_481),
.B2(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_476),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_473),
.A2(n_476),
.B1(n_477),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_473),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_481),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_487),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_483),
.B(n_488),
.C(n_490),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_490),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_533),
.B(n_538),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_517),
.B(n_532),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_494),
.B(n_506),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_494),
.B(n_506),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_495),
.A2(n_496),
.B1(n_503),
.B2(n_504),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_500),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_497),
.B(n_500),
.C(n_503),
.Y(n_534)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_512),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_507),
.A2(n_508),
.B1(n_512),
.B2(n_513),
.Y(n_530)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx3_ASAP7_75t_SL g509 ( 
.A(n_510),
.Y(n_509)
);

INVx8_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_518),
.A2(n_524),
.B(n_531),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_520),
.Y(n_518)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx5_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_530),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_530),
.Y(n_531)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_535),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_534),
.B(n_535),
.Y(n_538)
);

NOR2x1p5_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_543),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_543),
.B(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);


endmodule