module real_aes_8982_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_476;
wire n_599;
wire n_887;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_592;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_870;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_795;
wire n_400;
wire n_1160;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_796;
wire n_874;
wire n_1126;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_417;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_552;
wire n_590;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_859;
wire n_685;
wire n_1080;
wire n_917;
wire n_501;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1003;
wire n_749;
wire n_914;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_873;
wire n_438;
wire n_446;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1161;
wire n_686;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_837;
wire n_829;
wire n_1030;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1129;
wire n_1014;
wire n_742;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_994;
wire n_1128;
wire n_1098;
wire n_824;
wire n_992;
wire n_813;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1062;
wire n_651;
wire n_801;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1163;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1162;
wire n_762;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_459;
wire n_1172;
wire n_998;
wire n_836;
wire n_1184;
wire n_583;
wire n_414;
wire n_776;
wire n_1138;
wire n_890;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1055;
wire n_611;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_905;
wire n_878;
wire n_577;
wire n_759;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_937;
wire n_773;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_816;
wire n_625;
wire n_953;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_609;
wire n_1006;
wire n_561;
wire n_437;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1050;
wire n_426;
wire n_1134;
wire n_616;
wire n_880;
wire n_1103;
wire n_832;
wire n_1060;
wire n_1154;
wire n_632;
wire n_714;
wire n_1222;
wire n_1041;
wire n_957;
wire n_995;
wire n_1124;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1033;
wire n_1028;
wire n_727;
wire n_1083;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1191;
wire n_705;
wire n_1206;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_1101;
wire n_1076;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_1096;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_974;
wire n_857;
wire n_491;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_1021;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_408;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1198;
wire n_993;
wire n_819;
wire n_737;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_986;
wire n_451;
wire n_1037;
wire n_790;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_768;
wire n_412;
wire n_542;
wire n_1077;
wire n_1111;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1132;
wire n_843;
wire n_579;
wire n_533;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1057;
wire n_907;
wire n_1005;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_698;
wire n_587;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_483;
wire n_729;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_603;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_SL g852 ( .A1(n_0), .A2(n_58), .B1(n_853), .B2(n_855), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_1), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_2), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g602 ( .A(n_3), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_4), .A2(n_52), .B1(n_580), .B2(n_857), .Y(n_1076) );
AOI221xp5_ASAP7_75t_L g1122 ( .A1(n_5), .A2(n_13), .B1(n_905), .B2(n_1009), .C(n_1123), .Y(n_1122) );
AOI221xp5_ASAP7_75t_L g1109 ( .A1(n_6), .A2(n_282), .B1(n_1020), .B2(n_1110), .C(n_1111), .Y(n_1109) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_7), .Y(n_724) );
AO22x2_ASAP7_75t_L g434 ( .A1(n_8), .A2(n_235), .B1(n_426), .B2(n_431), .Y(n_434) );
INVx1_ASAP7_75t_L g1166 ( .A(n_8), .Y(n_1166) );
CKINVDCx20_ASAP7_75t_R g1088 ( .A(n_9), .Y(n_1088) );
CKINVDCx20_ASAP7_75t_R g1194 ( .A(n_10), .Y(n_1194) );
CKINVDCx20_ASAP7_75t_R g1219 ( .A(n_11), .Y(n_1219) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_12), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_14), .A2(n_102), .B1(n_766), .B2(n_768), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_15), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_16), .Y(n_831) );
AOI222xp33_ASAP7_75t_L g856 ( .A1(n_17), .A2(n_53), .B1(n_155), .B2(n_484), .C1(n_501), .C2(n_857), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_18), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g1211 ( .A1(n_19), .A2(n_333), .B1(n_594), .B2(n_939), .Y(n_1211) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_20), .A2(n_163), .B1(n_512), .B2(n_582), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_21), .Y(n_813) );
CKINVDCx20_ASAP7_75t_R g1069 ( .A(n_22), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_23), .A2(n_376), .B1(n_754), .B2(n_878), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_24), .A2(n_381), .B1(n_568), .B2(n_680), .Y(n_1044) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_25), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_26), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_27), .Y(n_826) );
AOI222xp33_ASAP7_75t_L g967 ( .A1(n_28), .A2(n_57), .B1(n_362), .B2(n_578), .C1(n_855), .C2(n_968), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_29), .A2(n_128), .B1(n_518), .B2(n_746), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_30), .Y(n_873) );
AO22x2_ASAP7_75t_L g436 ( .A1(n_31), .A2(n_113), .B1(n_426), .B2(n_427), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g1107 ( .A1(n_32), .A2(n_1108), .B1(n_1127), .B2(n_1128), .Y(n_1107) );
INVx1_ASAP7_75t_L g1127 ( .A(n_32), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_33), .A2(n_392), .B1(n_604), .B2(n_751), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_34), .A2(n_222), .B1(n_957), .B2(n_1023), .Y(n_1048) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_35), .A2(n_590), .B1(n_631), .B2(n_632), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_35), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_36), .A2(n_258), .B1(n_518), .B2(n_596), .Y(n_965) );
INVx1_ASAP7_75t_L g983 ( .A(n_37), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_38), .A2(n_117), .B1(n_540), .B2(n_595), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_39), .A2(n_54), .B1(n_456), .B2(n_694), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_40), .A2(n_168), .B1(n_845), .B2(n_1064), .Y(n_1063) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_41), .A2(n_288), .B1(n_420), .B2(n_437), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g1026 ( .A(n_42), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_43), .B(n_905), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g1210 ( .A(n_44), .Y(n_1210) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_45), .A2(n_204), .B1(n_594), .B2(n_596), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_46), .A2(n_308), .B1(n_491), .B2(n_513), .Y(n_811) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_47), .A2(n_230), .B1(n_487), .B2(n_491), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_48), .A2(n_352), .B1(n_525), .B2(n_992), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_49), .B(n_679), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g1190 ( .A(n_50), .Y(n_1190) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_51), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_55), .Y(n_784) );
AOI22xp33_ASAP7_75t_SL g685 ( .A1(n_56), .A2(n_396), .B1(n_547), .B2(n_686), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_59), .A2(n_760), .B1(n_794), .B2(n_795), .Y(n_759) );
INVx1_ASAP7_75t_L g794 ( .A(n_59), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_60), .A2(n_134), .B1(n_774), .B2(n_1183), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_61), .A2(n_336), .B1(n_600), .B2(n_773), .Y(n_1065) );
AOI22xp33_ASAP7_75t_SL g519 ( .A1(n_62), .A2(n_284), .B1(n_520), .B2(n_521), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_63), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_64), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_65), .A2(n_314), .B1(n_883), .B2(n_995), .Y(n_994) );
CKINVDCx20_ASAP7_75t_R g975 ( .A(n_66), .Y(n_975) );
CKINVDCx20_ASAP7_75t_R g1215 ( .A(n_67), .Y(n_1215) );
AOI22xp33_ASAP7_75t_SL g689 ( .A1(n_68), .A2(n_200), .B1(n_690), .B2(n_691), .Y(n_689) );
INVx1_ASAP7_75t_L g927 ( .A(n_69), .Y(n_927) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_70), .Y(n_607) );
CKINVDCx20_ASAP7_75t_R g1025 ( .A(n_71), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_72), .A2(n_107), .B1(n_518), .B2(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_73), .A2(n_359), .B1(n_547), .B2(n_773), .Y(n_935) );
CKINVDCx20_ASAP7_75t_R g1006 ( .A(n_74), .Y(n_1006) );
INVx1_ASAP7_75t_L g849 ( .A(n_75), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_76), .A2(n_103), .B1(n_878), .B2(n_880), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g1084 ( .A(n_77), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_78), .A2(n_261), .B1(n_677), .B2(n_729), .Y(n_1010) );
AOI222xp33_ASAP7_75t_L g577 ( .A1(n_79), .A2(n_294), .B1(n_358), .B2(n_578), .C1(n_580), .C2(n_583), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_80), .A2(n_269), .B1(n_491), .B2(n_513), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_81), .A2(n_306), .B1(n_517), .B2(n_610), .Y(n_966) );
AOI22xp33_ASAP7_75t_SL g674 ( .A1(n_82), .A2(n_330), .B1(n_501), .B2(n_584), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_83), .A2(n_226), .B1(n_584), .B2(n_855), .Y(n_900) );
INVx1_ASAP7_75t_L g416 ( .A(n_84), .Y(n_416) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_85), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g1089 ( .A(n_86), .Y(n_1089) );
CKINVDCx20_ASAP7_75t_R g1112 ( .A(n_87), .Y(n_1112) );
CKINVDCx20_ASAP7_75t_R g1186 ( .A(n_88), .Y(n_1186) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_89), .A2(n_137), .B1(n_707), .B2(n_1081), .Y(n_1080) );
AO22x2_ASAP7_75t_L g430 ( .A1(n_90), .A2(n_262), .B1(n_426), .B2(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g1163 ( .A(n_90), .Y(n_1163) );
CKINVDCx20_ASAP7_75t_R g1135 ( .A(n_91), .Y(n_1135) );
CKINVDCx20_ASAP7_75t_R g1204 ( .A(n_92), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_93), .A2(n_94), .B1(n_460), .B2(n_610), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_95), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_96), .A2(n_111), .B1(n_455), .B2(n_457), .Y(n_454) );
OA22x2_ASAP7_75t_L g800 ( .A1(n_97), .A2(n_801), .B1(n_802), .B2(n_803), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_97), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_98), .A2(n_156), .B1(n_878), .B2(n_1023), .Y(n_1022) );
AOI222xp33_ASAP7_75t_L g1126 ( .A1(n_99), .A2(n_110), .B1(n_140), .B2(n_578), .C1(n_621), .C2(n_968), .Y(n_1126) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_100), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_101), .Y(n_792) );
AOI221xp5_ASAP7_75t_L g567 ( .A1(n_104), .A2(n_348), .B1(n_568), .B2(n_569), .C(n_570), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_105), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_106), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_108), .A2(n_196), .B1(n_512), .B2(n_815), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_109), .A2(n_227), .B1(n_693), .B2(n_764), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_112), .A2(n_158), .B1(n_461), .B2(n_521), .Y(n_716) );
INVx1_ASAP7_75t_L g1167 ( .A(n_113), .Y(n_1167) );
CKINVDCx20_ASAP7_75t_R g1075 ( .A(n_114), .Y(n_1075) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_115), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_116), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_118), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_119), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_120), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g1180 ( .A(n_121), .Y(n_1180) );
CKINVDCx20_ASAP7_75t_R g1041 ( .A(n_122), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_123), .A2(n_302), .B1(n_517), .B2(n_713), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_124), .A2(n_281), .B1(n_690), .B2(n_771), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g1187 ( .A(n_125), .Y(n_1187) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_126), .A2(n_325), .B1(n_561), .B2(n_1020), .Y(n_1019) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_127), .A2(n_239), .B1(n_773), .B2(n_774), .Y(n_772) );
AOI22xp33_ASAP7_75t_SL g678 ( .A1(n_129), .A2(n_246), .B1(n_679), .B2(n_680), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_130), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_131), .B(n_1009), .Y(n_1008) );
AOI22xp33_ASAP7_75t_SL g1140 ( .A1(n_132), .A2(n_190), .B1(n_582), .B2(n_646), .Y(n_1140) );
AOI22xp33_ASAP7_75t_SL g1143 ( .A1(n_133), .A2(n_316), .B1(n_460), .B2(n_754), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_135), .A2(n_184), .B1(n_845), .B2(n_846), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_136), .A2(n_351), .B1(n_492), .B2(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_138), .A2(n_326), .B1(n_487), .B2(n_677), .Y(n_1092) );
AOI22xp33_ASAP7_75t_SL g511 ( .A1(n_139), .A2(n_343), .B1(n_512), .B2(n_513), .Y(n_511) );
AOI22xp33_ASAP7_75t_SL g1043 ( .A1(n_141), .A2(n_206), .B1(n_677), .B2(n_855), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_142), .A2(n_349), .B1(n_956), .B2(n_957), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_143), .A2(n_324), .B1(n_910), .B2(n_995), .Y(n_1178) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_144), .A2(n_327), .B1(n_693), .B2(n_694), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_145), .A2(n_211), .B1(n_525), .B2(n_911), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_146), .A2(n_219), .B1(n_449), .B2(n_766), .Y(n_916) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_147), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g1217 ( .A(n_148), .Y(n_1217) );
CKINVDCx20_ASAP7_75t_R g1125 ( .A(n_149), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_150), .B(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_151), .A2(n_216), .B1(n_420), .B2(n_748), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_152), .A2(n_250), .B1(n_540), .B2(n_840), .Y(n_839) );
CKINVDCx20_ASAP7_75t_R g1002 ( .A(n_153), .Y(n_1002) );
AND2x6_ASAP7_75t_L g401 ( .A(n_154), .B(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g1160 ( .A(n_154), .Y(n_1160) );
AOI22xp33_ASAP7_75t_SL g682 ( .A1(n_157), .A2(n_179), .B1(n_610), .B2(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_SL g1078 ( .A1(n_159), .A2(n_290), .B1(n_729), .B2(n_1079), .Y(n_1078) );
CKINVDCx20_ASAP7_75t_R g1222 ( .A(n_160), .Y(n_1222) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_161), .A2(n_188), .B1(n_443), .B2(n_517), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_162), .A2(n_272), .B1(n_455), .B2(n_655), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_164), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g1124 ( .A(n_165), .Y(n_1124) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_166), .A2(n_271), .B1(n_456), .B2(n_599), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_167), .A2(n_198), .B1(n_910), .B2(n_911), .Y(n_909) );
AOI22xp5_ASAP7_75t_SL g918 ( .A1(n_169), .A2(n_919), .B1(n_944), .B2(n_945), .Y(n_918) );
INVx1_ASAP7_75t_L g945 ( .A(n_169), .Y(n_945) );
CKINVDCx20_ASAP7_75t_R g978 ( .A(n_170), .Y(n_978) );
AOI22xp33_ASAP7_75t_SL g500 ( .A1(n_171), .A2(n_293), .B1(n_491), .B2(n_501), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g1095 ( .A(n_172), .Y(n_1095) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_173), .A2(n_399), .B(n_407), .C(n_1168), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_174), .A2(n_321), .B1(n_443), .B2(n_449), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g1139 ( .A(n_175), .B(n_568), .Y(n_1139) );
INVx1_ASAP7_75t_L g922 ( .A(n_176), .Y(n_922) );
AO22x2_ASAP7_75t_L g425 ( .A1(n_177), .A2(n_251), .B1(n_426), .B2(n_427), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g1164 ( .A(n_177), .B(n_1165), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_178), .B(n_786), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g1192 ( .A(n_180), .Y(n_1192) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_181), .A2(n_194), .B1(n_774), .B2(n_957), .Y(n_989) );
AOI22xp33_ASAP7_75t_SL g1147 ( .A1(n_182), .A2(n_268), .B1(n_825), .B2(n_1064), .Y(n_1147) );
CKINVDCx20_ASAP7_75t_R g1029 ( .A(n_183), .Y(n_1029) );
AOI211xp5_ASAP7_75t_L g1004 ( .A1(n_185), .A2(n_483), .B(n_1005), .C(n_1011), .Y(n_1004) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_186), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g1099 ( .A1(n_187), .A2(n_375), .B1(n_883), .B2(n_1100), .Y(n_1099) );
AOI22xp33_ASAP7_75t_SL g1136 ( .A1(n_189), .A2(n_279), .B1(n_513), .B2(n_584), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_191), .A2(n_199), .B1(n_525), .B2(n_838), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_192), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_193), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_195), .Y(n_866) );
CKINVDCx20_ASAP7_75t_R g1013 ( .A(n_197), .Y(n_1013) );
AOI22xp33_ASAP7_75t_SL g711 ( .A1(n_201), .A2(n_238), .B1(n_457), .B2(n_562), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g1145 ( .A1(n_202), .A2(n_215), .B1(n_457), .B2(n_1146), .Y(n_1145) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_203), .A2(n_241), .B1(n_460), .B2(n_463), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g970 ( .A1(n_205), .A2(n_971), .B1(n_996), .B2(n_997), .Y(n_970) );
INVx1_ASAP7_75t_L g996 ( .A(n_205), .Y(n_996) );
CKINVDCx20_ASAP7_75t_R g1121 ( .A(n_207), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_208), .A2(n_397), .B1(n_461), .B2(n_562), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_209), .B(n_624), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_210), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g969 ( .A(n_212), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_213), .A2(n_386), .B1(n_460), .B2(n_821), .Y(n_959) );
CKINVDCx20_ASAP7_75t_R g1039 ( .A(n_214), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_217), .A2(n_305), .B1(n_566), .B2(n_821), .Y(n_820) );
AOI22xp33_ASAP7_75t_SL g715 ( .A1(n_218), .A2(n_315), .B1(n_456), .B2(n_520), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g1142 ( .A1(n_220), .A2(n_373), .B1(n_604), .B2(n_957), .Y(n_1142) );
CKINVDCx20_ASAP7_75t_R g961 ( .A(n_221), .Y(n_961) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_223), .A2(n_265), .B1(n_517), .B2(n_518), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_224), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g1177 ( .A(n_225), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_228), .A2(n_234), .B1(n_584), .B2(n_869), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g1101 ( .A1(n_229), .A2(n_350), .B1(n_439), .B2(n_1102), .Y(n_1101) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_231), .Y(n_554) );
XNOR2x2_ASAP7_75t_L g834 ( .A(n_232), .B(n_835), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_233), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g1094 ( .A(n_236), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_237), .A2(n_365), .B1(n_566), .B2(n_838), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_240), .A2(n_283), .B1(n_939), .B2(n_942), .Y(n_938) );
OA22x2_ASAP7_75t_L g634 ( .A1(n_242), .A2(n_635), .B1(n_636), .B2(n_659), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_242), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_243), .A2(n_391), .B1(n_600), .B2(n_687), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_244), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_245), .B(n_569), .Y(n_1138) );
XNOR2x2_ASAP7_75t_L g1059 ( .A(n_247), .B(n_1060), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_248), .A2(n_384), .B1(n_463), .B2(n_1020), .Y(n_1047) );
INVx2_ASAP7_75t_L g406 ( .A(n_249), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g882 ( .A1(n_252), .A2(n_264), .B1(n_746), .B2(n_883), .Y(n_882) );
CKINVDCx20_ASAP7_75t_R g1205 ( .A(n_253), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_254), .B(n_707), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_255), .Y(n_783) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_256), .A2(n_285), .B1(n_478), .B2(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g527 ( .A1(n_257), .A2(n_393), .B1(n_461), .B2(n_463), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g1067 ( .A(n_259), .Y(n_1067) );
AOI22xp33_ASAP7_75t_SL g524 ( .A1(n_260), .A2(n_389), .B1(n_437), .B2(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_263), .A2(n_367), .B1(n_473), .B2(n_501), .Y(n_906) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_266), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g1113 ( .A(n_267), .Y(n_1113) );
CKINVDCx20_ASAP7_75t_R g622 ( .A(n_270), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_273), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_274), .A2(n_390), .B1(n_748), .B2(n_825), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_275), .A2(n_533), .B1(n_585), .B2(n_586), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_275), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_276), .A2(n_371), .B1(n_598), .B2(n_600), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_277), .B(n_903), .Y(n_902) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_278), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_280), .Y(n_639) );
OA22x2_ASAP7_75t_L g667 ( .A1(n_286), .A2(n_668), .B1(n_669), .B2(n_695), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_286), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_287), .B(n_508), .Y(n_851) );
OA22x2_ASAP7_75t_L g1031 ( .A1(n_289), .A2(n_1032), .B1(n_1033), .B2(n_1052), .Y(n_1031) );
CKINVDCx20_ASAP7_75t_R g1032 ( .A(n_289), .Y(n_1032) );
INVx1_ASAP7_75t_L g925 ( .A(n_291), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_292), .A2(n_317), .B1(n_753), .B2(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g930 ( .A(n_295), .Y(n_930) );
XNOR2xp5_ASAP7_75t_L g1169 ( .A(n_296), .B(n_1170), .Y(n_1169) );
INVx1_ASAP7_75t_L g426 ( .A(n_297), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_297), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_298), .A2(n_388), .B1(n_455), .B2(n_518), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_299), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g1195 ( .A(n_300), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1206 ( .A1(n_301), .A2(n_379), .B1(n_600), .B2(n_1183), .Y(n_1206) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_303), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g1028 ( .A(n_304), .Y(n_1028) );
AOI22xp5_ASAP7_75t_L g1200 ( .A1(n_307), .A2(n_1201), .B1(n_1223), .B2(n_1224), .Y(n_1200) );
INVx1_ASAP7_75t_L g1223 ( .A(n_307), .Y(n_1223) );
AOI221xp5_ASAP7_75t_L g1115 ( .A1(n_309), .A2(n_329), .B1(n_883), .B2(n_1116), .C(n_1119), .Y(n_1115) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_310), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_311), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g1189 ( .A(n_312), .Y(n_1189) );
CKINVDCx20_ASAP7_75t_R g1037 ( .A(n_313), .Y(n_1037) );
INVx1_ASAP7_75t_L g777 ( .A(n_318), .Y(n_777) );
CKINVDCx20_ASAP7_75t_R g1214 ( .A(n_319), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_320), .B(n_903), .Y(n_962) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_322), .Y(n_807) );
AOI22xp33_ASAP7_75t_SL g914 ( .A1(n_323), .A2(n_383), .B1(n_553), .B2(n_915), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_328), .A2(n_347), .B1(n_439), .B2(n_594), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_331), .A2(n_357), .B1(n_473), .B2(n_477), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g980 ( .A(n_332), .Y(n_980) );
INVx1_ASAP7_75t_L g405 ( .A(n_334), .Y(n_405) );
INVx1_ASAP7_75t_L g984 ( .A(n_335), .Y(n_984) );
CKINVDCx20_ASAP7_75t_R g1209 ( .A(n_337), .Y(n_1209) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_338), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g1148 ( .A(n_339), .Y(n_1148) );
INVx1_ASAP7_75t_L g402 ( .A(n_340), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g1071 ( .A(n_341), .Y(n_1071) );
CKINVDCx20_ASAP7_75t_R g1120 ( .A(n_342), .Y(n_1120) );
OA22x2_ASAP7_75t_L g494 ( .A1(n_344), .A2(n_495), .B1(n_496), .B2(n_528), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_344), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_345), .A2(n_380), .B1(n_610), .B2(n_690), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_346), .B(n_508), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g1091 ( .A(n_353), .Y(n_1091) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_354), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_355), .B(n_857), .Y(n_928) );
CKINVDCx20_ASAP7_75t_R g1072 ( .A(n_356), .Y(n_1072) );
CKINVDCx20_ASAP7_75t_R g1174 ( .A(n_360), .Y(n_1174) );
CKINVDCx20_ASAP7_75t_R g1012 ( .A(n_361), .Y(n_1012) );
CKINVDCx20_ASAP7_75t_R g899 ( .A(n_363), .Y(n_899) );
INVx1_ASAP7_75t_L g885 ( .A(n_364), .Y(n_885) );
CKINVDCx20_ASAP7_75t_R g1221 ( .A(n_366), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_368), .B(n_729), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_369), .Y(n_789) );
INVx1_ASAP7_75t_L g923 ( .A(n_370), .Y(n_923) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_372), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_374), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g1218 ( .A(n_377), .Y(n_1218) );
CKINVDCx20_ASAP7_75t_R g1181 ( .A(n_378), .Y(n_1181) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_382), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g917 ( .A(n_385), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_387), .B(n_584), .Y(n_981) );
CKINVDCx20_ASAP7_75t_R g974 ( .A(n_394), .Y(n_974) );
INVx1_ASAP7_75t_L g931 ( .A(n_395), .Y(n_931) );
INVx2_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_401), .B(n_403), .Y(n_400) );
HB1xp67_ASAP7_75t_L g1159 ( .A(n_402), .Y(n_1159) );
OA21x2_ASAP7_75t_L g1228 ( .A1(n_403), .A2(n_1158), .B(n_1229), .Y(n_1228) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_889), .B1(n_1153), .B2(n_1154), .C(n_1155), .Y(n_407) );
INVx1_ASAP7_75t_L g1153 ( .A(n_408), .Y(n_1153) );
XNOR2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_663), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_587), .B1(n_588), .B2(n_662), .Y(n_409) );
INVx1_ASAP7_75t_L g662 ( .A(n_410), .Y(n_662) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI22xp5_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_414), .B1(n_531), .B2(n_532), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_494), .B1(n_529), .B2(n_530), .Y(n_414) );
INVx2_ASAP7_75t_SL g529 ( .A(n_415), .Y(n_529) );
XNOR2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
NOR4xp75_ASAP7_75t_L g417 ( .A(n_418), .B(n_453), .C(n_465), .D(n_481), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_419), .B(n_442), .Y(n_418) );
INVxp67_ASAP7_75t_L g537 ( .A(n_420), .Y(n_537) );
INVx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx3_ASAP7_75t_L g517 ( .A(n_421), .Y(n_517) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_422), .Y(n_595) );
BUFx2_ASAP7_75t_SL g825 ( .A(n_422), .Y(n_825) );
BUFx2_ASAP7_75t_SL g1102 ( .A(n_422), .Y(n_1102) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_432), .Y(n_422) );
AND2x6_ASAP7_75t_L g439 ( .A(n_423), .B(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g456 ( .A(n_423), .B(n_448), .Y(n_456) );
AND2x6_ASAP7_75t_L g484 ( .A(n_423), .B(n_480), .Y(n_484) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_429), .Y(n_423) );
AND2x2_ASAP7_75t_L g462 ( .A(n_424), .B(n_430), .Y(n_462) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g446 ( .A(n_425), .B(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_425), .B(n_430), .Y(n_452) );
AND2x2_ASAP7_75t_L g476 ( .A(n_425), .B(n_434), .Y(n_476) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g431 ( .A(n_428), .Y(n_431) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g447 ( .A(n_430), .Y(n_447) );
INVx1_ASAP7_75t_L g490 ( .A(n_430), .Y(n_490) );
AND2x2_ASAP7_75t_L g458 ( .A(n_432), .B(n_446), .Y(n_458) );
AND2x4_ASAP7_75t_L g461 ( .A(n_432), .B(n_462), .Y(n_461) );
AND2x4_ASAP7_75t_L g464 ( .A(n_432), .B(n_451), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_432), .B(n_446), .Y(n_557) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_435), .Y(n_432) );
OR2x2_ASAP7_75t_L g441 ( .A(n_433), .B(n_436), .Y(n_441) );
AND2x2_ASAP7_75t_L g448 ( .A(n_433), .B(n_436), .Y(n_448) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g480 ( .A(n_434), .B(n_436), .Y(n_480) );
INVx1_ASAP7_75t_L g450 ( .A(n_435), .Y(n_450) );
AND2x2_ASAP7_75t_L g489 ( .A(n_435), .B(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g475 ( .A(n_436), .Y(n_475) );
INVx4_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI21xp33_ASAP7_75t_SL g643 ( .A1(n_438), .A2(n_644), .B(n_645), .Y(n_643) );
INVx2_ASAP7_75t_SL g746 ( .A(n_438), .Y(n_746) );
INVx3_ASAP7_75t_L g771 ( .A(n_438), .Y(n_771) );
INVx4_ASAP7_75t_L g1146 ( .A(n_438), .Y(n_1146) );
INVx11_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx11_ASAP7_75t_L g563 ( .A(n_439), .Y(n_563) );
AND2x4_ASAP7_75t_L g510 ( .A(n_440), .B(n_462), .Y(n_510) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g466 ( .A(n_441), .B(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g751 ( .A(n_443), .Y(n_751) );
BUFx2_ASAP7_75t_L g1183 ( .A(n_443), .Y(n_1183) );
INVx5_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx4_ASAP7_75t_L g520 ( .A(n_444), .Y(n_520) );
INVx1_ASAP7_75t_L g599 ( .A(n_444), .Y(n_599) );
INVx2_ASAP7_75t_L g687 ( .A(n_444), .Y(n_687) );
INVx3_ASAP7_75t_L g915 ( .A(n_444), .Y(n_915) );
BUFx3_ASAP7_75t_L g958 ( .A(n_444), .Y(n_958) );
INVx8_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_446), .B(n_448), .Y(n_544) );
INVx1_ASAP7_75t_L g479 ( .A(n_447), .Y(n_479) );
NAND2x1p5_ASAP7_75t_L g470 ( .A(n_448), .B(n_462), .Y(n_470) );
AND2x6_ASAP7_75t_L g506 ( .A(n_448), .B(n_462), .Y(n_506) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
NAND2x1p5_ASAP7_75t_L g572 ( .A(n_450), .B(n_476), .Y(n_572) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR2x6_ASAP7_75t_L g522 ( .A(n_452), .B(n_475), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_454), .B(n_459), .Y(n_453) );
BUFx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx6_ASAP7_75t_L g526 ( .A(n_456), .Y(n_526) );
BUFx3_ASAP7_75t_L g693 ( .A(n_456), .Y(n_693) );
BUFx3_ASAP7_75t_L g941 ( .A(n_456), .Y(n_941) );
BUFx3_ASAP7_75t_L g694 ( .A(n_457), .Y(n_694) );
BUFx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx3_ASAP7_75t_L g518 ( .A(n_458), .Y(n_518) );
BUFx3_ASAP7_75t_L g846 ( .A(n_458), .Y(n_846) );
BUFx3_ASAP7_75t_L g911 ( .A(n_458), .Y(n_911) );
HB1xp67_ASAP7_75t_L g1176 ( .A(n_460), .Y(n_1176) );
BUFx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx3_ASAP7_75t_L g566 ( .A(n_461), .Y(n_566) );
BUFx3_ASAP7_75t_L g753 ( .A(n_461), .Y(n_753) );
INVx2_ASAP7_75t_L g767 ( .A(n_461), .Y(n_767) );
BUFx6f_ASAP7_75t_L g842 ( .A(n_461), .Y(n_842) );
INVx1_ASAP7_75t_L g467 ( .A(n_462), .Y(n_467) );
BUFx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx3_ASAP7_75t_L g540 ( .A(n_464), .Y(n_540) );
BUFx3_ASAP7_75t_L g610 ( .A(n_464), .Y(n_610) );
BUFx3_ASAP7_75t_L g713 ( .A(n_464), .Y(n_713) );
BUFx2_ASAP7_75t_SL g748 ( .A(n_464), .Y(n_748) );
BUFx2_ASAP7_75t_SL g1064 ( .A(n_464), .Y(n_1064) );
BUFx3_ASAP7_75t_L g1110 ( .A(n_464), .Y(n_1110) );
OAI221xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_468), .B1(n_469), .B2(n_471), .C(n_472), .Y(n_465) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_466), .Y(n_627) );
BUFx3_ASAP7_75t_L g640 ( .A(n_466), .Y(n_640) );
INVx2_ASAP7_75t_L g779 ( .A(n_466), .Y(n_779) );
INVx2_ASAP7_75t_L g737 ( .A(n_469), .Y(n_737) );
BUFx3_ASAP7_75t_L g1007 ( .A(n_469), .Y(n_1007) );
BUFx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g630 ( .A(n_470), .Y(n_630) );
BUFx3_ASAP7_75t_L g512 ( .A(n_473), .Y(n_512) );
BUFx2_ASAP7_75t_L g646 ( .A(n_473), .Y(n_646) );
BUFx2_ASAP7_75t_L g677 ( .A(n_473), .Y(n_677) );
INVx1_ASAP7_75t_L g854 ( .A(n_473), .Y(n_854) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_476), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x4_ASAP7_75t_L g488 ( .A(n_476), .B(n_489), .Y(n_488) );
AND2x4_ASAP7_75t_L g492 ( .A(n_476), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_SL g730 ( .A(n_477), .Y(n_730) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx2_ASAP7_75t_SL g513 ( .A(n_478), .Y(n_513) );
BUFx2_ASAP7_75t_SL g855 ( .A(n_478), .Y(n_855) );
AND2x4_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g576 ( .A(n_479), .Y(n_576) );
INVx1_ASAP7_75t_L g575 ( .A(n_480), .Y(n_575) );
OAI21xp5_ASAP7_75t_SL g481 ( .A1(n_482), .A2(n_485), .B(n_486), .Y(n_481) );
OAI21xp5_ASAP7_75t_SL g498 ( .A1(n_482), .A2(n_499), .B(n_500), .Y(n_498) );
OAI21xp33_ASAP7_75t_L g809 ( .A1(n_482), .A2(n_810), .B(n_811), .Y(n_809) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx4_ASAP7_75t_L g579 ( .A(n_484), .Y(n_579) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_484), .Y(n_653) );
INVx2_ASAP7_75t_L g672 ( .A(n_484), .Y(n_672) );
INVx2_ASAP7_75t_SL g782 ( .A(n_484), .Y(n_782) );
INVx2_ASAP7_75t_L g977 ( .A(n_484), .Y(n_977) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_487), .Y(n_621) );
INVx1_ASAP7_75t_L g740 ( .A(n_487), .Y(n_740) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx4f_ASAP7_75t_SL g501 ( .A(n_488), .Y(n_501) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_488), .Y(n_582) );
BUFx2_ASAP7_75t_L g655 ( .A(n_488), .Y(n_655) );
BUFx6f_ASAP7_75t_L g815 ( .A(n_488), .Y(n_815) );
INVx1_ASAP7_75t_L g493 ( .A(n_490), .Y(n_493) );
BUFx4f_ASAP7_75t_SL g968 ( .A(n_491), .Y(n_968) );
INVx2_ASAP7_75t_L g1016 ( .A(n_491), .Y(n_1016) );
BUFx12f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_492), .Y(n_584) );
BUFx6f_ASAP7_75t_L g726 ( .A(n_492), .Y(n_726) );
INVx1_ASAP7_75t_L g530 ( .A(n_494), .Y(n_530) );
XOR2x2_ASAP7_75t_L g633 ( .A(n_494), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g528 ( .A(n_496), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_514), .Y(n_496) );
NOR2xp67_ASAP7_75t_L g497 ( .A(n_498), .B(n_502), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g502 ( .A(n_503), .B(n_507), .C(n_511), .Y(n_502) );
INVx1_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_SL g680 ( .A(n_505), .Y(n_680) );
INVx1_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g569 ( .A(n_506), .Y(n_569) );
BUFx2_ASAP7_75t_L g707 ( .A(n_506), .Y(n_707) );
BUFx4f_ASAP7_75t_L g905 ( .A(n_506), .Y(n_905) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_508), .Y(n_568) );
INVx5_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g679 ( .A(n_509), .Y(n_679) );
INVx2_ASAP7_75t_L g903 ( .A(n_509), .Y(n_903) );
INVx2_ASAP7_75t_L g1081 ( .A(n_509), .Y(n_1081) );
INVx4_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NOR2x1_ASAP7_75t_L g514 ( .A(n_515), .B(n_523), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_519), .Y(n_515) );
BUFx2_ASAP7_75t_L g764 ( .A(n_518), .Y(n_764) );
INVx1_ASAP7_75t_L g993 ( .A(n_518), .Y(n_993) );
BUFx6f_ASAP7_75t_L g773 ( .A(n_520), .Y(n_773) );
INVx2_ASAP7_75t_L g879 ( .A(n_520), .Y(n_879) );
INVx1_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
INVx6_ASAP7_75t_SL g548 ( .A(n_522), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_522), .A2(n_574), .B1(n_648), .B2(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g880 ( .A(n_522), .Y(n_880) );
INVx1_ASAP7_75t_SL g1023 ( .A(n_522), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_527), .Y(n_523) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g553 ( .A(n_526), .Y(n_553) );
INVx2_ASAP7_75t_L g604 ( .A(n_526), .Y(n_604) );
INVx2_ASAP7_75t_L g956 ( .A(n_526), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g1070 ( .A1(n_526), .A2(n_832), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g586 ( .A(n_533), .Y(n_586) );
AND4x1_ASAP7_75t_L g533 ( .A(n_534), .B(n_549), .C(n_567), .D(n_577), .Y(n_533) );
NOR2xp33_ASAP7_75t_SL g534 ( .A(n_535), .B(n_541), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_537), .B1(n_538), .B2(n_539), .Y(n_535) );
INVx2_ASAP7_75t_L g1100 ( .A(n_539), .Y(n_1100) );
OAI221xp5_ASAP7_75t_SL g1203 ( .A1(n_539), .A2(n_555), .B1(n_1204), .B2(n_1205), .C(n_1206), .Y(n_1203) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
HB1xp67_ASAP7_75t_L g995 ( .A(n_540), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B1(n_545), .B2(n_546), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g1111 ( .A1(n_543), .A2(n_1112), .B1(n_1113), .B2(n_1114), .Y(n_1111) );
BUFx2_ASAP7_75t_R g543 ( .A(n_544), .Y(n_543) );
INVxp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx2_ASAP7_75t_L g600 ( .A(n_548), .Y(n_600) );
BUFx2_ASAP7_75t_L g754 ( .A(n_548), .Y(n_754) );
BUFx4f_ASAP7_75t_SL g774 ( .A(n_548), .Y(n_774) );
BUFx2_ASAP7_75t_L g821 ( .A(n_548), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_558), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_552), .B1(n_554), .B2(n_555), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_552), .A2(n_555), .B1(n_1025), .B2(n_1026), .Y(n_1024) );
INVxp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_555), .A2(n_602), .B1(n_603), .B2(n_605), .Y(n_601) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g832 ( .A(n_556), .Y(n_832) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B1(n_564), .B2(n_565), .Y(n_558) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g1068 ( .A(n_562), .Y(n_1068) );
INVx5_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g596 ( .A(n_563), .Y(n_596) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_563), .Y(n_684) );
INVx2_ASAP7_75t_L g838 ( .A(n_563), .Y(n_838) );
INVx4_ASAP7_75t_L g910 ( .A(n_563), .Y(n_910) );
INVx2_ASAP7_75t_SL g1118 ( .A(n_563), .Y(n_1118) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_565), .A2(n_607), .B1(n_608), .B2(n_609), .Y(n_606) );
INVx1_ASAP7_75t_L g691 ( .A(n_565), .Y(n_691) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_572), .B1(n_573), .B2(n_574), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_572), .A2(n_613), .B1(n_614), .B2(n_615), .Y(n_612) );
BUFx3_ASAP7_75t_L g742 ( .A(n_572), .Y(n_742) );
INVx4_ASAP7_75t_L g791 ( .A(n_572), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_572), .A2(n_615), .B1(n_930), .B2(n_931), .Y(n_929) );
CKINVDCx16_ASAP7_75t_R g616 ( .A(n_574), .Y(n_616) );
BUFx2_ASAP7_75t_L g985 ( .A(n_574), .Y(n_985) );
OR2x6_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx2_ASAP7_75t_L g618 ( .A(n_578), .Y(n_618) );
INVx4_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx2_ASAP7_75t_L g867 ( .A(n_579), .Y(n_867) );
INVx3_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx4_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
BUFx2_ASAP7_75t_L g869 ( .A(n_582), .Y(n_869) );
INVx2_ASAP7_75t_L g1036 ( .A(n_582), .Y(n_1036) );
INVx2_ASAP7_75t_L g1191 ( .A(n_583), .Y(n_1191) );
BUFx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx2_ASAP7_75t_L g624 ( .A(n_584), .Y(n_624) );
INVx2_ASAP7_75t_L g787 ( .A(n_584), .Y(n_787) );
INVx2_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
OA22x2_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_633), .B1(n_660), .B2(n_661), .Y(n_588) );
INVx1_ASAP7_75t_L g660 ( .A(n_589), .Y(n_660) );
INVx1_ASAP7_75t_L g632 ( .A(n_590), .Y(n_632) );
AND2x2_ASAP7_75t_SL g590 ( .A(n_591), .B(n_611), .Y(n_590) );
NOR3xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_601), .C(n_606), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_597), .Y(n_592) );
BUFx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx3_ASAP7_75t_L g690 ( .A(n_595), .Y(n_690) );
BUFx6f_ASAP7_75t_L g845 ( .A(n_595), .Y(n_845) );
INVx3_ASAP7_75t_L g1021 ( .A(n_595), .Y(n_1021) );
INVx2_ASAP7_75t_L g829 ( .A(n_596), .Y(n_829) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g1114 ( .A(n_600), .Y(n_1114) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVxp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR3xp33_ASAP7_75t_SL g611 ( .A(n_612), .B(n_617), .C(n_625), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_615), .A2(n_871), .B1(n_872), .B2(n_873), .Y(n_870) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g793 ( .A(n_616), .Y(n_793) );
OAI221xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_619), .B1(n_620), .B2(n_622), .C(n_623), .Y(n_617) );
OAI221xp5_ASAP7_75t_SL g924 ( .A1(n_618), .A2(n_925), .B1(n_926), .B2(n_927), .C(n_928), .Y(n_924) );
OAI21xp33_ASAP7_75t_SL g1090 ( .A1(n_618), .A2(n_1091), .B(n_1092), .Y(n_1090) );
OAI221xp5_ASAP7_75t_L g781 ( .A1(n_620), .A2(n_782), .B1(n_783), .B2(n_784), .C(n_785), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g1011 ( .A1(n_620), .A2(n_1012), .B1(n_1013), .B2(n_1014), .Y(n_1011) );
OAI222xp33_ASAP7_75t_L g1188 ( .A1(n_620), .A2(n_1038), .B1(n_1189), .B2(n_1190), .C1(n_1191), .C2(n_1192), .Y(n_1188) );
OAI222xp33_ASAP7_75t_L g1216 ( .A1(n_620), .A2(n_723), .B1(n_1191), .B2(n_1217), .C1(n_1218), .C2(n_1219), .Y(n_1216) );
INVx2_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_SL g979 ( .A(n_621), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B1(n_628), .B2(n_629), .Y(n_625) );
INVx1_ASAP7_75t_L g734 ( .A(n_627), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_629), .A2(n_733), .B1(n_1088), .B2(n_1089), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1213 ( .A1(n_629), .A2(n_806), .B1(n_1214), .B2(n_1215), .Y(n_1213) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g642 ( .A(n_630), .Y(n_642) );
INVx1_ASAP7_75t_L g850 ( .A(n_630), .Y(n_850) );
INVx1_ASAP7_75t_L g661 ( .A(n_633), .Y(n_661) );
INVx2_ASAP7_75t_L g659 ( .A(n_636), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_650), .Y(n_636) );
NOR3xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_643), .C(n_647), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B1(n_641), .B2(n_642), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g973 ( .A1(n_640), .A2(n_736), .B1(n_974), .B2(n_975), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_642), .A2(n_777), .B1(n_778), .B2(n_780), .Y(n_776) );
OA211x2_ASAP7_75t_L g960 ( .A1(n_642), .A2(n_961), .B(n_962), .C(n_963), .Y(n_960) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_656), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx2_ASAP7_75t_L g723 ( .A(n_653), .Y(n_723) );
INVx2_ASAP7_75t_SL g1038 ( .A(n_653), .Y(n_1038) );
INVx1_ASAP7_75t_L g926 ( .A(n_655), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
XNOR2xp5_ASAP7_75t_SL g663 ( .A(n_664), .B(n_757), .Y(n_663) );
BUFx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B1(n_696), .B2(n_697), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g695 ( .A(n_669), .Y(n_695) );
NAND3x1_ASAP7_75t_L g669 ( .A(n_670), .B(n_681), .C(n_688), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_675), .Y(n_670) );
OAI21xp5_ASAP7_75t_SL g671 ( .A1(n_672), .A2(n_673), .B(n_674), .Y(n_671) );
OAI21xp5_ASAP7_75t_SL g701 ( .A1(n_672), .A2(n_702), .B(n_703), .Y(n_701) );
OAI21xp5_ASAP7_75t_SL g1074 ( .A1(n_672), .A2(n_1075), .B(n_1076), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
BUFx2_ASAP7_75t_L g1009 ( .A(n_679), .Y(n_1009) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_685), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_692), .Y(n_688) );
INVx2_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
AO22x2_ASAP7_75t_SL g697 ( .A1(n_698), .A2(n_718), .B1(n_719), .B2(n_756), .Y(n_697) );
INVx3_ASAP7_75t_L g756 ( .A(n_698), .Y(n_756) );
XOR2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_717), .Y(n_698) );
NAND2x1_ASAP7_75t_SL g699 ( .A(n_700), .B(n_709), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_704), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .C(n_708), .Y(n_704) );
NOR2x1_ASAP7_75t_L g709 ( .A(n_710), .B(n_714), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
BUFx2_ASAP7_75t_L g768 ( .A(n_713), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
XOR2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_755), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_743), .Y(n_720) );
NOR3xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_731), .C(n_738), .Y(n_721) );
OAI221xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B1(n_725), .B2(n_727), .C(n_728), .Y(n_722) );
OAI21xp5_ASAP7_75t_L g898 ( .A1(n_723), .A2(n_899), .B(n_900), .Y(n_898) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
BUFx4f_ASAP7_75t_L g857 ( .A(n_726), .Y(n_857) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B1(n_735), .B2(n_736), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g1185 ( .A1(n_733), .A2(n_736), .B1(n_1186), .B2(n_1187), .Y(n_1185) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI22xp5_ASAP7_75t_SL g805 ( .A1(n_736), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_736), .A2(n_862), .B1(n_863), .B2(n_864), .Y(n_861) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_738) );
OAI22xp33_ASAP7_75t_L g812 ( .A1(n_742), .A2(n_813), .B1(n_814), .B2(n_816), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_749), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
INVx1_ASAP7_75t_SL g827 ( .A(n_748), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_752), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_796), .B1(n_887), .B2(n_888), .Y(n_757) );
INVx2_ASAP7_75t_L g887 ( .A(n_758), .Y(n_887) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g795 ( .A(n_760), .Y(n_795) );
AND2x2_ASAP7_75t_SL g760 ( .A(n_761), .B(n_775), .Y(n_760) );
NOR2xp33_ASAP7_75t_SL g761 ( .A(n_762), .B(n_769), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_765), .Y(n_762) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g1027 ( .A1(n_767), .A2(n_1028), .B1(n_1029), .B2(n_1030), .Y(n_1027) );
INVx1_ASAP7_75t_L g1030 ( .A(n_768), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
NOR3xp33_ASAP7_75t_L g775 ( .A(n_776), .B(n_781), .C(n_788), .Y(n_775) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g806 ( .A(n_779), .Y(n_806) );
INVx1_ASAP7_75t_SL g863 ( .A(n_779), .Y(n_863) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
OAI22xp5_ASAP7_75t_SL g1093 ( .A1(n_787), .A2(n_985), .B1(n_1094), .B2(n_1095), .Y(n_1093) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_790), .B1(n_792), .B2(n_793), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_790), .A2(n_793), .B1(n_1124), .B2(n_1125), .Y(n_1123) );
OAI22xp5_ASAP7_75t_L g1193 ( .A1(n_790), .A2(n_793), .B1(n_1194), .B2(n_1195), .Y(n_1193) );
OAI22xp5_ASAP7_75t_L g1220 ( .A1(n_790), .A2(n_793), .B1(n_1221), .B2(n_1222), .Y(n_1220) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx3_ASAP7_75t_SL g872 ( .A(n_791), .Y(n_872) );
INVx1_ASAP7_75t_L g888 ( .A(n_796), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_798), .B1(n_858), .B2(n_886), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_800), .B1(n_833), .B2(n_834), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_SL g802 ( .A(n_803), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_817), .Y(n_803) );
NOR3xp33_ASAP7_75t_L g804 ( .A(n_805), .B(n_809), .C(n_812), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g921 ( .A1(n_806), .A2(n_850), .B1(n_922), .B2(n_923), .Y(n_921) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
NOR3xp33_ASAP7_75t_L g817 ( .A(n_818), .B(n_822), .C(n_828), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_824), .B1(n_826), .B2(n_827), .Y(n_822) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_830), .B1(n_831), .B2(n_832), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g1119 ( .A1(n_832), .A2(n_940), .B1(n_1120), .B2(n_1121), .Y(n_1119) );
OAI221xp5_ASAP7_75t_SL g1179 ( .A1(n_832), .A2(n_940), .B1(n_1180), .B2(n_1181), .C(n_1182), .Y(n_1179) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
NAND4xp75_ASAP7_75t_L g835 ( .A(n_836), .B(n_843), .C(n_848), .D(n_856), .Y(n_835) );
AND2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_839), .Y(n_836) );
INVx3_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx4_ASAP7_75t_L g883 ( .A(n_841), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g1066 ( .A1(n_841), .A2(n_1067), .B1(n_1068), .B2(n_1069), .Y(n_1066) );
INVx4_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
AND2x2_ASAP7_75t_L g843 ( .A(n_844), .B(n_847), .Y(n_843) );
OA211x2_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_850), .B(n_851), .C(n_852), .Y(n_848) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g1079 ( .A(n_854), .Y(n_1079) );
INVx1_ASAP7_75t_L g1040 ( .A(n_857), .Y(n_1040) );
INVx1_ASAP7_75t_L g886 ( .A(n_858), .Y(n_886) );
XOR2x2_ASAP7_75t_L g858 ( .A(n_859), .B(n_885), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_860), .B(n_874), .Y(n_859) );
NOR3xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_865), .C(n_870), .Y(n_860) );
OAI21xp33_ASAP7_75t_L g865 ( .A1(n_866), .A2(n_867), .B(n_868), .Y(n_865) );
OAI22xp5_ASAP7_75t_L g982 ( .A1(n_872), .A2(n_983), .B1(n_984), .B2(n_985), .Y(n_982) );
NOR2xp33_ASAP7_75t_L g874 ( .A(n_875), .B(n_881), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_876), .B(n_877), .Y(n_875) );
INVx3_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_882), .B(n_884), .Y(n_881) );
INVx1_ASAP7_75t_L g1154 ( .A(n_889), .Y(n_1154) );
AOI22xp5_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_1056), .B1(n_1057), .B2(n_1152), .Y(n_889) );
INVx1_ASAP7_75t_L g1152 ( .A(n_890), .Y(n_1152) );
XOR2xp5_ASAP7_75t_L g890 ( .A(n_891), .B(n_946), .Y(n_890) );
INVx4_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
XOR2x2_ASAP7_75t_L g892 ( .A(n_893), .B(n_918), .Y(n_892) );
INVx2_ASAP7_75t_SL g893 ( .A(n_894), .Y(n_893) );
INVx3_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
XOR2x2_ASAP7_75t_L g895 ( .A(n_896), .B(n_917), .Y(n_895) );
NAND2xp5_ASAP7_75t_SL g896 ( .A(n_897), .B(n_907), .Y(n_896) );
NOR2xp33_ASAP7_75t_L g897 ( .A(n_898), .B(n_901), .Y(n_897) );
NAND3xp33_ASAP7_75t_L g901 ( .A(n_902), .B(n_904), .C(n_906), .Y(n_901) );
NOR2x1_ASAP7_75t_L g907 ( .A(n_908), .B(n_913), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_909), .B(n_912), .Y(n_908) );
INVx1_ASAP7_75t_SL g1208 ( .A(n_910), .Y(n_1208) );
INVx1_ASAP7_75t_L g943 ( .A(n_911), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_914), .B(n_916), .Y(n_913) );
INVx1_ASAP7_75t_SL g944 ( .A(n_919), .Y(n_944) );
AND2x2_ASAP7_75t_SL g919 ( .A(n_920), .B(n_932), .Y(n_919) );
NOR3xp33_ASAP7_75t_L g920 ( .A(n_921), .B(n_924), .C(n_929), .Y(n_920) );
NOR2xp33_ASAP7_75t_L g932 ( .A(n_933), .B(n_936), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_934), .B(n_935), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_937), .B(n_938), .Y(n_936) );
INVx2_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx3_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
OAI22xp5_ASAP7_75t_SL g946 ( .A1(n_947), .A2(n_999), .B1(n_1000), .B2(n_1055), .Y(n_946) );
BUFx2_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g1055 ( .A(n_948), .Y(n_1055) );
OAI22xp5_ASAP7_75t_SL g948 ( .A1(n_949), .A2(n_950), .B1(n_970), .B2(n_998), .Y(n_948) );
INVx1_ASAP7_75t_SL g949 ( .A(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
XNOR2xp5_ASAP7_75t_L g1082 ( .A(n_951), .B(n_1083), .Y(n_1082) );
INVx2_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
XOR2x2_ASAP7_75t_L g952 ( .A(n_953), .B(n_969), .Y(n_952) );
NAND4xp75_ASAP7_75t_L g953 ( .A(n_954), .B(n_960), .C(n_964), .D(n_967), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_955), .B(n_959), .Y(n_954) );
INVx3_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
AND2x2_ASAP7_75t_L g964 ( .A(n_965), .B(n_966), .Y(n_964) );
INVx1_ASAP7_75t_L g998 ( .A(n_970), .Y(n_998) );
INVx2_ASAP7_75t_L g997 ( .A(n_971), .Y(n_997) );
AND2x2_ASAP7_75t_SL g971 ( .A(n_972), .B(n_986), .Y(n_971) );
NOR3xp33_ASAP7_75t_L g972 ( .A(n_973), .B(n_976), .C(n_982), .Y(n_972) );
OAI221xp5_ASAP7_75t_L g976 ( .A1(n_977), .A2(n_978), .B1(n_979), .B2(n_980), .C(n_981), .Y(n_976) );
OAI21xp5_ASAP7_75t_SL g1134 ( .A1(n_977), .A2(n_1135), .B(n_1136), .Y(n_1134) );
NOR2xp33_ASAP7_75t_L g986 ( .A(n_987), .B(n_990), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_988), .B(n_989), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_991), .B(n_994), .Y(n_990) );
INVx2_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVx1_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
AOI22xp5_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1031), .B1(n_1053), .B2(n_1054), .Y(n_1000) );
INVx2_ASAP7_75t_L g1054 ( .A(n_1001), .Y(n_1054) );
XNOR2x1_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1003), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1017), .Y(n_1003) );
OAI211xp5_ASAP7_75t_L g1005 ( .A1(n_1006), .A2(n_1007), .B(n_1008), .C(n_1010), .Y(n_1005) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx3_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
NOR3xp33_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1024), .C(n_1027), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1022), .Y(n_1018) );
INVx2_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
OAI221xp5_ASAP7_75t_SL g1173 ( .A1(n_1021), .A2(n_1174), .B1(n_1175), .B2(n_1177), .C(n_1178), .Y(n_1173) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1031), .Y(n_1053) );
INVx1_ASAP7_75t_SL g1052 ( .A(n_1033), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1045), .Y(n_1033) );
NOR2x1_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1042), .Y(n_1034) );
OAI222xp33_ASAP7_75t_L g1035 ( .A1(n_1036), .A2(n_1037), .B1(n_1038), .B2(n_1039), .C1(n_1040), .C2(n_1041), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1044), .Y(n_1042) );
NOR2xp33_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1049), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1048), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1051), .Y(n_1049) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
AOI22xp5_ASAP7_75t_L g1057 ( .A1(n_1058), .A2(n_1105), .B1(n_1150), .B2(n_1151), .Y(n_1057) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1058), .Y(n_1151) );
AOI22xp5_ASAP7_75t_L g1058 ( .A1(n_1059), .A2(n_1082), .B1(n_1103), .B2(n_1104), .Y(n_1058) );
INVx2_ASAP7_75t_L g1103 ( .A(n_1059), .Y(n_1103) );
OAI22xp5_ASAP7_75t_L g1129 ( .A1(n_1059), .A2(n_1103), .B1(n_1130), .B2(n_1131), .Y(n_1129) );
NAND2xp5_ASAP7_75t_SL g1060 ( .A(n_1061), .B(n_1073), .Y(n_1060) );
NOR3xp33_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1066), .C(n_1070), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1065), .Y(n_1062) );
NOR2xp33_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1077), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1080), .Y(n_1077) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1082), .Y(n_1104) );
XNOR2x1_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1085), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1096), .Y(n_1085) );
NOR3xp33_ASAP7_75t_L g1086 ( .A(n_1087), .B(n_1090), .C(n_1093), .Y(n_1086) );
AND4x1_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1098), .C(n_1099), .D(n_1101), .Y(n_1096) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1105), .Y(n_1150) );
OAI22xp5_ASAP7_75t_SL g1105 ( .A1(n_1106), .A2(n_1107), .B1(n_1129), .B2(n_1149), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1108), .Y(n_1128) );
AND4x1_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1115), .C(n_1122), .D(n_1126), .Y(n_1108) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1129), .Y(n_1149) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
XOR2x2_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1148), .Y(n_1131) );
NAND3x1_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1141), .C(n_1144), .Y(n_1132) );
NOR2xp33_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1137), .Y(n_1133) );
NAND3xp33_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1139), .C(n_1140), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1143), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1147), .Y(n_1144) );
INVx1_ASAP7_75t_SL g1155 ( .A(n_1156), .Y(n_1155) );
NOR2x1_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1161), .Y(n_1156) );
OR2x2_ASAP7_75t_SL g1227 ( .A(n_1157), .B(n_1162), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1160), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1158), .B(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1159), .B(n_1197), .Y(n_1229) );
CKINVDCx16_ASAP7_75t_R g1197 ( .A(n_1160), .Y(n_1197) );
CKINVDCx20_ASAP7_75t_R g1161 ( .A(n_1162), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1164), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1167), .Y(n_1165) );
OAI222xp33_ASAP7_75t_L g1168 ( .A1(n_1169), .A2(n_1196), .B1(n_1198), .B2(n_1223), .C1(n_1225), .C2(n_1228), .Y(n_1168) );
INVx1_ASAP7_75t_SL g1170 ( .A(n_1171), .Y(n_1170) );
AND2x2_ASAP7_75t_SL g1171 ( .A(n_1172), .B(n_1184), .Y(n_1171) );
NOR2xp33_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1179), .Y(n_1172) );
OAI221xp5_ASAP7_75t_SL g1207 ( .A1(n_1175), .A2(n_1208), .B1(n_1209), .B2(n_1210), .C(n_1211), .Y(n_1207) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
NOR3xp33_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1188), .C(n_1193), .Y(n_1184) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1201), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1202), .B(n_1212), .Y(n_1201) );
NOR2xp33_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1207), .Y(n_1202) );
NOR3xp33_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1216), .C(n_1220), .Y(n_1212) );
CKINVDCx20_ASAP7_75t_R g1225 ( .A(n_1226), .Y(n_1225) );
CKINVDCx20_ASAP7_75t_R g1226 ( .A(n_1227), .Y(n_1226) );
endmodule