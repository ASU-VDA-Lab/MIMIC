module fake_ibex_707_n_924 (n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_924);

input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_924;

wire n_151;
wire n_599;
wire n_822;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_153;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_412;
wire n_357;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_375;
wire n_340;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_154;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_170;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_158;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_791;
wire n_715;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_580;
wire n_543;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_849;
wire n_857;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_648;
wire n_229;
wire n_209;
wire n_472;
wire n_571;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_456;
wire n_368;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_817;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_881;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_700;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_247;
wire n_285;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_148;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_807;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_164;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_794;
wire n_260;
wire n_620;
wire n_836;
wire n_683;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_816;
wire n_874;
wire n_890;
wire n_697;
wire n_912;
wire n_921;
wire n_149;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_895;
wire n_687;
wire n_159;
wire n_231;
wire n_298;
wire n_202;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_812;
wire n_855;
wire n_649;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_23),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_12),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_63),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_104),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_53),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_47),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_73),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_118),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_67),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_55),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_107),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_20),
.Y(n_160)
);

BUFx2_ASAP7_75t_SL g161 ( 
.A(n_33),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_71),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

NOR2xp67_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_89),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_61),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_108),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_86),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_85),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_27),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_35),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_8),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_105),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_109),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_56),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_10),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_43),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_7),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_45),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_48),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_69),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_91),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_50),
.Y(n_189)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_122),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_40),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_143),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_90),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_97),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_103),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_102),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_125),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

NOR2xp67_ASAP7_75t_L g200 ( 
.A(n_62),
.B(n_70),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_28),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_119),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_74),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_3),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_120),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_128),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_124),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_66),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_94),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_47),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_137),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_18),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_35),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_123),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_135),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_0),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_14),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_8),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_145),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_19),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_44),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_126),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_87),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_4),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_130),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_110),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_21),
.B(n_72),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_17),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_33),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_64),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_93),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_101),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_18),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_23),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_57),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_88),
.B(n_31),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_147),
.Y(n_238)
);

INVxp33_ASAP7_75t_SL g239 ( 
.A(n_84),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_24),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_92),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_13),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_100),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_99),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_51),
.Y(n_245)
);

CKINVDCx11_ASAP7_75t_R g246 ( 
.A(n_45),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_116),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_60),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_17),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_5),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_16),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_140),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_176),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_220),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_174),
.Y(n_255)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_195),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_177),
.B(n_209),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g258 ( 
.A(n_195),
.Y(n_258)
);

CKINVDCx6p67_ASAP7_75t_R g259 ( 
.A(n_195),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_157),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_157),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_160),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_167),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_167),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_239),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_162),
.Y(n_269)
);

INVxp33_ASAP7_75t_SL g270 ( 
.A(n_154),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_179),
.B(n_9),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_162),
.Y(n_272)
);

AND2x4_ASAP7_75t_L g273 ( 
.A(n_173),
.B(n_10),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_167),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_171),
.B(n_11),
.Y(n_275)
);

OAI21x1_ASAP7_75t_L g276 ( 
.A1(n_170),
.A2(n_77),
.B(n_144),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g277 ( 
.A(n_173),
.B(n_12),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_191),
.Y(n_278)
);

AOI22x1_ASAP7_75t_SL g279 ( 
.A1(n_160),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_208),
.B(n_15),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_170),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_167),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_180),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_216),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_171),
.B(n_19),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_216),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_152),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_216),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_154),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_231),
.B(n_22),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_180),
.Y(n_291)
);

NOR2x1_ASAP7_75t_L g292 ( 
.A(n_234),
.B(n_54),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_187),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_233),
.B(n_24),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_152),
.Y(n_295)
);

BUFx8_ASAP7_75t_SL g296 ( 
.A(n_222),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_216),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_187),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_221),
.B(n_25),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_234),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_245),
.B(n_26),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_249),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_245),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_196),
.B(n_29),
.Y(n_304)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_151),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_150),
.Y(n_306)
);

AND2x6_ASAP7_75t_L g307 ( 
.A(n_151),
.B(n_58),
.Y(n_307)
);

BUFx8_ASAP7_75t_L g308 ( 
.A(n_185),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_196),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_185),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g311 ( 
.A(n_153),
.B(n_32),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_163),
.B(n_34),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_198),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_205),
.B(n_36),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_165),
.B(n_36),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_198),
.B(n_203),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_203),
.B(n_37),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_213),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_217),
.B(n_37),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_149),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_264),
.Y(n_321)
);

AO21x2_ASAP7_75t_L g322 ( 
.A1(n_294),
.A2(n_304),
.B(n_276),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_256),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_255),
.B(n_155),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_264),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

INVx8_ASAP7_75t_L g327 ( 
.A(n_307),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_267),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_267),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_262),
.B(n_158),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_267),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_274),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_253),
.B(n_148),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_260),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_261),
.Y(n_336)
);

AOI21x1_ASAP7_75t_L g337 ( 
.A1(n_304),
.A2(n_292),
.B(n_280),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_274),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_262),
.B(n_204),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_274),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_261),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_269),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_282),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_282),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_269),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_277),
.Y(n_347)
);

INVx8_ASAP7_75t_L g348 ( 
.A(n_307),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_272),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_286),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_270),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_286),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_272),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_311),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_288),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_311),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_281),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_281),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_297),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_283),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_257),
.B(n_244),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_307),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_283),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_SL g366 ( 
.A(n_275),
.B(n_156),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_289),
.B(n_247),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_289),
.B(n_247),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_284),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_291),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_259),
.B(n_225),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_270),
.B(n_156),
.Y(n_373)
);

NOR2x1p5_ASAP7_75t_L g374 ( 
.A(n_258),
.B(n_265),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_284),
.Y(n_375)
);

INVx5_ASAP7_75t_L g376 ( 
.A(n_284),
.Y(n_376)
);

OR2x6_ASAP7_75t_L g377 ( 
.A(n_263),
.B(n_161),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_284),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_293),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_293),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_298),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_309),
.Y(n_382)
);

BUFx6f_ASAP7_75t_SL g383 ( 
.A(n_319),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_309),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_313),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_320),
.B(n_181),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_313),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_266),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_306),
.B(n_168),
.Y(n_389)
);

BUFx10_ASAP7_75t_L g390 ( 
.A(n_285),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_308),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_312),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_271),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_290),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_308),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_300),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_302),
.Y(n_397)
);

NAND3xp33_ASAP7_75t_L g398 ( 
.A(n_285),
.B(n_183),
.C(n_182),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_318),
.B(n_178),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_317),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_299),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_278),
.B(n_184),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_314),
.Y(n_404)
);

NAND2xp33_ASAP7_75t_L g405 ( 
.A(n_305),
.B(n_207),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_315),
.Y(n_406)
);

AO21x2_ASAP7_75t_L g407 ( 
.A1(n_301),
.A2(n_237),
.B(n_228),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_268),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_303),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_254),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_279),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_295),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_296),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_296),
.Y(n_414)
);

NOR2x1p5_ASAP7_75t_L g415 ( 
.A(n_259),
.B(n_235),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_257),
.B(n_189),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_264),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_270),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_273),
.Y(n_419)
);

NAND2xp33_ASAP7_75t_L g420 ( 
.A(n_307),
.B(n_207),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_260),
.Y(n_421)
);

BUFx6f_ASAP7_75t_SL g422 ( 
.A(n_307),
.Y(n_422)
);

BUFx6f_ASAP7_75t_SL g423 ( 
.A(n_414),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_404),
.B(n_190),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_364),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_388),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_404),
.B(n_166),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_393),
.B(n_169),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_394),
.B(n_172),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_175),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_388),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_331),
.B(n_194),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_339),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_339),
.B(n_363),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_418),
.B(n_246),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_395),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_408),
.A2(n_159),
.B1(n_212),
.B2(n_215),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_416),
.B(n_201),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_408),
.A2(n_159),
.B1(n_197),
.B2(n_212),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_351),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_395),
.Y(n_441)
);

AOI221xp5_ASAP7_75t_L g442 ( 
.A1(n_409),
.A2(n_229),
.B1(n_214),
.B2(n_251),
.C(n_211),
.Y(n_442)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_416),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_403),
.B(n_223),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_403),
.B(n_224),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_391),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_391),
.B(n_227),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_351),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_367),
.B(n_369),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_410),
.A2(n_197),
.B1(n_232),
.B2(n_238),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_407),
.B(n_186),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_407),
.B(n_188),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_401),
.Y(n_453)
);

O2A1O1Ixp33_ASAP7_75t_L g454 ( 
.A1(n_410),
.A2(n_252),
.B(n_192),
.C(n_193),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_323),
.B(n_241),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_327),
.Y(n_456)
);

BUFx12f_ASAP7_75t_L g457 ( 
.A(n_415),
.Y(n_457)
);

A2O1A1Ixp33_ASAP7_75t_L g458 ( 
.A1(n_400),
.A2(n_248),
.B(n_199),
.C(n_202),
.Y(n_458)
);

NOR3xp33_ASAP7_75t_L g459 ( 
.A(n_366),
.B(n_219),
.C(n_218),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_401),
.B(n_230),
.Y(n_460)
);

OR2x6_ASAP7_75t_L g461 ( 
.A(n_413),
.B(n_242),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_402),
.B(n_240),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_347),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_392),
.B(n_206),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_355),
.B(n_210),
.Y(n_465)
);

OR2x6_ASAP7_75t_L g466 ( 
.A(n_413),
.B(n_242),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_386),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_372),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_358),
.Y(n_469)
);

INVx8_ASAP7_75t_L g470 ( 
.A(n_348),
.Y(n_470)
);

OR2x6_ASAP7_75t_L g471 ( 
.A(n_374),
.B(n_164),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_396),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_397),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_348),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_412),
.B(n_226),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_419),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_322),
.B(n_334),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_329),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_324),
.B(n_236),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_412),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_335),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_335),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_336),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_322),
.B(n_200),
.Y(n_484)
);

NOR3xp33_ASAP7_75t_L g485 ( 
.A(n_411),
.B(n_38),
.C(n_39),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_322),
.B(n_59),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_383),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_336),
.B(n_65),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_390),
.B(n_38),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_398),
.B(n_68),
.Y(n_490)
);

A2O1A1Ixp33_ASAP7_75t_L g491 ( 
.A1(n_449),
.A2(n_420),
.B(n_365),
.C(n_360),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_443),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_453),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_434),
.B(n_389),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_477),
.A2(n_405),
.B(n_399),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_467),
.B(n_383),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_424),
.B(n_341),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_460),
.B(n_377),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_435),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_468),
.A2(n_377),
.B1(n_411),
.B2(n_422),
.Y(n_500)
);

OAI21xp33_ASAP7_75t_L g501 ( 
.A1(n_438),
.A2(n_377),
.B(n_337),
.Y(n_501)
);

O2A1O1Ixp33_ASAP7_75t_L g502 ( 
.A1(n_451),
.A2(n_377),
.B(n_345),
.C(n_349),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_427),
.B(n_342),
.Y(n_503)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_456),
.B(n_422),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_451),
.A2(n_353),
.B(n_349),
.Y(n_505)
);

O2A1O1Ixp33_ASAP7_75t_L g506 ( 
.A1(n_452),
.A2(n_359),
.B(n_362),
.C(n_421),
.Y(n_506)
);

O2A1O1Ixp33_ASAP7_75t_L g507 ( 
.A1(n_452),
.A2(n_382),
.B(n_371),
.C(n_379),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_487),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_448),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_446),
.Y(n_510)
);

NOR3xp33_ASAP7_75t_L g511 ( 
.A(n_437),
.B(n_381),
.C(n_380),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_430),
.A2(n_384),
.B(n_381),
.Y(n_512)
);

O2A1O1Ixp33_ASAP7_75t_SL g513 ( 
.A1(n_488),
.A2(n_385),
.B(n_387),
.C(n_370),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_427),
.B(n_385),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_486),
.A2(n_387),
.B(n_378),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_428),
.B(n_40),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_428),
.B(n_41),
.Y(n_517)
);

O2A1O1Ixp33_ASAP7_75t_L g518 ( 
.A1(n_458),
.A2(n_454),
.B(n_433),
.C(n_429),
.Y(n_518)
);

OA22x2_ASAP7_75t_L g519 ( 
.A1(n_437),
.A2(n_42),
.B1(n_43),
.B2(n_46),
.Y(n_519)
);

AO21x1_ASAP7_75t_L g520 ( 
.A1(n_486),
.A2(n_368),
.B(n_417),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_429),
.B(n_469),
.Y(n_521)
);

AOI21x1_ASAP7_75t_L g522 ( 
.A1(n_488),
.A2(n_346),
.B(n_325),
.Y(n_522)
);

OAI21xp33_ASAP7_75t_L g523 ( 
.A1(n_444),
.A2(n_375),
.B(n_321),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_470),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_426),
.A2(n_350),
.B(n_328),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_431),
.A2(n_481),
.B(n_478),
.Y(n_526)
);

AOI33xp33_ASAP7_75t_L g527 ( 
.A1(n_442),
.A2(n_356),
.A3(n_330),
.B1(n_332),
.B2(n_333),
.B3(n_338),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_482),
.A2(n_352),
.B(n_328),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_459),
.A2(n_375),
.B1(n_376),
.B2(n_361),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_470),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_440),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_483),
.A2(n_344),
.B(n_357),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_425),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_480),
.B(n_49),
.Y(n_534)
);

NOR2x1_ASAP7_75t_R g535 ( 
.A(n_457),
.B(n_376),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_436),
.B(n_51),
.Y(n_536)
);

OAI21xp33_ASAP7_75t_L g537 ( 
.A1(n_445),
.A2(n_343),
.B(n_340),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_432),
.B(n_475),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_R g539 ( 
.A(n_441),
.B(n_52),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_463),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_439),
.B(n_53),
.Y(n_541)
);

AOI21x1_ASAP7_75t_L g542 ( 
.A1(n_490),
.A2(n_354),
.B(n_326),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_439),
.B(n_354),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_489),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_544)
);

O2A1O1Ixp33_ASAP7_75t_L g545 ( 
.A1(n_464),
.A2(n_79),
.B(n_80),
.C(n_81),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_476),
.A2(n_82),
.B(n_83),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_462),
.B(n_95),
.Y(n_547)
);

O2A1O1Ixp33_ASAP7_75t_L g548 ( 
.A1(n_465),
.A2(n_142),
.B(n_96),
.C(n_98),
.Y(n_548)
);

INVx8_ASAP7_75t_L g549 ( 
.A(n_461),
.Y(n_549)
);

OR2x6_ASAP7_75t_L g550 ( 
.A(n_466),
.B(n_111),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_447),
.B(n_138),
.Y(n_551)
);

NOR2x1_ASAP7_75t_L g552 ( 
.A(n_471),
.B(n_129),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_479),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_553)
);

INVx3_ASAP7_75t_SL g554 ( 
.A(n_471),
.Y(n_554)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_515),
.A2(n_472),
.B(n_473),
.Y(n_555)
);

OAI21xp33_ASAP7_75t_L g556 ( 
.A1(n_538),
.A2(n_541),
.B(n_517),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_516),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_494),
.B(n_485),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_519),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_498),
.B(n_455),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_531),
.Y(n_561)
);

OR2x6_ASAP7_75t_L g562 ( 
.A(n_549),
.B(n_474),
.Y(n_562)
);

BUFx12f_ASAP7_75t_L g563 ( 
.A(n_509),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_499),
.B(n_423),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_L g565 ( 
.A(n_504),
.B(n_549),
.Y(n_565)
);

AND3x4_ASAP7_75t_L g566 ( 
.A(n_552),
.B(n_536),
.C(n_551),
.Y(n_566)
);

A2O1A1Ixp33_ASAP7_75t_L g567 ( 
.A1(n_501),
.A2(n_495),
.B(n_527),
.C(n_526),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_554),
.Y(n_568)
);

OAI21x1_ASAP7_75t_L g569 ( 
.A1(n_528),
.A2(n_532),
.B(n_525),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_512),
.A2(n_507),
.B(n_506),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_500),
.B(n_496),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_537),
.A2(n_523),
.B(n_547),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_551),
.A2(n_534),
.B(n_511),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_539),
.B(n_508),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_524),
.B(n_530),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_533),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_524),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_530),
.Y(n_578)
);

NAND3xp33_ASAP7_75t_L g579 ( 
.A(n_545),
.B(n_544),
.C(n_548),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_535),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_533),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_540),
.Y(n_582)
);

NAND3xp33_ASAP7_75t_L g583 ( 
.A(n_553),
.B(n_546),
.C(n_529),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_535),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_510),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_499),
.B(n_418),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_L g587 ( 
.A(n_504),
.B(n_470),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_521),
.B(n_443),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_524),
.B(n_530),
.Y(n_589)
);

OAI22x1_ASAP7_75t_L g590 ( 
.A1(n_536),
.A2(n_450),
.B1(n_287),
.B2(n_295),
.Y(n_590)
);

OAI22x1_ASAP7_75t_L g591 ( 
.A1(n_536),
.A2(n_450),
.B1(n_287),
.B2(n_295),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g592 ( 
.A1(n_491),
.A2(n_477),
.B(n_505),
.Y(n_592)
);

OAI21x1_ASAP7_75t_L g593 ( 
.A1(n_515),
.A2(n_522),
.B(n_542),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_521),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_521),
.Y(n_595)
);

OAI21x1_ASAP7_75t_L g596 ( 
.A1(n_515),
.A2(n_522),
.B(n_542),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_513),
.A2(n_420),
.B(n_477),
.Y(n_597)
);

A2O1A1Ixp33_ASAP7_75t_L g598 ( 
.A1(n_518),
.A2(n_449),
.B(n_502),
.C(n_516),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_524),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_521),
.A2(n_503),
.B1(n_514),
.B2(n_497),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_515),
.A2(n_522),
.B(n_542),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_521),
.B(n_443),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_493),
.B(n_437),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_531),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_499),
.B(n_418),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_499),
.B(n_418),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_491),
.A2(n_477),
.B(n_505),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_L g608 ( 
.A1(n_491),
.A2(n_477),
.B(n_505),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_531),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_521),
.B(n_443),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_L g611 ( 
.A1(n_491),
.A2(n_477),
.B(n_505),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_521),
.B(n_443),
.Y(n_612)
);

AOI21xp33_ASAP7_75t_L g613 ( 
.A1(n_496),
.A2(n_418),
.B(n_443),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_492),
.B(n_418),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_L g615 ( 
.A1(n_491),
.A2(n_477),
.B(n_505),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_491),
.A2(n_477),
.B(n_505),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_493),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_492),
.Y(n_618)
);

OAI22x1_ASAP7_75t_L g619 ( 
.A1(n_536),
.A2(n_450),
.B1(n_287),
.B2(n_295),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_521),
.A2(n_503),
.B1(n_514),
.B2(n_497),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_521),
.A2(n_503),
.B1(n_514),
.B2(n_497),
.Y(n_621)
);

CKINVDCx6p67_ASAP7_75t_R g622 ( 
.A(n_554),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_493),
.Y(n_623)
);

AO21x1_ASAP7_75t_L g624 ( 
.A1(n_545),
.A2(n_484),
.B(n_477),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_491),
.A2(n_477),
.B(n_505),
.Y(n_625)
);

OR2x6_ASAP7_75t_L g626 ( 
.A(n_549),
.B(n_550),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_491),
.A2(n_477),
.B(n_505),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_521),
.B(n_443),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_493),
.B(n_443),
.Y(n_629)
);

A2O1A1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_518),
.A2(n_449),
.B(n_502),
.C(n_516),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_521),
.B(n_443),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_493),
.B(n_443),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_493),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_492),
.B(n_418),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_492),
.B(n_418),
.Y(n_635)
);

A2O1A1Ixp33_ASAP7_75t_L g636 ( 
.A1(n_518),
.A2(n_449),
.B(n_502),
.C(n_516),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_499),
.B(n_418),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_521),
.B(n_443),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_524),
.B(n_530),
.Y(n_639)
);

NOR2xp67_ASAP7_75t_L g640 ( 
.A(n_524),
.B(n_530),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_521),
.A2(n_503),
.B1(n_514),
.B2(n_497),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_521),
.B(n_443),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_493),
.B(n_443),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_524),
.B(n_530),
.Y(n_644)
);

AOI21xp33_ASAP7_75t_L g645 ( 
.A1(n_496),
.A2(n_418),
.B(n_443),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_492),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_521),
.B(n_443),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_491),
.A2(n_477),
.B(n_505),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_609),
.Y(n_649)
);

BUFx5_ASAP7_75t_L g650 ( 
.A(n_575),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_600),
.B(n_620),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_577),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_575),
.B(n_589),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_582),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_584),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_641),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_594),
.B(n_595),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g658 ( 
.A1(n_598),
.A2(n_636),
.B(n_630),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_559),
.A2(n_603),
.B1(n_566),
.B2(n_557),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_617),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_626),
.Y(n_661)
);

INVx8_ASAP7_75t_L g662 ( 
.A(n_577),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_577),
.Y(n_663)
);

AO21x2_ASAP7_75t_L g664 ( 
.A1(n_624),
.A2(n_567),
.B(n_572),
.Y(n_664)
);

AND2x6_ASAP7_75t_L g665 ( 
.A(n_576),
.B(n_581),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_626),
.Y(n_666)
);

BUFx2_ASAP7_75t_SL g667 ( 
.A(n_640),
.Y(n_667)
);

A2O1A1Ixp33_ASAP7_75t_L g668 ( 
.A1(n_556),
.A2(n_573),
.B(n_570),
.C(n_648),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g669 ( 
.A1(n_592),
.A2(n_608),
.B(n_607),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_592),
.A2(n_608),
.B(n_607),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_626),
.Y(n_671)
);

AO21x2_ASAP7_75t_L g672 ( 
.A1(n_611),
.A2(n_615),
.B(n_616),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_588),
.B(n_602),
.Y(n_673)
);

INVx8_ASAP7_75t_L g674 ( 
.A(n_639),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_571),
.A2(n_558),
.B1(n_619),
.B2(n_590),
.Y(n_675)
);

NAND2x1p5_ASAP7_75t_L g676 ( 
.A(n_644),
.B(n_640),
.Y(n_676)
);

AO21x2_ASAP7_75t_L g677 ( 
.A1(n_611),
.A2(n_625),
.B(n_627),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_627),
.A2(n_570),
.B(n_579),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_610),
.B(n_612),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_579),
.A2(n_583),
.B(n_569),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_578),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_623),
.Y(n_682)
);

INVx6_ASAP7_75t_L g683 ( 
.A(n_563),
.Y(n_683)
);

AOI22x1_ASAP7_75t_L g684 ( 
.A1(n_599),
.A2(n_560),
.B1(n_585),
.B2(n_591),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_628),
.B(n_647),
.Y(n_685)
);

CKINVDCx11_ASAP7_75t_R g686 ( 
.A(n_622),
.Y(n_686)
);

OR2x6_ASAP7_75t_L g687 ( 
.A(n_562),
.B(n_580),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_631),
.B(n_642),
.Y(n_688)
);

BUFx12f_ASAP7_75t_L g689 ( 
.A(n_568),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_638),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_629),
.B(n_632),
.Y(n_691)
);

BUFx4f_ASAP7_75t_L g692 ( 
.A(n_574),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_613),
.A2(n_645),
.B(n_587),
.Y(n_693)
);

OAI211xp5_ASAP7_75t_L g694 ( 
.A1(n_633),
.A2(n_606),
.B(n_637),
.C(n_605),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_565),
.A2(n_614),
.B(n_635),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_643),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_618),
.Y(n_697)
);

NOR2x1_ASAP7_75t_R g698 ( 
.A(n_604),
.B(n_634),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_586),
.B(n_561),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_646),
.Y(n_700)
);

INVx6_ASAP7_75t_L g701 ( 
.A(n_564),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_584),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_586),
.A2(n_437),
.B1(n_439),
.B2(n_373),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_582),
.Y(n_704)
);

OAI21xp5_ASAP7_75t_L g705 ( 
.A1(n_598),
.A2(n_636),
.B(n_630),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_600),
.A2(n_621),
.B(n_620),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_603),
.B(n_443),
.Y(n_707)
);

AO31x2_ASAP7_75t_L g708 ( 
.A1(n_567),
.A2(n_624),
.A3(n_520),
.B(n_597),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_600),
.A2(n_541),
.B1(n_543),
.B2(n_519),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_600),
.A2(n_541),
.B1(n_543),
.B2(n_519),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_600),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_576),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_594),
.B(n_443),
.Y(n_713)
);

BUFx12f_ASAP7_75t_L g714 ( 
.A(n_568),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_577),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_577),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_600),
.A2(n_541),
.B1(n_543),
.B2(n_519),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_600),
.B(n_620),
.Y(n_718)
);

BUFx6f_ASAP7_75t_SL g719 ( 
.A(n_626),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_600),
.B(n_620),
.Y(n_720)
);

OA21x2_ASAP7_75t_L g721 ( 
.A1(n_593),
.A2(n_601),
.B(n_596),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_582),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_598),
.A2(n_636),
.B(n_630),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_582),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_555),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_656),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_686),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_656),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_711),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_651),
.B(n_718),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_711),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_725),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_721),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_674),
.Y(n_734)
);

AO21x2_ASAP7_75t_L g735 ( 
.A1(n_680),
.A2(n_678),
.B(n_658),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_720),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_720),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_703),
.B(n_694),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_674),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_654),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_704),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_665),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_722),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_SL g744 ( 
.A1(n_719),
.A2(n_684),
.B1(n_661),
.B2(n_706),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_SL g745 ( 
.A1(n_719),
.A2(n_661),
.B1(n_706),
.B2(n_671),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_662),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_724),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_672),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_677),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_665),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_673),
.B(n_679),
.Y(n_751)
);

BUFx10_ASAP7_75t_L g752 ( 
.A(n_653),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_662),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_685),
.B(n_657),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_677),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_686),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_705),
.Y(n_757)
);

OA21x2_ASAP7_75t_L g758 ( 
.A1(n_668),
.A2(n_678),
.B(n_669),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_662),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_705),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_723),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_SL g762 ( 
.A1(n_666),
.A2(n_650),
.B1(n_667),
.B2(n_694),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_723),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_712),
.Y(n_764)
);

CKINVDCx6p67_ASAP7_75t_R g765 ( 
.A(n_689),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_660),
.Y(n_766)
);

BUFx2_ASAP7_75t_R g767 ( 
.A(n_655),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_664),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_733),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_730),
.B(n_670),
.Y(n_770)
);

INVxp67_ASAP7_75t_SL g771 ( 
.A(n_732),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_735),
.B(n_670),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_742),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_742),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_738),
.A2(n_659),
.B1(n_710),
.B2(n_709),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_728),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_730),
.B(n_709),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_750),
.Y(n_778)
);

OAI221xp5_ASAP7_75t_SL g779 ( 
.A1(n_754),
.A2(n_659),
.B1(n_675),
.B2(n_717),
.C(n_660),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_731),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_726),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_758),
.B(n_664),
.Y(n_782)
);

INVx5_ASAP7_75t_L g783 ( 
.A(n_764),
.Y(n_783)
);

NOR2x1_ASAP7_75t_L g784 ( 
.A(n_746),
.B(n_663),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_750),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_726),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_SL g787 ( 
.A1(n_762),
.A2(n_676),
.B(n_675),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_757),
.B(n_708),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_757),
.B(n_760),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_729),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_729),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_776),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_776),
.Y(n_793)
);

AOI221xp5_ASAP7_75t_L g794 ( 
.A1(n_779),
.A2(n_707),
.B1(n_688),
.B2(n_696),
.C(n_690),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_770),
.B(n_751),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_775),
.A2(n_761),
.B1(n_763),
.B2(n_745),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_772),
.B(n_748),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_769),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_776),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_772),
.B(n_749),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_780),
.Y(n_801)
);

INVxp67_ASAP7_75t_SL g802 ( 
.A(n_771),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_781),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_783),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_781),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_775),
.A2(n_763),
.B1(n_737),
.B2(n_736),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_772),
.B(n_755),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_784),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_770),
.B(n_751),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_789),
.B(n_737),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_782),
.B(n_768),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_798),
.Y(n_812)
);

AND2x4_ASAP7_75t_SL g813 ( 
.A(n_805),
.B(n_752),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_795),
.B(n_790),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_792),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_804),
.B(n_773),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_792),
.B(n_788),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_793),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_795),
.B(n_790),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_809),
.B(n_791),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_809),
.B(n_791),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_810),
.B(n_786),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_810),
.B(n_786),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_793),
.B(n_788),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_804),
.B(n_773),
.Y(n_825)
);

INVx3_ASAP7_75t_R g826 ( 
.A(n_803),
.Y(n_826)
);

OR2x2_ASAP7_75t_L g827 ( 
.A(n_803),
.B(n_805),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_802),
.B(n_789),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_797),
.B(n_774),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_799),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_797),
.B(n_774),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_829),
.B(n_811),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_815),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_814),
.B(n_800),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_831),
.B(n_811),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_821),
.B(n_811),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_818),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_813),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_830),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_813),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_828),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_819),
.B(n_800),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_817),
.B(n_807),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_817),
.B(n_807),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_827),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_820),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_812),
.Y(n_847)
);

INVxp67_ASAP7_75t_SL g848 ( 
.A(n_847),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_847),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_838),
.A2(n_787),
.B(n_794),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_838),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_841),
.B(n_824),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_833),
.Y(n_853)
);

AO21x1_ASAP7_75t_L g854 ( 
.A1(n_833),
.A2(n_787),
.B(n_837),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_837),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_839),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_839),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_841),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_834),
.B(n_822),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_834),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_845),
.A2(n_779),
.B(n_766),
.C(n_794),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_832),
.Y(n_862)
);

OA222x2_ASAP7_75t_L g863 ( 
.A1(n_840),
.A2(n_826),
.B1(n_804),
.B2(n_778),
.C1(n_773),
.C2(n_785),
.Y(n_863)
);

OAI221xp5_ASAP7_75t_SL g864 ( 
.A1(n_861),
.A2(n_796),
.B1(n_846),
.B2(n_806),
.C(n_840),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_862),
.Y(n_865)
);

OAI31xp33_ASAP7_75t_SL g866 ( 
.A1(n_850),
.A2(n_854),
.A3(n_863),
.B(n_848),
.Y(n_866)
);

OAI221xp5_ASAP7_75t_L g867 ( 
.A1(n_851),
.A2(n_744),
.B1(n_823),
.B2(n_842),
.C(n_824),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_851),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_851),
.A2(n_832),
.B1(n_835),
.B2(n_843),
.Y(n_869)
);

INVxp67_ASAP7_75t_SL g870 ( 
.A(n_854),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_859),
.A2(n_835),
.B1(n_844),
.B2(n_843),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_849),
.B(n_816),
.Y(n_872)
);

AOI221xp5_ASAP7_75t_L g873 ( 
.A1(n_870),
.A2(n_858),
.B1(n_860),
.B2(n_852),
.C(n_855),
.Y(n_873)
);

AOI222xp33_ASAP7_75t_L g874 ( 
.A1(n_870),
.A2(n_860),
.B1(n_858),
.B2(n_855),
.C1(n_856),
.C2(n_862),
.Y(n_874)
);

O2A1O1Ixp5_ASAP7_75t_SL g875 ( 
.A1(n_866),
.A2(n_856),
.B(n_693),
.C(n_715),
.Y(n_875)
);

NAND3xp33_ASAP7_75t_L g876 ( 
.A(n_864),
.B(n_857),
.C(n_853),
.Y(n_876)
);

OAI221xp5_ASAP7_75t_SL g877 ( 
.A1(n_867),
.A2(n_859),
.B1(n_777),
.B2(n_808),
.C(n_844),
.Y(n_877)
);

NAND3xp33_ASAP7_75t_SL g878 ( 
.A(n_868),
.B(n_756),
.C(n_727),
.Y(n_878)
);

OAI32xp33_ASAP7_75t_L g879 ( 
.A1(n_869),
.A2(n_808),
.A3(n_853),
.B1(n_857),
.B2(n_746),
.Y(n_879)
);

AOI221xp5_ASAP7_75t_L g880 ( 
.A1(n_871),
.A2(n_849),
.B1(n_836),
.B2(n_682),
.C(n_649),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_865),
.B(n_836),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_872),
.A2(n_825),
.B1(n_816),
.B2(n_773),
.Y(n_882)
);

AOI21xp33_ASAP7_75t_L g883 ( 
.A1(n_876),
.A2(n_698),
.B(n_682),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_878),
.B(n_765),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_880),
.B(n_873),
.Y(n_885)
);

NAND4xp25_ASAP7_75t_L g886 ( 
.A(n_877),
.B(n_753),
.C(n_734),
.D(n_739),
.Y(n_886)
);

NOR3xp33_ASAP7_75t_L g887 ( 
.A(n_879),
.B(n_702),
.C(n_693),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_882),
.A2(n_825),
.B1(n_816),
.B2(n_765),
.Y(n_888)
);

NOR3xp33_ASAP7_75t_L g889 ( 
.A(n_875),
.B(n_707),
.C(n_695),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_874),
.B(n_799),
.Y(n_890)
);

NOR3xp33_ASAP7_75t_L g891 ( 
.A(n_885),
.B(n_652),
.C(n_695),
.Y(n_891)
);

OAI322xp33_ASAP7_75t_L g892 ( 
.A1(n_890),
.A2(n_881),
.A3(n_754),
.B1(n_740),
.B2(n_747),
.C1(n_743),
.C2(n_741),
.Y(n_892)
);

NAND3xp33_ASAP7_75t_L g893 ( 
.A(n_887),
.B(n_700),
.C(n_697),
.Y(n_893)
);

NOR3x1_ASAP7_75t_L g894 ( 
.A(n_886),
.B(n_888),
.C(n_884),
.Y(n_894)
);

NOR2x1_ASAP7_75t_L g895 ( 
.A(n_883),
.B(n_753),
.Y(n_895)
);

NAND3x1_ASAP7_75t_L g896 ( 
.A(n_889),
.B(n_767),
.C(n_784),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_885),
.B(n_801),
.Y(n_897)
);

NOR2x1_ASAP7_75t_L g898 ( 
.A(n_895),
.B(n_753),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_892),
.B(n_897),
.Y(n_899)
);

NOR2x1_ASAP7_75t_L g900 ( 
.A(n_893),
.B(n_663),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_891),
.A2(n_683),
.B1(n_714),
.B2(n_701),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_894),
.B(n_759),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_896),
.B(n_683),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_893),
.Y(n_904)
);

INVxp67_ASAP7_75t_SL g905 ( 
.A(n_891),
.Y(n_905)
);

NAND4xp75_ASAP7_75t_L g906 ( 
.A(n_902),
.B(n_683),
.C(n_759),
.D(n_699),
.Y(n_906)
);

INVxp33_ASAP7_75t_SL g907 ( 
.A(n_901),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_903),
.B(n_825),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_906),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_907),
.A2(n_905),
.B(n_904),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_908),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_911),
.B(n_899),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_909),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_913),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_912),
.Y(n_915)
);

INVx1_ASAP7_75t_SL g916 ( 
.A(n_913),
.Y(n_916)
);

AOI211xp5_ASAP7_75t_SL g917 ( 
.A1(n_914),
.A2(n_910),
.B(n_713),
.C(n_898),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_916),
.A2(n_900),
.B1(n_701),
.B2(n_687),
.Y(n_918)
);

OAI21x1_ASAP7_75t_SL g919 ( 
.A1(n_915),
.A2(n_691),
.B(n_681),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_917),
.A2(n_716),
.B(n_692),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_920),
.A2(n_919),
.B(n_918),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_921),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_922),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_923),
.A2(n_687),
.B(n_692),
.Y(n_924)
);


endmodule