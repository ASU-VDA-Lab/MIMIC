module fake_jpeg_20406_n_110 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_55),
.Y(n_63)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_53),
.Y(n_69)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_49),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_61),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_56),
.B(n_46),
.Y(n_61)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_51),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_41),
.B1(n_47),
.B2(n_44),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_50),
.B1(n_42),
.B2(n_39),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_79),
.B1(n_7),
.B2(n_8),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_73),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_21),
.C(n_35),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_63),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_20),
.B1(n_34),
.B2(n_33),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_9),
.Y(n_89)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_10),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_91),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_4),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_88),
.B1(n_91),
.B2(n_87),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_89),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_74),
.B1(n_12),
.B2(n_13),
.Y(n_93)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_94),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_95),
.A2(n_85),
.B(n_15),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_99),
.C(n_11),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_22),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_24),
.B(n_25),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_27),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_100),
.C(n_101),
.Y(n_106)
);

NOR2x1_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_28),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_107),
.A2(n_29),
.B(n_31),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_32),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_37),
.Y(n_110)
);


endmodule