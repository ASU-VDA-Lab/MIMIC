module fake_netlist_6_2089_n_1846 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_186, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1846);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_186;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1846;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_268;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g188 ( 
.A(n_15),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_102),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_51),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_42),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_103),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_95),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_164),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_47),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_78),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_48),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_99),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_106),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_177),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_56),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_109),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_18),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_79),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_13),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_119),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_54),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_137),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_83),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_141),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_31),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_59),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_82),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_38),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_133),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_172),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_163),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_84),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_183),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_46),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_86),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_107),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_166),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_26),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_66),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_60),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_169),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_11),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_98),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_74),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_87),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_162),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_29),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_77),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_101),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_158),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_44),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_57),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_152),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_46),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_117),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_65),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_155),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_71),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_142),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_178),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_170),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_62),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_181),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_136),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_116),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_29),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_132),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_58),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_149),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_93),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_23),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_50),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_50),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_64),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_147),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_115),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_88),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_129),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_122),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_33),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_89),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_81),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_43),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_138),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_185),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_134),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_176),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_80),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_30),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_20),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_126),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_30),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_153),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_105),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_173),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_144),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_154),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_146),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_21),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_13),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_53),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_63),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_161),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_121),
.Y(n_294)
);

BUFx8_ASAP7_75t_SL g295 ( 
.A(n_143),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_28),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_17),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_112),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_15),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_125),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_165),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_111),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_150),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_21),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_113),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_97),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_1),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_73),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_40),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_33),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_90),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_5),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_38),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_3),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_42),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_7),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_9),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_20),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_110),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_69),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_174),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_17),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_175),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_36),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_51),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_140),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_53),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_182),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_19),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_49),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_131),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_8),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_19),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_167),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_39),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_171),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_44),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_35),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_76),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_12),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_35),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_151),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_39),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_118),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_91),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_37),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_94),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_68),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_70),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_5),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_145),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_40),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_148),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_23),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_22),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_45),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_157),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_7),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_18),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_12),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_61),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_37),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_27),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_75),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_6),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_135),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_34),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_55),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_36),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_43),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_186),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_124),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_67),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_4),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_261),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_261),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_261),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_208),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_261),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_263),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_216),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_220),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_261),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_292),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_228),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_261),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_261),
.Y(n_387)
);

INVxp33_ASAP7_75t_SL g388 ( 
.A(n_290),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_254),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_261),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_196),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_260),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_359),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_361),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_213),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_274),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_196),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_196),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_196),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_277),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g401 ( 
.A(n_289),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_289),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_309),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_233),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_233),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_309),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_372),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_318),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_295),
.Y(n_409)
);

INVxp33_ASAP7_75t_L g410 ( 
.A(n_188),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_196),
.Y(n_411)
);

BUFx2_ASAP7_75t_SL g412 ( 
.A(n_337),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_318),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_190),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_207),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_289),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_209),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_240),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_279),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_232),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_241),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_279),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g423 ( 
.A(n_316),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_339),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_227),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_229),
.Y(n_426)
);

BUFx6f_ASAP7_75t_SL g427 ( 
.A(n_240),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_237),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_256),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_297),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_299),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_304),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_310),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_291),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_291),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_244),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_268),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_262),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_268),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_273),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_280),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_282),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_296),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_332),
.Y(n_444)
);

INVxp33_ASAP7_75t_SL g445 ( 
.A(n_191),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_234),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_307),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_312),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_315),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_332),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_313),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_314),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_343),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_343),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_317),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_358),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_324),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_363),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_363),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_322),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_235),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_325),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_191),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_330),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_333),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_236),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_287),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_239),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_391),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_375),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_409),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_391),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_404),
.B(n_281),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_397),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_464),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_375),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_399),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_406),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_405),
.B(n_189),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_399),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_418),
.B(n_281),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_397),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_411),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_398),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_411),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_376),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_437),
.B(n_281),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_386),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_386),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_439),
.B(n_189),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_387),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_426),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_446),
.Y(n_494)
);

AND2x6_ASAP7_75t_L g495 ( 
.A(n_387),
.B(n_201),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_388),
.A2(n_338),
.B1(n_270),
.B2(n_198),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_377),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_398),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_390),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_419),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_388),
.A2(n_356),
.B1(n_205),
.B2(n_370),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_468),
.B(n_287),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_378),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_390),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_419),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_395),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_381),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_379),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_434),
.Y(n_509)
);

OA21x2_ASAP7_75t_L g510 ( 
.A1(n_383),
.A2(n_346),
.B(n_335),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_395),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_434),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_435),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_462),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_468),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_435),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_444),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_412),
.B(n_194),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_406),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_444),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_422),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_422),
.Y(n_522)
);

INVx6_ASAP7_75t_L g523 ( 
.A(n_427),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_403),
.B(n_194),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_408),
.B(n_200),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_467),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_412),
.B(n_200),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_413),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_450),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_450),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_453),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_414),
.B(n_192),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_393),
.B(n_316),
.Y(n_533)
);

BUFx8_ASAP7_75t_L g534 ( 
.A(n_427),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_453),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_454),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_454),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_456),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_456),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_457),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_382),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_380),
.A2(n_369),
.B1(n_205),
.B2(n_370),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_415),
.B(n_192),
.Y(n_543)
);

OA21x2_ASAP7_75t_L g544 ( 
.A1(n_457),
.A2(n_355),
.B(n_350),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_417),
.B(n_193),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_459),
.B(n_206),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_393),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_459),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_499),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_489),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_499),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_510),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_474),
.B(n_384),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_477),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_519),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_477),
.Y(n_556)
);

INVxp33_ASAP7_75t_L g557 ( 
.A(n_519),
.Y(n_557)
);

BUFx10_ASAP7_75t_L g558 ( 
.A(n_523),
.Y(n_558)
);

CKINVDCx6p67_ASAP7_75t_R g559 ( 
.A(n_503),
.Y(n_559)
);

AND2x6_ASAP7_75t_L g560 ( 
.A(n_518),
.B(n_206),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_499),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_474),
.B(n_394),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_489),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_477),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_499),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_510),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_478),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_480),
.B(n_445),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_499),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_487),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_487),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_478),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_534),
.B(n_420),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_487),
.Y(n_574)
);

NAND3xp33_ASAP7_75t_L g575 ( 
.A(n_510),
.B(n_428),
.C(n_425),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_SL g576 ( 
.A1(n_496),
.A2(n_423),
.B1(n_401),
.B2(n_424),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_497),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_474),
.B(n_420),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_489),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_534),
.B(n_421),
.Y(n_580)
);

NAND3xp33_ASAP7_75t_L g581 ( 
.A(n_510),
.B(n_438),
.C(n_436),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_478),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_482),
.B(n_421),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_497),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_493),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_489),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_534),
.B(n_429),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_481),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_515),
.B(n_210),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_489),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_481),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_497),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_482),
.B(n_429),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_489),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_481),
.Y(n_595)
);

CKINVDCx11_ASAP7_75t_R g596 ( 
.A(n_507),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_508),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_489),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_484),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_484),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_480),
.B(n_445),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_508),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_508),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_479),
.A2(n_469),
.B1(n_491),
.B2(n_533),
.Y(n_604)
);

OR2x6_ASAP7_75t_L g605 ( 
.A(n_515),
.B(n_210),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_490),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_482),
.B(n_460),
.Y(n_607)
);

INVxp33_ASAP7_75t_L g608 ( 
.A(n_476),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_484),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_510),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_490),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_470),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_534),
.B(n_430),
.Y(n_613)
);

BUFx4f_ASAP7_75t_L g614 ( 
.A(n_544),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_470),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_490),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_534),
.B(n_430),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_502),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_541),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_486),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_473),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_490),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_515),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_479),
.B(n_431),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_488),
.A2(n_337),
.B1(n_368),
.B2(n_367),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_486),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_473),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_475),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_491),
.B(n_431),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_486),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_488),
.A2(n_365),
.B1(n_374),
.B2(n_336),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_475),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_494),
.B(n_385),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_488),
.B(n_432),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_517),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_517),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_502),
.Y(n_637)
);

AOI22x1_ASAP7_75t_L g638 ( 
.A1(n_518),
.A2(n_527),
.B1(n_502),
.B2(n_525),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_490),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_483),
.Y(n_640)
);

CKINVDCx16_ASAP7_75t_R g641 ( 
.A(n_547),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_518),
.B(n_432),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_527),
.A2(n_336),
.B1(n_306),
.B2(n_463),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_483),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_485),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_485),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_527),
.A2(n_306),
.B1(n_465),
.B2(n_461),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_517),
.Y(n_648)
);

AOI21x1_ASAP7_75t_L g649 ( 
.A1(n_498),
.A2(n_212),
.B(n_199),
.Y(n_649)
);

NAND2xp33_ASAP7_75t_L g650 ( 
.A(n_532),
.B(n_543),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_490),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_517),
.Y(n_652)
);

AOI21x1_ASAP7_75t_L g653 ( 
.A1(n_498),
.A2(n_222),
.B(n_214),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_533),
.B(n_433),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_476),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_517),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_490),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_492),
.B(n_433),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_492),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_517),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_492),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_532),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_492),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_517),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_524),
.B(n_460),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_492),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_543),
.B(n_451),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_492),
.B(n_451),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_471),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_492),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_523),
.B(n_231),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_504),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_471),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_L g674 ( 
.A(n_545),
.B(n_452),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_545),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_506),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_504),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_544),
.A2(n_466),
.B1(n_449),
.B2(n_448),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_514),
.Y(n_679)
);

INVxp67_ASAP7_75t_SL g680 ( 
.A(n_504),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_504),
.Y(n_681)
);

INVxp33_ASAP7_75t_L g682 ( 
.A(n_501),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_528),
.B(n_452),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_528),
.B(n_455),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_504),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_547),
.B(n_455),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_504),
.B(n_458),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_471),
.B(n_230),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_524),
.B(n_440),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_471),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_524),
.B(n_301),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_544),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_495),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_R g694 ( 
.A(n_472),
.B(n_389),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_535),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_506),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_L g697 ( 
.A(n_495),
.B(n_201),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_544),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_535),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_662),
.B(n_544),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_662),
.B(n_528),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_675),
.B(n_511),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_568),
.A2(n_407),
.B1(n_400),
.B2(n_396),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_619),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_601),
.B(n_511),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_642),
.B(n_501),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_554),
.Y(n_707)
);

NAND2xp33_ASAP7_75t_L g708 ( 
.A(n_560),
.B(n_242),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_623),
.B(n_521),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_578),
.A2(n_392),
.B1(n_344),
.B2(n_345),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_658),
.A2(n_525),
.B(n_524),
.Y(n_711)
);

BUFx6f_ASAP7_75t_SL g712 ( 
.A(n_589),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_623),
.B(n_521),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_667),
.B(n_526),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_650),
.B(n_521),
.Y(n_715)
);

OR2x6_ASAP7_75t_L g716 ( 
.A(n_696),
.B(n_655),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_554),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_618),
.B(n_521),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_556),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_583),
.B(n_321),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_L g721 ( 
.A(n_560),
.B(n_243),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_614),
.A2(n_524),
.B(n_525),
.C(n_284),
.Y(n_722)
);

NAND2xp33_ASAP7_75t_L g723 ( 
.A(n_560),
.B(n_245),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_618),
.B(n_525),
.Y(n_724)
);

AO221x1_ASAP7_75t_L g725 ( 
.A1(n_604),
.A2(n_496),
.B1(n_542),
.B2(n_302),
.C(n_224),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_637),
.B(n_441),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_637),
.B(n_607),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_607),
.B(n_546),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_556),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_593),
.B(n_402),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_665),
.Y(n_731)
);

INVx4_ASAP7_75t_L g732 ( 
.A(n_563),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_668),
.B(n_546),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_655),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_552),
.A2(n_542),
.B1(n_302),
.B2(n_224),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_634),
.B(n_416),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_555),
.B(n_410),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_687),
.B(n_535),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_553),
.B(n_193),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_564),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_629),
.B(n_427),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_665),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_564),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_552),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_562),
.B(n_195),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_557),
.B(n_195),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_696),
.Y(n_747)
);

NOR2xp67_ASAP7_75t_L g748 ( 
.A(n_575),
.B(n_522),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_589),
.B(n_535),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_566),
.A2(n_201),
.B1(n_224),
.B2(n_302),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_624),
.B(n_197),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_567),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_608),
.B(n_676),
.Y(n_753)
);

HB1xp67_ASAP7_75t_L g754 ( 
.A(n_691),
.Y(n_754)
);

NOR2xp67_ASAP7_75t_L g755 ( 
.A(n_575),
.B(n_522),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_614),
.A2(n_537),
.B(n_530),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_674),
.A2(n_523),
.B1(n_264),
.B2(n_253),
.Y(n_757)
);

O2A1O1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_692),
.A2(n_443),
.B(n_442),
.C(n_447),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_683),
.B(n_197),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_612),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_560),
.B(n_249),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_615),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_615),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_621),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_684),
.B(n_202),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_689),
.B(n_581),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_654),
.B(n_566),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_689),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_621),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_567),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_627),
.B(n_202),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_638),
.B(n_203),
.Y(n_772)
);

NAND3xp33_ASAP7_75t_L g773 ( 
.A(n_625),
.B(n_329),
.C(n_327),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_638),
.B(n_203),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_698),
.A2(n_224),
.B1(n_201),
.B2(n_302),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_647),
.B(n_631),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_690),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_589),
.B(n_535),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_572),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_614),
.A2(n_271),
.B1(n_285),
.B2(n_373),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_698),
.A2(n_201),
.B1(n_224),
.B2(n_302),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_610),
.B(n_535),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_610),
.A2(n_258),
.B1(n_303),
.B2(n_238),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_563),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_643),
.B(n_204),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_627),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_572),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_628),
.B(n_523),
.Y(n_788)
);

AOI221xp5_ASAP7_75t_L g789 ( 
.A1(n_682),
.A2(n_217),
.B1(n_223),
.B2(n_340),
.C(n_341),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_688),
.B(n_204),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_573),
.B(n_211),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_641),
.B(n_316),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_560),
.A2(n_259),
.B1(n_326),
.B2(n_246),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_560),
.A2(n_257),
.B1(n_247),
.B2(n_248),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_632),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_581),
.A2(n_342),
.B1(n_357),
.B2(n_255),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_640),
.B(n_495),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_580),
.B(n_211),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_582),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_644),
.B(n_495),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_644),
.Y(n_801)
);

INVxp67_ASAP7_75t_SL g802 ( 
.A(n_645),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_582),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_587),
.B(n_215),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_645),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_646),
.B(n_495),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_L g807 ( 
.A(n_549),
.B(n_251),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_678),
.A2(n_646),
.B1(n_605),
.B2(n_571),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_613),
.B(n_215),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_549),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_551),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_551),
.B(n_495),
.Y(n_812)
);

AND3x4_ASAP7_75t_L g813 ( 
.A(n_576),
.B(n_540),
.C(n_530),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_686),
.B(n_218),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_561),
.B(n_495),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_561),
.B(n_495),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_605),
.A2(n_266),
.B1(n_252),
.B2(n_265),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_605),
.A2(n_269),
.B1(n_267),
.B2(n_272),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_L g819 ( 
.A(n_565),
.B(n_275),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_563),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_569),
.B(n_520),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_569),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_617),
.B(n_218),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_690),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_690),
.B(n_520),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_680),
.B(n_520),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_659),
.B(n_520),
.Y(n_827)
);

NOR3xp33_ASAP7_75t_L g828 ( 
.A(n_641),
.B(n_250),
.C(n_371),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_605),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_559),
.B(n_585),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_588),
.Y(n_831)
);

OAI22xp33_ASAP7_75t_L g832 ( 
.A1(n_605),
.A2(n_356),
.B1(n_352),
.B2(n_341),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_671),
.B(n_529),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_694),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_588),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_570),
.A2(n_592),
.B1(n_597),
.B2(n_571),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_659),
.B(n_530),
.Y(n_837)
);

AO221x1_ASAP7_75t_L g838 ( 
.A1(n_550),
.A2(n_606),
.B1(n_657),
.B2(n_598),
.C(n_663),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_661),
.B(n_219),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_661),
.A2(n_328),
.B1(n_276),
.B2(n_286),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_591),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_666),
.B(n_537),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_591),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_666),
.B(n_537),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_574),
.Y(n_845)
);

BUFx6f_ASAP7_75t_SL g846 ( 
.A(n_596),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_577),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_681),
.B(n_540),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_681),
.B(n_219),
.Y(n_849)
);

A2O1A1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_577),
.A2(n_548),
.B(n_529),
.C(n_539),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_550),
.B(n_221),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_671),
.A2(n_693),
.B1(n_597),
.B2(n_602),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_550),
.B(n_540),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_594),
.B(n_500),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_671),
.A2(n_334),
.B1(n_221),
.B2(n_225),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_585),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_693),
.B(n_225),
.Y(n_857)
);

OR2x6_ASAP7_75t_L g858 ( 
.A(n_559),
.B(n_531),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_720),
.B(n_679),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_810),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_744),
.B(n_584),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_811),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_753),
.B(n_679),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_SL g864 ( 
.A1(n_706),
.A2(n_360),
.B1(n_223),
.B2(n_217),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_750),
.A2(n_340),
.B1(n_354),
.B2(n_360),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_766),
.A2(n_602),
.B1(n_592),
.B2(n_603),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_702),
.B(n_579),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_777),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_736),
.B(n_531),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_744),
.B(n_603),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_802),
.B(n_594),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_768),
.B(n_671),
.Y(n_872)
);

BUFx12f_ASAP7_75t_L g873 ( 
.A(n_858),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_737),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_822),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_736),
.B(n_536),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_802),
.B(n_594),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_760),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_731),
.B(n_671),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_706),
.A2(n_606),
.B(n_598),
.C(n_611),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_727),
.A2(n_697),
.B(n_669),
.C(n_673),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_742),
.B(n_536),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_784),
.Y(n_883)
);

AO22x1_ASAP7_75t_L g884 ( 
.A1(n_813),
.A2(n_352),
.B1(n_354),
.B2(n_362),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_766),
.B(n_598),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_733),
.B(n_606),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_704),
.Y(n_887)
);

BUFx4f_ASAP7_75t_L g888 ( 
.A(n_716),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_738),
.A2(n_590),
.B(n_579),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_700),
.B(n_611),
.Y(n_890)
);

BUFx12f_ASAP7_75t_L g891 ( 
.A(n_858),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_716),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_726),
.B(n_538),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_720),
.B(n_611),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_762),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_716),
.Y(n_896)
);

NOR2xp67_ASAP7_75t_L g897 ( 
.A(n_834),
.B(n_695),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_777),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_763),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_750),
.A2(n_362),
.B1(n_538),
.B2(n_539),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_754),
.B(n_657),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_702),
.B(n_558),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_754),
.B(n_657),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_728),
.B(n_663),
.Y(n_904)
);

INVx5_ASAP7_75t_L g905 ( 
.A(n_784),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_764),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_769),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_707),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_767),
.B(n_663),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_786),
.Y(n_910)
);

INVxp67_ASAP7_75t_SL g911 ( 
.A(n_784),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_759),
.B(n_558),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_759),
.B(n_670),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_726),
.B(n_548),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_725),
.A2(n_669),
.B1(n_673),
.B2(n_699),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_730),
.B(n_558),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_717),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_746),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_719),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_767),
.B(n_775),
.Y(n_920)
);

BUFx8_ASAP7_75t_L g921 ( 
.A(n_846),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_792),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_795),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_735),
.A2(n_783),
.B1(n_776),
.B2(n_780),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_846),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_801),
.Y(n_926)
);

CKINVDCx16_ASAP7_75t_R g927 ( 
.A(n_703),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_856),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_805),
.Y(n_929)
);

NOR3xp33_ASAP7_75t_SL g930 ( 
.A(n_710),
.B(n_226),
.C(n_278),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_701),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_734),
.B(n_500),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_775),
.B(n_670),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_781),
.B(n_672),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_729),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_740),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_783),
.B(n_672),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_830),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_743),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_747),
.Y(n_940)
);

INVxp67_ASAP7_75t_SL g941 ( 
.A(n_784),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_734),
.B(n_505),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_781),
.B(n_672),
.Y(n_943)
);

O2A1O1Ixp5_ASAP7_75t_L g944 ( 
.A1(n_772),
.A2(n_649),
.B(n_653),
.C(n_636),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_748),
.B(n_635),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_752),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_755),
.B(n_635),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_845),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_714),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_747),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_735),
.B(n_718),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_770),
.Y(n_952)
);

AOI221xp5_ASAP7_75t_SL g953 ( 
.A1(n_758),
.A2(n_516),
.B1(n_513),
.B2(n_512),
.C(n_509),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_796),
.A2(n_699),
.B1(n_695),
.B2(n_636),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_808),
.B(n_724),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_833),
.B(n_648),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_847),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_705),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_779),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_813),
.Y(n_960)
);

AND2x6_ASAP7_75t_SL g961 ( 
.A(n_814),
.B(n_505),
.Y(n_961)
);

OR2x2_ASAP7_75t_SL g962 ( 
.A(n_773),
.B(n_509),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_751),
.A2(n_648),
.B(n_652),
.C(n_664),
.Y(n_963)
);

NOR3xp33_ASAP7_75t_SL g964 ( 
.A(n_789),
.B(n_283),
.C(n_278),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_787),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_808),
.B(n_652),
.Y(n_966)
);

INVx5_ASAP7_75t_L g967 ( 
.A(n_820),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_751),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_771),
.B(n_563),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_765),
.B(n_586),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_829),
.B(n_656),
.Y(n_971)
);

INVx4_ASAP7_75t_L g972 ( 
.A(n_712),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_829),
.A2(n_626),
.B(n_609),
.C(n_620),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_824),
.Y(n_974)
);

AND2x6_ASAP7_75t_L g975 ( 
.A(n_852),
.B(n_656),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_R g976 ( 
.A(n_712),
.B(n_226),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_771),
.B(n_563),
.Y(n_977)
);

NAND2xp33_ASAP7_75t_L g978 ( 
.A(n_796),
.B(n_616),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_782),
.B(n_660),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_709),
.B(n_713),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_832),
.B(n_283),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_790),
.Y(n_982)
);

NOR3xp33_ASAP7_75t_L g983 ( 
.A(n_791),
.B(n_353),
.C(n_331),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_756),
.A2(n_664),
.B(n_660),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_799),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_836),
.B(n_595),
.Y(n_986)
);

AND2x2_ASAP7_75t_SL g987 ( 
.A(n_828),
.B(n_586),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_741),
.Y(n_988)
);

NAND2x1p5_ASAP7_75t_L g989 ( 
.A(n_732),
.B(n_586),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_739),
.A2(n_685),
.B1(n_677),
.B2(n_590),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_820),
.Y(n_991)
);

AND2x6_ASAP7_75t_SL g992 ( 
.A(n_839),
.B(n_512),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_854),
.Y(n_993)
);

BUFx8_ASAP7_75t_L g994 ( 
.A(n_803),
.Y(n_994)
);

NAND2x1p5_ASAP7_75t_L g995 ( 
.A(n_732),
.B(n_590),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_820),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_745),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_836),
.B(n_595),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_793),
.A2(n_630),
.B1(n_620),
.B2(n_599),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_715),
.B(n_599),
.Y(n_1000)
);

INVx5_ASAP7_75t_L g1001 ( 
.A(n_820),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_839),
.B(n_616),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_831),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_835),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_798),
.B(n_804),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_809),
.B(n_677),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_828),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_823),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_849),
.B(n_616),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_832),
.B(n_677),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_817),
.B(n_331),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_711),
.B(n_600),
.Y(n_1012)
);

NOR3xp33_ASAP7_75t_SL g1013 ( 
.A(n_855),
.B(n_366),
.C(n_364),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_841),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_843),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_757),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_838),
.B(n_600),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_821),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_807),
.A2(n_685),
.B1(n_616),
.B2(n_651),
.Y(n_1019)
);

INVx5_ASAP7_75t_L g1020 ( 
.A(n_722),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_840),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_850),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_749),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_837),
.B(n_609),
.Y(n_1024)
);

OR2x6_ASAP7_75t_L g1025 ( 
.A(n_785),
.B(n_685),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_778),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_825),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_819),
.A2(n_849),
.B1(n_851),
.B2(n_708),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_818),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_812),
.A2(n_653),
.B(n_649),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_797),
.B(n_800),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_806),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_842),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_844),
.Y(n_1034)
);

INVxp67_ASAP7_75t_L g1035 ( 
.A(n_827),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_848),
.B(n_793),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_794),
.B(n_626),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_794),
.B(n_630),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_853),
.B(n_826),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_815),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_883),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_968),
.B(n_857),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_887),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_918),
.B(n_859),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_984),
.A2(n_774),
.B(n_816),
.Y(n_1045)
);

CKINVDCx11_ASAP7_75t_R g1046 ( 
.A(n_873),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_860),
.Y(n_1047)
);

INVx3_ASAP7_75t_SL g1048 ( 
.A(n_925),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_878),
.Y(n_1049)
);

NAND2x1p5_ASAP7_75t_L g1050 ( 
.A(n_928),
.B(n_616),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_994),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_908),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_863),
.B(n_513),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_920),
.A2(n_788),
.B(n_761),
.C(n_723),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_869),
.B(n_721),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_876),
.B(n_516),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_994),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_874),
.B(n_334),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_920),
.A2(n_347),
.B(n_348),
.C(n_349),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_960),
.A2(n_347),
.B1(n_349),
.B2(n_351),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_931),
.B(n_622),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_981),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_1010),
.A2(n_351),
.B1(n_353),
.B2(n_364),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_955),
.A2(n_366),
.B1(n_639),
.B2(n_622),
.Y(n_1064)
);

O2A1O1Ixp5_ASAP7_75t_L g1065 ( 
.A1(n_912),
.A2(n_916),
.B(n_867),
.C(n_902),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_949),
.B(n_319),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_940),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_950),
.B(n_311),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_905),
.A2(n_651),
.B(n_639),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_951),
.A2(n_651),
.B1(n_639),
.B2(n_622),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_921),
.Y(n_1071)
);

INVx4_ASAP7_75t_L g1072 ( 
.A(n_905),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_893),
.B(n_639),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1033),
.B(n_323),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_1007),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_1075)
);

NAND3xp33_ASAP7_75t_L g1076 ( 
.A(n_930),
.B(n_964),
.C(n_864),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_955),
.A2(n_320),
.B1(n_308),
.B2(n_305),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_1016),
.A2(n_300),
.B1(n_298),
.B2(n_294),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_893),
.B(n_123),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1034),
.B(n_293),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1035),
.B(n_288),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_895),
.B(n_4),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_899),
.B(n_6),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_951),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_1084)
);

AO21x1_ASAP7_75t_L g1085 ( 
.A1(n_1028),
.A2(n_10),
.B(n_11),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_967),
.A2(n_187),
.B(n_180),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_967),
.A2(n_179),
.B(n_160),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_883),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_958),
.B(n_14),
.Y(n_1089)
);

NAND2x1p5_ASAP7_75t_L g1090 ( 
.A(n_972),
.B(n_159),
.Y(n_1090)
);

BUFx8_ASAP7_75t_L g1091 ( 
.A(n_891),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_906),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_896),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_967),
.A2(n_156),
.B(n_130),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_907),
.B(n_14),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_910),
.B(n_16),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1001),
.A2(n_128),
.B(n_120),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_917),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_923),
.B(n_16),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_919),
.Y(n_1100)
);

O2A1O1Ixp5_ASAP7_75t_L g1101 ( 
.A1(n_970),
.A2(n_114),
.B(n_108),
.C(n_104),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_935),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_988),
.B(n_22),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_936),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_1021),
.B(n_100),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_888),
.Y(n_1106)
);

BUFx8_ASAP7_75t_L g1107 ( 
.A(n_892),
.Y(n_1107)
);

OR2x6_ASAP7_75t_L g1108 ( 
.A(n_972),
.B(n_938),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_927),
.B(n_24),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_969),
.A2(n_96),
.B1(n_92),
.B2(n_85),
.Y(n_1110)
);

NAND2x1p5_ASAP7_75t_L g1111 ( 
.A(n_1001),
.B(n_72),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_926),
.B(n_24),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_922),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_880),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_929),
.B(n_25),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_914),
.B(n_997),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1005),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_939),
.Y(n_1118)
);

AND2x6_ASAP7_75t_L g1119 ( 
.A(n_1032),
.B(n_879),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_921),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_978),
.A2(n_32),
.B1(n_34),
.B2(n_41),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1008),
.A2(n_41),
.B(n_45),
.C(n_47),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_914),
.B(n_48),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_1001),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_993),
.B(n_49),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_1001),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1012),
.A2(n_52),
.B(n_54),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_888),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1012),
.A2(n_52),
.B(n_55),
.Y(n_1129)
);

CKINVDCx20_ASAP7_75t_R g1130 ( 
.A(n_1029),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_948),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_946),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_883),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_966),
.A2(n_866),
.B1(n_998),
.B2(n_986),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1023),
.B(n_957),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_886),
.A2(n_1009),
.B(n_1002),
.Y(n_1136)
);

INVx4_ASAP7_75t_L g1137 ( 
.A(n_991),
.Y(n_1137)
);

BUFx10_ASAP7_75t_L g1138 ( 
.A(n_961),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_886),
.A2(n_1039),
.B(n_890),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_991),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1011),
.A2(n_865),
.B(n_983),
.C(n_982),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1039),
.A2(n_890),
.B(n_989),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_992),
.B(n_1005),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_R g1144 ( 
.A(n_987),
.B(n_868),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_991),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_962),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_932),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_956),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_989),
.A2(n_995),
.B(n_909),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_952),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_884),
.B(n_942),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1022),
.A2(n_1006),
.B(n_1027),
.C(n_875),
.Y(n_1152)
);

INVx3_ASAP7_75t_SL g1153 ( 
.A(n_882),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_862),
.A2(n_1018),
.B(n_894),
.C(n_1036),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_882),
.B(n_956),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_959),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1036),
.A2(n_1040),
.B(n_913),
.C(n_1026),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1003),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_966),
.A2(n_998),
.B1(n_986),
.B2(n_943),
.Y(n_1159)
);

BUFx8_ASAP7_75t_L g1160 ( 
.A(n_872),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_872),
.B(n_879),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1004),
.Y(n_1162)
);

NOR3xp33_ASAP7_75t_L g1163 ( 
.A(n_865),
.B(n_885),
.C(n_901),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_903),
.B(n_1032),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_868),
.B(n_1013),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_904),
.B(n_1026),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_904),
.A2(n_885),
.B(n_937),
.C(n_977),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_980),
.B(n_871),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_881),
.A2(n_974),
.B(n_1031),
.C(n_980),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_976),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_971),
.Y(n_1171)
);

AOI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1017),
.A2(n_909),
.B(n_979),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_933),
.A2(n_943),
.B1(n_934),
.B2(n_871),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1015),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_971),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_933),
.A2(n_934),
.B1(n_877),
.B2(n_1020),
.Y(n_1176)
);

CKINVDCx11_ASAP7_75t_R g1177 ( 
.A(n_1025),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1031),
.A2(n_973),
.B(n_1037),
.C(n_1038),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_877),
.B(n_979),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_900),
.A2(n_1017),
.B(n_963),
.C(n_945),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1032),
.B(n_898),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1014),
.B(n_985),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_944),
.A2(n_1030),
.B(n_984),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_861),
.B(n_870),
.Y(n_1184)
);

INVx5_ASAP7_75t_L g1185 ( 
.A(n_996),
.Y(n_1185)
);

NOR2x1_ASAP7_75t_L g1186 ( 
.A(n_897),
.B(n_996),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_889),
.A2(n_1030),
.B(n_870),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1037),
.A2(n_1038),
.B(n_947),
.C(n_945),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_947),
.A2(n_965),
.B(n_915),
.C(n_1020),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1014),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_911),
.B(n_941),
.Y(n_1191)
);

INVx4_ASAP7_75t_L g1192 ( 
.A(n_975),
.Y(n_1192)
);

OA21x2_ASAP7_75t_L g1193 ( 
.A1(n_1183),
.A2(n_953),
.B(n_1000),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1049),
.Y(n_1194)
);

INVx2_ASAP7_75t_SL g1195 ( 
.A(n_1067),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1187),
.A2(n_1024),
.B(n_995),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1147),
.B(n_975),
.Y(n_1197)
);

INVxp67_ASAP7_75t_SL g1198 ( 
.A(n_1168),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1139),
.A2(n_954),
.B(n_975),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1147),
.B(n_900),
.Y(n_1200)
);

AOI221x1_ASAP7_75t_L g1201 ( 
.A1(n_1084),
.A2(n_1127),
.B1(n_1129),
.B2(n_1176),
.C(n_1189),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1136),
.A2(n_1020),
.B(n_1019),
.Y(n_1202)
);

NAND2xp33_ASAP7_75t_R g1203 ( 
.A(n_1043),
.B(n_1025),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1045),
.A2(n_999),
.B(n_990),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1056),
.B(n_975),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1092),
.Y(n_1206)
);

AO31x2_ASAP7_75t_L g1207 ( 
.A1(n_1176),
.A2(n_1020),
.A3(n_1025),
.B(n_1152),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1142),
.A2(n_1054),
.B(n_1179),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1053),
.B(n_1151),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1044),
.B(n_1042),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_1093),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_SL g1212 ( 
.A1(n_1055),
.A2(n_1178),
.B(n_1169),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1143),
.A2(n_1146),
.B1(n_1076),
.B2(n_1121),
.Y(n_1213)
);

AND2x2_ASAP7_75t_SL g1214 ( 
.A(n_1121),
.B(n_1192),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1135),
.B(n_1164),
.Y(n_1215)
);

AOI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1172),
.A2(n_1070),
.B(n_1173),
.Y(n_1216)
);

AOI221xp5_ASAP7_75t_L g1217 ( 
.A1(n_1076),
.A2(n_1109),
.B1(n_1084),
.B2(n_1141),
.C(n_1103),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1183),
.A2(n_1184),
.B(n_1188),
.Y(n_1218)
);

NOR2xp67_ASAP7_75t_SL g1219 ( 
.A(n_1051),
.B(n_1057),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1171),
.B(n_1155),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1167),
.A2(n_1157),
.B(n_1180),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1070),
.A2(n_1069),
.B(n_1173),
.Y(n_1222)
);

BUFx4_ASAP7_75t_SL g1223 ( 
.A(n_1120),
.Y(n_1223)
);

NAND3xp33_ASAP7_75t_L g1224 ( 
.A(n_1063),
.B(n_1117),
.C(n_1077),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1072),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1154),
.A2(n_1065),
.B(n_1163),
.C(n_1062),
.Y(n_1226)
);

AOI21xp33_ASAP7_75t_L g1227 ( 
.A1(n_1114),
.A2(n_1077),
.B(n_1134),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1155),
.B(n_1161),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1166),
.A2(n_1159),
.B(n_1134),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1131),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1072),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1159),
.A2(n_1186),
.B(n_1101),
.Y(n_1232)
);

NAND2x1_ASAP7_75t_L g1233 ( 
.A(n_1124),
.B(n_1126),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1153),
.B(n_1175),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1192),
.A2(n_1125),
.B1(n_1171),
.B2(n_1079),
.Y(n_1235)
);

AO21x1_ASAP7_75t_L g1236 ( 
.A1(n_1110),
.A2(n_1165),
.B(n_1075),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1074),
.B(n_1081),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1061),
.A2(n_1064),
.B(n_1087),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1068),
.B(n_1060),
.Y(n_1239)
);

INVx8_ASAP7_75t_L g1240 ( 
.A(n_1119),
.Y(n_1240)
);

AOI221xp5_ASAP7_75t_L g1241 ( 
.A1(n_1089),
.A2(n_1123),
.B1(n_1122),
.B2(n_1085),
.C(n_1059),
.Y(n_1241)
);

OR2x6_ASAP7_75t_L g1242 ( 
.A(n_1108),
.B(n_1106),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1082),
.A2(n_1083),
.B(n_1099),
.Y(n_1243)
);

AO22x2_ASAP7_75t_L g1244 ( 
.A1(n_1095),
.A2(n_1096),
.B1(n_1112),
.B2(n_1115),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1047),
.B(n_1080),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1119),
.B(n_1182),
.Y(n_1246)
);

INVxp67_ASAP7_75t_SL g1247 ( 
.A(n_1148),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1181),
.A2(n_1158),
.B(n_1162),
.C(n_1174),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1052),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1119),
.B(n_1073),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1086),
.A2(n_1097),
.B(n_1094),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1107),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1050),
.A2(n_1111),
.B(n_1100),
.Y(n_1253)
);

INVx4_ASAP7_75t_L g1254 ( 
.A(n_1124),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1098),
.A2(n_1150),
.B(n_1118),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1126),
.A2(n_1191),
.B(n_1190),
.Y(n_1256)
);

A2O1A1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1102),
.A2(n_1104),
.B(n_1156),
.C(n_1132),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1116),
.Y(n_1258)
);

AND2x6_ASAP7_75t_SL g1259 ( 
.A(n_1108),
.B(n_1073),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1088),
.A2(n_1090),
.B(n_1105),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1119),
.B(n_1148),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1066),
.B(n_1078),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1058),
.A2(n_1185),
.B(n_1108),
.Y(n_1263)
);

NAND3xp33_ASAP7_75t_L g1264 ( 
.A(n_1177),
.B(n_1160),
.C(n_1107),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1144),
.A2(n_1137),
.B(n_1041),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1128),
.A2(n_1130),
.B1(n_1041),
.B2(n_1133),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1041),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1160),
.A2(n_1138),
.B1(n_1113),
.B2(n_1170),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1138),
.B(n_1145),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1133),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1140),
.B(n_1145),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1140),
.B(n_1145),
.Y(n_1272)
);

OA21x2_ASAP7_75t_L g1273 ( 
.A1(n_1071),
.A2(n_1091),
.B(n_1046),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1048),
.B(n_1091),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1147),
.B(n_927),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1136),
.A2(n_1142),
.B(n_1139),
.Y(n_1276)
);

NAND3x1_ASAP7_75t_L g1277 ( 
.A(n_1109),
.B(n_703),
.C(n_706),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1168),
.A2(n_924),
.B1(n_750),
.B2(n_781),
.Y(n_1278)
);

INVx4_ASAP7_75t_L g1279 ( 
.A(n_1072),
.Y(n_1279)
);

INVx4_ASAP7_75t_L g1280 ( 
.A(n_1072),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1147),
.B(n_1053),
.Y(n_1281)
);

AOI21x1_ASAP7_75t_SL g1282 ( 
.A1(n_1055),
.A2(n_1125),
.B(n_1005),
.Y(n_1282)
);

OA21x2_ASAP7_75t_L g1283 ( 
.A1(n_1183),
.A2(n_1189),
.B(n_1187),
.Y(n_1283)
);

AOI21xp33_ASAP7_75t_L g1284 ( 
.A1(n_1141),
.A2(n_706),
.B(n_759),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1093),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1147),
.B(n_869),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1147),
.B(n_1053),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1049),
.Y(n_1288)
);

NAND3xp33_ASAP7_75t_L g1289 ( 
.A(n_1076),
.B(n_759),
.C(n_968),
.Y(n_1289)
);

NAND3xp33_ASAP7_75t_L g1290 ( 
.A(n_1076),
.B(n_759),
.C(n_968),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1041),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1136),
.A2(n_1142),
.B(n_1139),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1067),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1072),
.Y(n_1294)
);

AOI21xp33_ASAP7_75t_L g1295 ( 
.A1(n_1141),
.A2(n_759),
.B(n_720),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1049),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1147),
.B(n_869),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1049),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1136),
.A2(n_1142),
.B(n_1139),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1049),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1136),
.A2(n_1142),
.B(n_1139),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1093),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1139),
.A2(n_1167),
.B(n_1157),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1067),
.Y(n_1304)
);

NAND2x1p5_ASAP7_75t_L g1305 ( 
.A(n_1072),
.B(n_1124),
.Y(n_1305)
);

BUFx8_ASAP7_75t_L g1306 ( 
.A(n_1120),
.Y(n_1306)
);

CKINVDCx14_ASAP7_75t_R g1307 ( 
.A(n_1071),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1147),
.B(n_1053),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1176),
.A2(n_1189),
.A3(n_1152),
.B(n_1173),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1147),
.B(n_869),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1147),
.B(n_927),
.Y(n_1311)
);

INVx6_ASAP7_75t_SL g1312 ( 
.A(n_1108),
.Y(n_1312)
);

OAI22x1_ASAP7_75t_L g1313 ( 
.A1(n_1121),
.A2(n_813),
.B1(n_1146),
.B2(n_1076),
.Y(n_1313)
);

NAND2x1_ASAP7_75t_L g1314 ( 
.A(n_1072),
.B(n_1124),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1147),
.B(n_869),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1136),
.A2(n_1142),
.B(n_1139),
.Y(n_1316)
);

BUFx8_ASAP7_75t_SL g1317 ( 
.A(n_1071),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1139),
.A2(n_1167),
.B(n_1157),
.Y(n_1318)
);

CKINVDCx11_ASAP7_75t_R g1319 ( 
.A(n_1048),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1168),
.A2(n_924),
.B1(n_750),
.B2(n_781),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1139),
.A2(n_1167),
.B(n_1157),
.Y(n_1321)
);

AO22x2_ASAP7_75t_L g1322 ( 
.A1(n_1084),
.A2(n_813),
.B1(n_1076),
.B2(n_1176),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1136),
.A2(n_1142),
.B(n_1139),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1147),
.B(n_869),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1147),
.B(n_869),
.Y(n_1325)
);

NOR2xp67_ASAP7_75t_L g1326 ( 
.A(n_1043),
.B(n_856),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1147),
.B(n_869),
.Y(n_1327)
);

AOI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1149),
.A2(n_1172),
.B(n_1142),
.Y(n_1328)
);

CKINVDCx11_ASAP7_75t_R g1329 ( 
.A(n_1048),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1147),
.B(n_869),
.Y(n_1330)
);

BUFx10_ASAP7_75t_L g1331 ( 
.A(n_1143),
.Y(n_1331)
);

AOI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1149),
.A2(n_1172),
.B(n_1142),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1147),
.B(n_869),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_SL g1334 ( 
.A1(n_1085),
.A2(n_1114),
.B(n_1121),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1141),
.A2(n_705),
.B(n_968),
.C(n_859),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1147),
.B(n_869),
.Y(n_1336)
);

A2O1A1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1141),
.A2(n_706),
.B(n_924),
.C(n_968),
.Y(n_1337)
);

AOI31xp67_ASAP7_75t_L g1338 ( 
.A1(n_1055),
.A2(n_1028),
.A3(n_774),
.B(n_772),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1136),
.A2(n_1142),
.B(n_1139),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1295),
.A2(n_1284),
.B(n_1337),
.Y(n_1340)
);

NAND2x1p5_ASAP7_75t_L g1341 ( 
.A(n_1260),
.B(n_1265),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1210),
.B(n_1198),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1277),
.A2(n_1217),
.B1(n_1289),
.B2(n_1290),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_SL g1344 ( 
.A(n_1317),
.B(n_1326),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1281),
.B(n_1287),
.Y(n_1345)
);

AO31x2_ASAP7_75t_L g1346 ( 
.A1(n_1201),
.A2(n_1339),
.A3(n_1323),
.B(n_1276),
.Y(n_1346)
);

AO21x2_ASAP7_75t_L g1347 ( 
.A1(n_1295),
.A2(n_1299),
.B(n_1292),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1335),
.B(n_1289),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1207),
.Y(n_1349)
);

CKINVDCx6p67_ASAP7_75t_R g1350 ( 
.A(n_1319),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1206),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1290),
.B(n_1275),
.Y(n_1352)
);

NOR2xp67_ASAP7_75t_L g1353 ( 
.A(n_1195),
.B(n_1211),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1308),
.B(n_1215),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1240),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1230),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1311),
.Y(n_1357)
);

AO32x2_ASAP7_75t_L g1358 ( 
.A1(n_1235),
.A2(n_1278),
.A3(n_1320),
.B1(n_1266),
.B2(n_1322),
.Y(n_1358)
);

AOI22x1_ASAP7_75t_L g1359 ( 
.A1(n_1244),
.A2(n_1322),
.B1(n_1313),
.B2(n_1334),
.Y(n_1359)
);

CKINVDCx6p67_ASAP7_75t_R g1360 ( 
.A(n_1329),
.Y(n_1360)
);

OA21x2_ASAP7_75t_L g1361 ( 
.A1(n_1303),
.A2(n_1321),
.B(n_1318),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1223),
.Y(n_1362)
);

OA21x2_ASAP7_75t_L g1363 ( 
.A1(n_1303),
.A2(n_1321),
.B(n_1318),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1224),
.A2(n_1239),
.B1(n_1227),
.B2(n_1241),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1194),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1224),
.A2(n_1227),
.B1(n_1214),
.B2(n_1244),
.Y(n_1366)
);

AO21x2_ASAP7_75t_L g1367 ( 
.A1(n_1301),
.A2(n_1316),
.B(n_1208),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1293),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_R g1369 ( 
.A(n_1213),
.B(n_1252),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1286),
.B(n_1297),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1204),
.A2(n_1202),
.B(n_1222),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1243),
.A2(n_1237),
.B(n_1226),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1251),
.A2(n_1282),
.B(n_1238),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1213),
.B(n_1209),
.Y(n_1374)
);

AOI221xp5_ASAP7_75t_L g1375 ( 
.A1(n_1278),
.A2(n_1320),
.B1(n_1324),
.B2(n_1315),
.C(n_1310),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1288),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1325),
.B(n_1327),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1240),
.Y(n_1378)
);

AOI221xp5_ASAP7_75t_L g1379 ( 
.A1(n_1330),
.A2(n_1333),
.B1(n_1336),
.B2(n_1243),
.C(n_1221),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_SL g1380 ( 
.A1(n_1199),
.A2(n_1248),
.B(n_1205),
.C(n_1251),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1212),
.A2(n_1218),
.B(n_1199),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1296),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1307),
.Y(n_1383)
);

A2O1A1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1221),
.A2(n_1262),
.B(n_1229),
.C(n_1245),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1298),
.Y(n_1385)
);

OR2x6_ASAP7_75t_L g1386 ( 
.A(n_1240),
.B(n_1263),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1235),
.A2(n_1232),
.B(n_1246),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1216),
.A2(n_1253),
.B(n_1283),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1304),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1283),
.A2(n_1193),
.B(n_1256),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1200),
.B(n_1220),
.Y(n_1391)
);

OR2x6_ASAP7_75t_L g1392 ( 
.A(n_1263),
.B(n_1242),
.Y(n_1392)
);

AO21x2_ASAP7_75t_L g1393 ( 
.A1(n_1236),
.A2(n_1197),
.B(n_1255),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1300),
.Y(n_1394)
);

AO31x2_ASAP7_75t_L g1395 ( 
.A1(n_1338),
.A2(n_1257),
.A3(n_1207),
.B(n_1309),
.Y(n_1395)
);

BUFx12f_ASAP7_75t_L g1396 ( 
.A(n_1306),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1258),
.B(n_1228),
.Y(n_1397)
);

AO31x2_ASAP7_75t_L g1398 ( 
.A1(n_1207),
.A2(n_1309),
.A3(n_1193),
.B(n_1249),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1255),
.A2(n_1314),
.B(n_1233),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1234),
.B(n_1302),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1305),
.A2(n_1294),
.B(n_1225),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1267),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1331),
.A2(n_1264),
.B1(n_1273),
.B2(n_1242),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1285),
.B(n_1247),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1312),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1270),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1254),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1231),
.A2(n_1294),
.B(n_1250),
.Y(n_1408)
);

INVx8_ASAP7_75t_L g1409 ( 
.A(n_1291),
.Y(n_1409)
);

AO21x2_ASAP7_75t_L g1410 ( 
.A1(n_1261),
.A2(n_1271),
.B(n_1272),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1331),
.Y(n_1411)
);

AO31x2_ASAP7_75t_L g1412 ( 
.A1(n_1279),
.A2(n_1280),
.A3(n_1259),
.B(n_1203),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1268),
.B(n_1269),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1291),
.Y(n_1414)
);

AOI22x1_ASAP7_75t_L g1415 ( 
.A1(n_1279),
.A2(n_1259),
.B1(n_1312),
.B2(n_1274),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1264),
.A2(n_1219),
.B(n_1273),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1284),
.A2(n_1337),
.B(n_1295),
.C(n_1217),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1240),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1196),
.A2(n_1332),
.B(n_1328),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1284),
.A2(n_1217),
.B1(n_725),
.B2(n_1224),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1210),
.A2(n_1277),
.B1(n_1198),
.B2(n_924),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_1317),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1319),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1196),
.A2(n_1332),
.B(n_1328),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1206),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1209),
.B(n_1281),
.Y(n_1426)
);

AO21x2_ASAP7_75t_L g1427 ( 
.A1(n_1295),
.A2(n_1292),
.B(n_1276),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1293),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1206),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1210),
.B(n_1284),
.Y(n_1430)
);

AO31x2_ASAP7_75t_L g1431 ( 
.A1(n_1201),
.A2(n_1276),
.A3(n_1299),
.B(n_1292),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1210),
.B(n_1284),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_SL g1433 ( 
.A(n_1317),
.B(n_585),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1206),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1277),
.A2(n_633),
.B1(n_1239),
.B2(n_1210),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1209),
.B(n_1281),
.Y(n_1436)
);

CKINVDCx20_ASAP7_75t_R g1437 ( 
.A(n_1317),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_SL g1438 ( 
.A1(n_1236),
.A2(n_1085),
.B(n_1334),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1277),
.A2(n_633),
.B1(n_1239),
.B2(n_1210),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1240),
.Y(n_1440)
);

NAND3x1_ASAP7_75t_L g1441 ( 
.A(n_1210),
.B(n_1109),
.C(n_1268),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1210),
.A2(n_1277),
.B1(n_1198),
.B2(n_924),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1201),
.A2(n_1318),
.B(n_1303),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_SL g1444 ( 
.A1(n_1236),
.A2(n_1085),
.B(n_1334),
.Y(n_1444)
);

OR2x6_ASAP7_75t_L g1445 ( 
.A(n_1240),
.B(n_1192),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1196),
.A2(n_1332),
.B(n_1328),
.Y(n_1446)
);

AO31x2_ASAP7_75t_L g1447 ( 
.A1(n_1201),
.A2(n_1276),
.A3(n_1299),
.B(n_1292),
.Y(n_1447)
);

O2A1O1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1284),
.A2(n_1337),
.B(n_1295),
.C(n_1217),
.Y(n_1448)
);

OA21x2_ASAP7_75t_L g1449 ( 
.A1(n_1201),
.A2(n_1318),
.B(n_1303),
.Y(n_1449)
);

OA21x2_ASAP7_75t_L g1450 ( 
.A1(n_1201),
.A2(n_1318),
.B(n_1303),
.Y(n_1450)
);

AOI221xp5_ASAP7_75t_L g1451 ( 
.A1(n_1284),
.A2(n_1217),
.B1(n_706),
.B2(n_1295),
.C(n_1210),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1196),
.A2(n_1332),
.B(n_1328),
.Y(n_1452)
);

INVx1_ASAP7_75t_SL g1453 ( 
.A(n_1275),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_SL g1454 ( 
.A(n_1284),
.B(n_1217),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1284),
.A2(n_1337),
.B(n_1295),
.C(n_1217),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1284),
.A2(n_1217),
.B1(n_725),
.B2(n_1224),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1304),
.Y(n_1457)
);

NOR2xp67_ASAP7_75t_L g1458 ( 
.A(n_1326),
.B(n_856),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1209),
.B(n_1281),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1295),
.A2(n_1292),
.B(n_1276),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1196),
.A2(n_1332),
.B(n_1328),
.Y(n_1461)
);

AOI222xp33_ASAP7_75t_L g1462 ( 
.A1(n_1217),
.A2(n_496),
.B1(n_706),
.B2(n_1224),
.C1(n_1239),
.C2(n_1210),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1201),
.A2(n_1318),
.B(n_1303),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1426),
.B(n_1436),
.Y(n_1464)
);

BUFx4f_ASAP7_75t_SL g1465 ( 
.A(n_1396),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1422),
.Y(n_1466)
);

O2A1O1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1454),
.A2(n_1462),
.B(n_1343),
.C(n_1432),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1459),
.B(n_1374),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1361),
.A2(n_1363),
.B(n_1367),
.Y(n_1469)
);

O2A1O1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1454),
.A2(n_1430),
.B(n_1348),
.C(n_1455),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1451),
.B(n_1375),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1365),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1451),
.B(n_1375),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1364),
.B(n_1372),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1368),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1374),
.B(n_1352),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1352),
.B(n_1345),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_SL g1478 ( 
.A1(n_1421),
.A2(n_1442),
.B(n_1417),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1428),
.Y(n_1479)
);

AND2x4_ASAP7_75t_SL g1480 ( 
.A(n_1437),
.B(n_1350),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1386),
.B(n_1355),
.Y(n_1481)
);

NOR2xp67_ASAP7_75t_L g1482 ( 
.A(n_1377),
.B(n_1458),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1361),
.A2(n_1363),
.B(n_1367),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1386),
.B(n_1418),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1364),
.A2(n_1435),
.B1(n_1439),
.B2(n_1441),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1354),
.B(n_1391),
.Y(n_1486)
);

CKINVDCx14_ASAP7_75t_R g1487 ( 
.A(n_1437),
.Y(n_1487)
);

O2A1O1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1348),
.A2(n_1448),
.B(n_1417),
.C(n_1455),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1410),
.Y(n_1489)
);

OA21x2_ASAP7_75t_L g1490 ( 
.A1(n_1340),
.A2(n_1390),
.B(n_1388),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1379),
.B(n_1366),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1366),
.A2(n_1420),
.B1(n_1456),
.B2(n_1413),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1357),
.B(n_1453),
.Y(n_1493)
);

OA21x2_ASAP7_75t_L g1494 ( 
.A1(n_1371),
.A2(n_1452),
.B(n_1461),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1403),
.A2(n_1359),
.B1(n_1411),
.B2(n_1397),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1370),
.B(n_1356),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1403),
.A2(n_1379),
.B1(n_1353),
.B2(n_1415),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1414),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1392),
.A2(n_1400),
.B1(n_1404),
.B2(n_1384),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1392),
.A2(n_1445),
.B1(n_1405),
.B2(n_1385),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1392),
.A2(n_1445),
.B1(n_1382),
.B2(n_1376),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1410),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1393),
.B(n_1443),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1445),
.A2(n_1394),
.B1(n_1457),
.B2(n_1389),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1362),
.Y(n_1505)
);

AOI221xp5_ASAP7_75t_L g1506 ( 
.A1(n_1438),
.A2(n_1444),
.B1(n_1380),
.B2(n_1387),
.C(n_1425),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1449),
.B(n_1450),
.Y(n_1507)
);

NOR2xp67_ASAP7_75t_L g1508 ( 
.A(n_1351),
.B(n_1434),
.Y(n_1508)
);

AOI21x1_ASAP7_75t_SL g1509 ( 
.A1(n_1349),
.A2(n_1369),
.B(n_1416),
.Y(n_1509)
);

CKINVDCx16_ASAP7_75t_R g1510 ( 
.A(n_1433),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1429),
.A2(n_1416),
.B1(n_1378),
.B2(n_1440),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1423),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1416),
.A2(n_1440),
.B1(n_1378),
.B2(n_1449),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1449),
.B(n_1463),
.Y(n_1514)
);

O2A1O1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1380),
.A2(n_1450),
.B(n_1406),
.C(n_1402),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1398),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1440),
.A2(n_1407),
.B1(n_1360),
.B2(n_1341),
.Y(n_1517)
);

O2A1O1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1341),
.A2(n_1460),
.B(n_1427),
.C(n_1347),
.Y(n_1518)
);

OA21x2_ASAP7_75t_L g1519 ( 
.A1(n_1419),
.A2(n_1424),
.B(n_1446),
.Y(n_1519)
);

O2A1O1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1344),
.A2(n_1358),
.B(n_1412),
.C(n_1447),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1412),
.B(n_1358),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1408),
.Y(n_1522)
);

BUFx3_ASAP7_75t_L g1523 ( 
.A(n_1396),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1401),
.Y(n_1524)
);

OAI211xp5_ASAP7_75t_L g1525 ( 
.A1(n_1383),
.A2(n_1373),
.B(n_1409),
.C(n_1399),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1395),
.B(n_1346),
.Y(n_1526)
);

OA22x2_ASAP7_75t_L g1527 ( 
.A1(n_1395),
.A2(n_1431),
.B1(n_1447),
.B2(n_813),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1431),
.B(n_1430),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_SL g1529 ( 
.A1(n_1451),
.A2(n_1198),
.B(n_1337),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1430),
.B(n_1432),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1381),
.A2(n_1320),
.B(n_1278),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1430),
.B(n_1432),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1364),
.A2(n_1277),
.B1(n_1210),
.B2(n_1430),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1364),
.A2(n_1277),
.B1(n_1210),
.B2(n_1430),
.Y(n_1534)
);

A2O1A1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1430),
.A2(n_1284),
.B(n_1432),
.C(n_1451),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1430),
.B(n_1432),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1430),
.B(n_1432),
.Y(n_1537)
);

O2A1O1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1454),
.A2(n_1284),
.B(n_1343),
.C(n_1462),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1364),
.A2(n_1277),
.B1(n_1210),
.B2(n_1430),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1342),
.B(n_378),
.Y(n_1540)
);

BUFx2_ASAP7_75t_SL g1541 ( 
.A(n_1353),
.Y(n_1541)
);

OR2x6_ASAP7_75t_L g1542 ( 
.A(n_1386),
.B(n_1381),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1426),
.B(n_1436),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_SL g1544 ( 
.A1(n_1451),
.A2(n_1198),
.B(n_1337),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1386),
.B(n_1355),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1522),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1521),
.B(n_1526),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1516),
.Y(n_1548)
);

AO21x1_ASAP7_75t_SL g1549 ( 
.A1(n_1471),
.A2(n_1473),
.B(n_1491),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1498),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1524),
.B(n_1542),
.Y(n_1551)
);

AOI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1467),
.A2(n_1538),
.B1(n_1470),
.B2(n_1488),
.C(n_1535),
.Y(n_1552)
);

OR2x6_ASAP7_75t_L g1553 ( 
.A(n_1542),
.B(n_1531),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1518),
.A2(n_1469),
.B(n_1483),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1472),
.Y(n_1555)
);

AOI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1497),
.A2(n_1513),
.B(n_1503),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1507),
.B(n_1514),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_SL g1558 ( 
.A1(n_1538),
.A2(n_1488),
.B(n_1470),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1507),
.B(n_1514),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1489),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1528),
.B(n_1502),
.Y(n_1561)
);

AO21x2_ASAP7_75t_L g1562 ( 
.A1(n_1471),
.A2(n_1473),
.B(n_1491),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1527),
.B(n_1542),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1490),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1490),
.B(n_1476),
.Y(n_1565)
);

AO21x2_ASAP7_75t_L g1566 ( 
.A1(n_1525),
.A2(n_1478),
.B(n_1474),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1519),
.B(n_1506),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1494),
.Y(n_1568)
);

OA21x2_ASAP7_75t_L g1569 ( 
.A1(n_1474),
.A2(n_1525),
.B(n_1499),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1494),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1477),
.B(n_1520),
.Y(n_1571)
);

NAND3xp33_ASAP7_75t_L g1572 ( 
.A(n_1533),
.B(n_1539),
.C(n_1534),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1511),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1508),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1481),
.B(n_1484),
.Y(n_1575)
);

BUFx5_ASAP7_75t_L g1576 ( 
.A(n_1484),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1501),
.Y(n_1577)
);

AO21x2_ASAP7_75t_L g1578 ( 
.A1(n_1492),
.A2(n_1520),
.B(n_1515),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_1487),
.Y(n_1579)
);

OR2x6_ASAP7_75t_L g1580 ( 
.A(n_1500),
.B(n_1544),
.Y(n_1580)
);

OR2x6_ASAP7_75t_L g1581 ( 
.A(n_1529),
.B(n_1545),
.Y(n_1581)
);

INVxp67_ASAP7_75t_SL g1582 ( 
.A(n_1496),
.Y(n_1582)
);

AO21x2_ASAP7_75t_L g1583 ( 
.A1(n_1530),
.A2(n_1536),
.B(n_1537),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1468),
.B(n_1532),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1537),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1548),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1548),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1560),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1555),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1561),
.B(n_1493),
.Y(n_1590)
);

INVx4_ASAP7_75t_L g1591 ( 
.A(n_1581),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1565),
.B(n_1557),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1561),
.B(n_1495),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1583),
.B(n_1585),
.Y(n_1594)
);

OA21x2_ASAP7_75t_L g1595 ( 
.A1(n_1554),
.A2(n_1485),
.B(n_1509),
.Y(n_1595)
);

INVxp67_ASAP7_75t_SL g1596 ( 
.A(n_1564),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1565),
.B(n_1557),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1583),
.B(n_1486),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1565),
.B(n_1543),
.Y(n_1599)
);

NOR2x1_ASAP7_75t_L g1600 ( 
.A(n_1583),
.B(n_1517),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1559),
.B(n_1464),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1558),
.B(n_1504),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1572),
.B(n_1479),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_1551),
.Y(n_1604)
);

INVx2_ASAP7_75t_SL g1605 ( 
.A(n_1574),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1551),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1568),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1576),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1546),
.B(n_1568),
.Y(n_1609)
);

INVx3_ASAP7_75t_L g1610 ( 
.A(n_1568),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1547),
.B(n_1475),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1602),
.A2(n_1572),
.B1(n_1552),
.B2(n_1562),
.Y(n_1612)
);

INVxp67_ASAP7_75t_SL g1613 ( 
.A(n_1596),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1588),
.Y(n_1614)
);

OR2x6_ASAP7_75t_L g1615 ( 
.A(n_1591),
.B(n_1581),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_L g1616 ( 
.A(n_1602),
.B(n_1552),
.C(n_1573),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1589),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1589),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1599),
.B(n_1575),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1609),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1604),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1598),
.B(n_1571),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1598),
.B(n_1571),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1586),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_SL g1625 ( 
.A1(n_1603),
.A2(n_1566),
.B1(n_1569),
.B2(n_1578),
.Y(n_1625)
);

BUFx12f_ASAP7_75t_L g1626 ( 
.A(n_1590),
.Y(n_1626)
);

NAND2xp33_ASAP7_75t_R g1627 ( 
.A(n_1595),
.B(n_1569),
.Y(n_1627)
);

OAI211xp5_ASAP7_75t_L g1628 ( 
.A1(n_1600),
.A2(n_1569),
.B(n_1573),
.C(n_1556),
.Y(n_1628)
);

INVx4_ASAP7_75t_SL g1629 ( 
.A(n_1605),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1599),
.B(n_1575),
.Y(n_1630)
);

A2O1A1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1603),
.A2(n_1600),
.B(n_1563),
.C(n_1571),
.Y(n_1631)
);

AO21x2_ASAP7_75t_L g1632 ( 
.A1(n_1596),
.A2(n_1564),
.B(n_1570),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_L g1633 ( 
.A(n_1594),
.B(n_1569),
.C(n_1577),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1593),
.A2(n_1562),
.B1(n_1549),
.B2(n_1566),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1593),
.A2(n_1562),
.B1(n_1549),
.B2(n_1566),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1592),
.B(n_1582),
.Y(n_1636)
);

OAI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1593),
.A2(n_1580),
.B1(n_1482),
.B2(n_1553),
.C(n_1540),
.Y(n_1637)
);

OAI211xp5_ASAP7_75t_L g1638 ( 
.A1(n_1595),
.A2(n_1569),
.B(n_1556),
.C(n_1577),
.Y(n_1638)
);

INVx3_ASAP7_75t_L g1639 ( 
.A(n_1609),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1611),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_L g1641 ( 
.A(n_1595),
.B(n_1553),
.C(n_1567),
.Y(n_1641)
);

OAI321xp33_ASAP7_75t_L g1642 ( 
.A1(n_1586),
.A2(n_1580),
.A3(n_1553),
.B1(n_1581),
.B2(n_1563),
.C(n_1567),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1587),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1588),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1624),
.Y(n_1645)
);

INVx4_ASAP7_75t_SL g1646 ( 
.A(n_1615),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1632),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1643),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1632),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1614),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1617),
.Y(n_1651)
);

NAND3xp33_ASAP7_75t_L g1652 ( 
.A(n_1616),
.B(n_1595),
.C(n_1553),
.Y(n_1652)
);

BUFx3_ASAP7_75t_L g1653 ( 
.A(n_1626),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1641),
.A2(n_1610),
.B(n_1607),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1620),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1620),
.B(n_1639),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1618),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1639),
.B(n_1592),
.Y(n_1658)
);

NAND3xp33_ASAP7_75t_SL g1659 ( 
.A(n_1612),
.B(n_1579),
.C(n_1550),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1619),
.B(n_1597),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1630),
.B(n_1597),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1614),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1644),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1644),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1621),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1629),
.Y(n_1666)
);

OR2x6_ASAP7_75t_L g1667 ( 
.A(n_1615),
.B(n_1580),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1629),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1613),
.Y(n_1669)
);

INVx5_ASAP7_75t_L g1670 ( 
.A(n_1615),
.Y(n_1670)
);

INVx4_ASAP7_75t_SL g1671 ( 
.A(n_1640),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1612),
.B(n_1584),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1654),
.B(n_1631),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1669),
.B(n_1622),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1645),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1653),
.B(n_1625),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1653),
.B(n_1523),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1647),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1669),
.B(n_1623),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1647),
.Y(n_1680)
);

INVxp67_ASAP7_75t_L g1681 ( 
.A(n_1650),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1647),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1659),
.A2(n_1625),
.B1(n_1553),
.B2(n_1566),
.Y(n_1683)
);

OAI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1659),
.A2(n_1633),
.B(n_1628),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_SL g1685 ( 
.A(n_1653),
.B(n_1642),
.Y(n_1685)
);

NOR2x1_ASAP7_75t_L g1686 ( 
.A(n_1652),
.B(n_1638),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1665),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1646),
.B(n_1608),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1649),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1671),
.B(n_1606),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1662),
.B(n_1601),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1671),
.B(n_1606),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1649),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1650),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1671),
.B(n_1606),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1648),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1649),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1671),
.B(n_1636),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1658),
.B(n_1656),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1670),
.B(n_1634),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1658),
.B(n_1656),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1664),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1646),
.B(n_1608),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1694),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1699),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1687),
.B(n_1672),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1687),
.B(n_1660),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1698),
.B(n_1690),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1694),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1676),
.B(n_1660),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1686),
.B(n_1646),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1686),
.B(n_1646),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1698),
.B(n_1666),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1696),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1676),
.B(n_1660),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1696),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1699),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1678),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1696),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1702),
.B(n_1664),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1684),
.B(n_1661),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1699),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1698),
.B(n_1666),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1690),
.B(n_1692),
.Y(n_1724)
);

A2O1A1Ixp33_ASAP7_75t_L g1725 ( 
.A1(n_1684),
.A2(n_1652),
.B(n_1634),
.C(n_1635),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_L g1726 ( 
.A(n_1685),
.B(n_1627),
.C(n_1635),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1677),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1690),
.B(n_1666),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1692),
.B(n_1668),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1685),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1692),
.B(n_1668),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1702),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1675),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1695),
.B(n_1668),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1674),
.B(n_1662),
.Y(n_1735)
);

OR2x6_ASAP7_75t_L g1736 ( 
.A(n_1700),
.B(n_1688),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1683),
.A2(n_1637),
.B1(n_1667),
.B2(n_1580),
.Y(n_1737)
);

AO221x1_ASAP7_75t_L g1738 ( 
.A1(n_1681),
.A2(n_1655),
.B1(n_1663),
.B2(n_1651),
.C(n_1657),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1675),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1701),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1727),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1720),
.B(n_1681),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1738),
.Y(n_1743)
);

INVx1_ASAP7_75t_SL g1744 ( 
.A(n_1727),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1708),
.B(n_1695),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1720),
.B(n_1674),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1727),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1704),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1708),
.B(n_1695),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1730),
.B(n_1677),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1724),
.B(n_1673),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1732),
.B(n_1679),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1724),
.B(n_1673),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1711),
.B(n_1465),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1711),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1711),
.B(n_1466),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1732),
.B(n_1691),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1721),
.B(n_1691),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1711),
.B(n_1480),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1712),
.B(n_1683),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1713),
.B(n_1673),
.Y(n_1761)
);

BUFx2_ASAP7_75t_SL g1762 ( 
.A(n_1712),
.Y(n_1762)
);

AO21x2_ASAP7_75t_L g1763 ( 
.A1(n_1738),
.A2(n_1700),
.B(n_1680),
.Y(n_1763)
);

INVx1_ASAP7_75t_SL g1764 ( 
.A(n_1712),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1713),
.B(n_1688),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1718),
.Y(n_1766)
);

AOI21xp33_ASAP7_75t_SL g1767 ( 
.A1(n_1760),
.A2(n_1726),
.B(n_1712),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1744),
.B(n_1723),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1744),
.B(n_1723),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1741),
.B(n_1706),
.Y(n_1770)
);

INVx2_ASAP7_75t_SL g1771 ( 
.A(n_1765),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1756),
.B(n_1707),
.Y(n_1772)
);

AOI221x1_ASAP7_75t_SL g1773 ( 
.A1(n_1743),
.A2(n_1726),
.B1(n_1710),
.B2(n_1715),
.C(n_1704),
.Y(n_1773)
);

NAND3xp33_ASAP7_75t_L g1774 ( 
.A(n_1747),
.B(n_1725),
.C(n_1736),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1763),
.A2(n_1737),
.B1(n_1736),
.B2(n_1703),
.Y(n_1775)
);

BUFx6f_ASAP7_75t_L g1776 ( 
.A(n_1754),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1742),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1763),
.A2(n_1736),
.B(n_1709),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1750),
.B(n_1512),
.Y(n_1779)
);

XNOR2x2_ASAP7_75t_L g1780 ( 
.A(n_1755),
.B(n_1709),
.Y(n_1780)
);

INVxp33_ASAP7_75t_L g1781 ( 
.A(n_1759),
.Y(n_1781)
);

AOI21xp33_ASAP7_75t_L g1782 ( 
.A1(n_1763),
.A2(n_1736),
.B(n_1729),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1742),
.Y(n_1783)
);

INVxp67_ASAP7_75t_L g1784 ( 
.A(n_1762),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1745),
.A2(n_1736),
.B1(n_1731),
.B2(n_1734),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1743),
.A2(n_1729),
.B(n_1728),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1777),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1781),
.B(n_1755),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1783),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1771),
.B(n_1745),
.Y(n_1790)
);

NAND2xp33_ASAP7_75t_R g1791 ( 
.A(n_1767),
.B(n_1505),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1773),
.B(n_1764),
.Y(n_1792)
);

INVxp67_ASAP7_75t_SL g1793 ( 
.A(n_1780),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1784),
.B(n_1764),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1768),
.B(n_1762),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1769),
.B(n_1761),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1776),
.B(n_1758),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1776),
.B(n_1746),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1776),
.B(n_1749),
.Y(n_1799)
);

AOI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1793),
.A2(n_1774),
.B1(n_1772),
.B2(n_1743),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1793),
.B(n_1770),
.Y(n_1801)
);

NAND4xp25_ASAP7_75t_L g1802 ( 
.A(n_1788),
.B(n_1775),
.C(n_1785),
.D(n_1786),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1799),
.B(n_1749),
.Y(n_1803)
);

OAI31xp33_ASAP7_75t_L g1804 ( 
.A1(n_1792),
.A2(n_1782),
.A3(n_1778),
.B(n_1751),
.Y(n_1804)
);

AOI221xp5_ASAP7_75t_L g1805 ( 
.A1(n_1798),
.A2(n_1748),
.B1(n_1757),
.B2(n_1761),
.C(n_1751),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1797),
.B(n_1746),
.Y(n_1806)
);

AOI32xp33_ASAP7_75t_L g1807 ( 
.A1(n_1790),
.A2(n_1753),
.A3(n_1765),
.B1(n_1748),
.B2(n_1734),
.Y(n_1807)
);

AOI211xp5_ASAP7_75t_SL g1808 ( 
.A1(n_1794),
.A2(n_1779),
.B(n_1753),
.C(n_1752),
.Y(n_1808)
);

NAND4xp75_ASAP7_75t_L g1809 ( 
.A(n_1787),
.B(n_1766),
.C(n_1731),
.D(n_1728),
.Y(n_1809)
);

NAND3xp33_ASAP7_75t_L g1810 ( 
.A(n_1795),
.B(n_1752),
.C(n_1766),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1800),
.B(n_1789),
.Y(n_1811)
);

XNOR2xp5_ASAP7_75t_L g1812 ( 
.A(n_1802),
.B(n_1796),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1808),
.B(n_1705),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1803),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1810),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1809),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1815),
.B(n_1804),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1816),
.B(n_1801),
.Y(n_1818)
);

NOR2x1_ASAP7_75t_L g1819 ( 
.A(n_1811),
.B(n_1806),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1814),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1813),
.B(n_1805),
.Y(n_1821)
);

INVx1_ASAP7_75t_SL g1822 ( 
.A(n_1812),
.Y(n_1822)
);

NAND3xp33_ASAP7_75t_L g1823 ( 
.A(n_1815),
.B(n_1807),
.C(n_1791),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1822),
.B(n_1705),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1818),
.Y(n_1825)
);

NOR2xp67_ASAP7_75t_L g1826 ( 
.A(n_1823),
.B(n_1820),
.Y(n_1826)
);

XNOR2x2_ASAP7_75t_SL g1827 ( 
.A(n_1821),
.B(n_1735),
.Y(n_1827)
);

AOI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1819),
.A2(n_1717),
.B1(n_1740),
.B2(n_1722),
.Y(n_1828)
);

NOR3xp33_ASAP7_75t_L g1829 ( 
.A(n_1817),
.B(n_1510),
.C(n_1766),
.Y(n_1829)
);

AOI21xp33_ASAP7_75t_L g1830 ( 
.A1(n_1824),
.A2(n_1825),
.B(n_1826),
.Y(n_1830)
);

OAI21xp5_ASAP7_75t_SL g1831 ( 
.A1(n_1828),
.A2(n_1722),
.B(n_1717),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1827),
.Y(n_1832)
);

NAND5xp2_ASAP7_75t_L g1833 ( 
.A(n_1832),
.B(n_1829),
.C(n_1733),
.D(n_1739),
.E(n_1714),
.Y(n_1833)
);

AOI322xp5_ASAP7_75t_L g1834 ( 
.A1(n_1833),
.A2(n_1830),
.A3(n_1740),
.B1(n_1831),
.B2(n_1718),
.C1(n_1714),
.C2(n_1719),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1834),
.Y(n_1835)
);

OR3x2_ASAP7_75t_L g1836 ( 
.A(n_1834),
.B(n_1739),
.C(n_1733),
.Y(n_1836)
);

OAI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1835),
.A2(n_1718),
.B(n_1716),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1836),
.B(n_1701),
.Y(n_1838)
);

OAI22xp5_ASAP7_75t_SL g1839 ( 
.A1(n_1837),
.A2(n_1541),
.B1(n_1719),
.B2(n_1716),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1838),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1840),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1841),
.A2(n_1839),
.B1(n_1678),
.B2(n_1680),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1842),
.B(n_1678),
.Y(n_1843)
);

AOI322xp5_ASAP7_75t_L g1844 ( 
.A1(n_1843),
.A2(n_1682),
.A3(n_1680),
.B1(n_1678),
.B2(n_1689),
.C1(n_1693),
.C2(n_1697),
.Y(n_1844)
);

AOI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1844),
.A2(n_1697),
.B1(n_1680),
.B2(n_1693),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1845),
.A2(n_1697),
.B1(n_1689),
.B2(n_1693),
.Y(n_1846)
);


endmodule