module fake_jpeg_10541_n_336 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_40),
.B(n_31),
.Y(n_64)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_46),
.Y(n_51)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_8),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_60),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_56),
.B1(n_68),
.B2(n_30),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_34),
.B(n_32),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_42),
.B(n_18),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_57),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_32),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_37),
.A2(n_30),
.B1(n_29),
.B2(n_24),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_70),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_72),
.A2(n_82),
.B1(n_92),
.B2(n_62),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_40),
.B1(n_30),
.B2(n_41),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_97),
.B1(n_69),
.B2(n_25),
.Y(n_102)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_77),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_26),
.B1(n_29),
.B2(n_21),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_19),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_59),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_79),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_85),
.Y(n_103)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_60),
.Y(n_124)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_18),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_63),
.B(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_34),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_50),
.B(n_33),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_34),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_34),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_49),
.A2(n_19),
.B1(n_20),
.B2(n_33),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_106),
.Y(n_140)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_17),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_118),
.Y(n_131)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_109),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_71),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_107),
.Y(n_150)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_115),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_72),
.A2(n_49),
.B1(n_62),
.B2(n_52),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_76),
.B1(n_73),
.B2(n_97),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_19),
.C(n_20),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_16),
.Y(n_143)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_126),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_75),
.B(n_81),
.Y(n_133)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_105),
.B1(n_109),
.B2(n_78),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_0),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_136),
.B1(n_145),
.B2(n_148),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_133),
.A2(n_134),
.B(n_138),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_92),
.B(n_84),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_119),
.A2(n_78),
.B1(n_83),
.B2(n_80),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_32),
.B(n_34),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_44),
.C(n_58),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_146),
.C(n_100),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_83),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_143),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_83),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_153),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_48),
.C(n_36),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_121),
.A2(n_78),
.B1(n_80),
.B2(n_54),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_106),
.A2(n_54),
.B1(n_39),
.B2(n_20),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_152),
.A2(n_154),
.B1(n_113),
.B2(n_126),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_0),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_39),
.B1(n_19),
.B2(n_20),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_155),
.B(n_156),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_131),
.B(n_110),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_157),
.B(n_159),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_144),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_162),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_118),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_164),
.C(n_179),
.Y(n_189)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_114),
.B1(n_101),
.B2(n_122),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_173),
.B1(n_135),
.B2(n_123),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_103),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_127),
.A2(n_111),
.B1(n_103),
.B2(n_113),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_165),
.A2(n_154),
.B1(n_151),
.B2(n_139),
.Y(n_199)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_167),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_131),
.B(n_108),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_125),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_168),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_169),
.A2(n_177),
.B(n_153),
.Y(n_200)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_170),
.A2(n_178),
.B1(n_180),
.B2(n_183),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_143),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_130),
.A2(n_113),
.B1(n_123),
.B2(n_80),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_132),
.B1(n_148),
.B2(n_128),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_150),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_100),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_SL g181 ( 
.A(n_145),
.B(n_108),
.C(n_104),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_181),
.A2(n_128),
.B1(n_135),
.B2(n_130),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_102),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_182),
.Y(n_193)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_185),
.A2(n_187),
.B1(n_190),
.B2(n_205),
.Y(n_218)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_197),
.C(n_158),
.Y(n_224)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_194),
.B(n_203),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_196),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_151),
.C(n_139),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_199),
.A2(n_206),
.B1(n_174),
.B2(n_194),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_202),
.B(n_210),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_153),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_167),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_204),
.B(n_9),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_143),
.B1(n_104),
.B2(n_91),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_175),
.A2(n_91),
.B1(n_61),
.B2(n_48),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_212),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_171),
.A2(n_115),
.B(n_96),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_209),
.A2(n_160),
.B(n_178),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_162),
.A2(n_32),
.B(n_91),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_175),
.B1(n_180),
.B2(n_166),
.Y(n_214)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_214),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_179),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_221),
.C(n_224),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_217),
.A2(n_232),
.B1(n_236),
.B2(n_237),
.Y(n_253)
);

BUFx8_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_220),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_172),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_209),
.B(n_187),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_192),
.B(n_171),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_210),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_164),
.C(n_158),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_202),
.C(n_4),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_211),
.A2(n_177),
.B1(n_182),
.B2(n_181),
.Y(n_228)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_226),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_230)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_235),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_193),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_185),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_233)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_195),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_193),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_199),
.A2(n_203),
.B1(n_207),
.B2(n_191),
.Y(n_237)
);

INVxp33_ASAP7_75t_SL g238 ( 
.A(n_208),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_238),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_241),
.A2(n_259),
.B(n_243),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_201),
.Y(n_244)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_201),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

XNOR2x1_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_215),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_254),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_186),
.Y(n_250)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_252),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_219),
.B(n_200),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_220),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_5),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_260),
.C(n_236),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_222),
.A2(n_202),
.B(n_11),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_3),
.C(n_5),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_231),
.B1(n_218),
.B2(n_228),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_264),
.A2(n_273),
.B1(n_242),
.B2(n_248),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_216),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_279),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_224),
.C(n_225),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_274),
.C(n_277),
.Y(n_282)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_244),
.B(n_217),
.CI(n_232),
.CON(n_270),
.SN(n_270)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_240),
.A2(n_213),
.B1(n_233),
.B2(n_7),
.Y(n_271)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_272),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_261),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_12),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_12),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_12),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_278),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_276),
.A2(n_249),
.B1(n_240),
.B2(n_255),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_280),
.A2(n_284),
.B1(n_285),
.B2(n_279),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_262),
.A2(n_253),
.B1(n_255),
.B2(n_243),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_253),
.B1(n_248),
.B2(n_242),
.Y(n_285)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_264),
.B(n_241),
.CI(n_259),
.CON(n_287),
.SN(n_287)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_288),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_277),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_239),
.B(n_257),
.Y(n_292)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_292),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_298),
.B(n_306),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_239),
.B(n_275),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_301),
.C(n_305),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_295),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_269),
.C(n_266),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_303),
.B(n_307),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_294),
.A2(n_256),
.B1(n_273),
.B2(n_272),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_304),
.A2(n_280),
.B1(n_283),
.B2(n_287),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_274),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_291),
.B(n_258),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_256),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_293),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_308),
.B(n_311),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_282),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_314),
.Y(n_320)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_313),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_299),
.B(n_258),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_282),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_265),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_324),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_317),
.A2(n_302),
.B(n_297),
.Y(n_321)
);

AO21x1_ASAP7_75t_L g329 ( 
.A1(n_321),
.A2(n_322),
.B(n_325),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_296),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_263),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_317),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_318),
.A2(n_312),
.B1(n_310),
.B2(n_287),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_326),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_323),
.A2(n_265),
.B(n_260),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_328),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_320),
.C(n_323),
.Y(n_332)
);

OAI321xp33_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_327),
.A3(n_329),
.B1(n_330),
.B2(n_11),
.C(n_14),
.Y(n_333)
);

OAI21xp33_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_9),
.B(n_10),
.Y(n_334)
);

O2A1O1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_6),
.B(n_10),
.C(n_15),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_16),
.B(n_333),
.Y(n_336)
);


endmodule