module fake_jpeg_9627_n_126 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_96;

INVx13_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_0),
.B(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_30),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_63),
.Y(n_69)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_61),
.B(n_64),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_68),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_86),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_38),
.B1(n_55),
.B2(n_44),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_102)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_80),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_63),
.B(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_83),
.B(n_88),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_0),
.Y(n_87)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_89),
.CI(n_90),
.CON(n_94),
.SN(n_94)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_56),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_1),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_50),
.A3(n_47),
.B1(n_39),
.B2(n_43),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_101),
.B1(n_102),
.B2(n_78),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_46),
.B1(n_48),
.B2(n_51),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_99),
.B1(n_103),
.B2(n_85),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_49),
.B1(n_56),
.B2(n_52),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_75),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_110),
.B1(n_101),
.B2(n_69),
.Y(n_111)
);

OAI32xp33_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_110),
.A3(n_107),
.B1(n_94),
.B2(n_71),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_112),
.A2(n_94),
.B(n_105),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_113),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_114),
.A2(n_103),
.B1(n_104),
.B2(n_89),
.Y(n_115)
);

AOI321xp33_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_93),
.A3(n_106),
.B1(n_72),
.B2(n_108),
.C(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_98),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_95),
.B1(n_5),
.B2(n_6),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_4),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_119),
.A2(n_100),
.B1(n_7),
.B2(n_9),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_8),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_10),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_11),
.Y(n_123)
);

OAI321xp33_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_12),
.A3(n_16),
.B1(n_17),
.B2(n_18),
.C(n_20),
.Y(n_124)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_124),
.B(n_21),
.CI(n_24),
.CON(n_125),
.SN(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_26),
.B(n_27),
.Y(n_126)
);


endmodule