module fake_netlist_6_27_n_1738 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1738);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1738;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_133),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_29),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_9),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_126),
.Y(n_160)
);

BUFx2_ASAP7_75t_R g161 ( 
.A(n_81),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_149),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_53),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_34),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_95),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_89),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_83),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_20),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_86),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_16),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_33),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_42),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_75),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_128),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_59),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_82),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_125),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_92),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_62),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_6),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_2),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_118),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_106),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_70),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_63),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_67),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_61),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_20),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_14),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_145),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_7),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_21),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_36),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_55),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_30),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_101),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_74),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_34),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_87),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_109),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_56),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_5),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_60),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_153),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_51),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_79),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_13),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_48),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_10),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_102),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_40),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_33),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_57),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_115),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_112),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_143),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_138),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_132),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_98),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_90),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_72),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_12),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_44),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_141),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_45),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_22),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_53),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_103),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_19),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_42),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_38),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_32),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_37),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_108),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_27),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_121),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_100),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_52),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_39),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_40),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_134),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_94),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_43),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_64),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_117),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_96),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_130),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_110),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_15),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_58),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_111),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_16),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_154),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_38),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_2),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_30),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_93),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_29),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_150),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_48),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_19),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_4),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_135),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_137),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_21),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_47),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_142),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_7),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_17),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_43),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_32),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_10),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_124),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_85),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_123),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_80),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_46),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_31),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_36),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_146),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_104),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_54),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_71),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_136),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_1),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_24),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_14),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_52),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_0),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_152),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_0),
.Y(n_301)
);

BUFx5_ASAP7_75t_L g302 ( 
.A(n_51),
.Y(n_302)
);

BUFx10_ASAP7_75t_L g303 ( 
.A(n_23),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_114),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_27),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_41),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_24),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_155),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_9),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_17),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_183),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_181),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_302),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_302),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_182),
.Y(n_317)
);

INVxp33_ASAP7_75t_SL g318 ( 
.A(n_158),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_302),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_302),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_184),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_303),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_212),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_212),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_212),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_211),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_212),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_158),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_212),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_185),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_165),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_168),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_192),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_240),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_278),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_278),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_240),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_244),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_303),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_240),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_240),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_244),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_240),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_278),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_237),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_237),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_189),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_266),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_266),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_191),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_159),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_186),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_213),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_200),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_165),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_207),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_219),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_303),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_195),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_196),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_199),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_168),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_221),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_222),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_235),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_205),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_230),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_210),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_214),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_241),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_216),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_248),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_243),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_250),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_253),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_279),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_227),
.Y(n_380)
);

INVxp33_ASAP7_75t_SL g381 ( 
.A(n_177),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_325),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_325),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_203),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_344),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_326),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_344),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_344),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_311),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_344),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_326),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_340),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_344),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_327),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_329),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_340),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_340),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_337),
.B(n_203),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_313),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_323),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_332),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_314),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_314),
.Y(n_406)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_337),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_329),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_334),
.B(n_273),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_312),
.A2(n_262),
.B1(n_176),
.B2(n_201),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_331),
.B(n_273),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_335),
.A2(n_236),
.B1(n_288),
.B2(n_265),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_336),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_315),
.Y(n_415)
);

BUFx8_ASAP7_75t_L g416 ( 
.A(n_334),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_318),
.A2(n_166),
.B1(n_242),
.B2(n_174),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_315),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_316),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_317),
.A2(n_239),
.B1(n_197),
.B2(n_307),
.Y(n_420)
);

BUFx8_ASAP7_75t_L g421 ( 
.A(n_334),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_316),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_346),
.B(n_231),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_336),
.B(n_157),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_319),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_376),
.B(n_171),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_339),
.B(n_157),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_346),
.B(n_231),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_319),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_320),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_342),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_342),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_343),
.B(n_160),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_343),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_324),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_338),
.B(n_298),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_345),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_345),
.B(n_160),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_349),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_L g441 ( 
.A(n_338),
.B(n_298),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_320),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_368),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_321),
.B(n_162),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_321),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_322),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_403),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_436),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_409),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_403),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_384),
.A2(n_444),
.B1(n_446),
.B2(n_445),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_445),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_416),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_385),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_403),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_390),
.B(n_376),
.Y(n_457)
);

CKINVDCx6p67_ASAP7_75t_R g458 ( 
.A(n_426),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_446),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_401),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_403),
.Y(n_461)
);

NAND3xp33_ASAP7_75t_L g462 ( 
.A(n_444),
.B(n_322),
.C(n_370),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_405),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_401),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_401),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_402),
.B(n_352),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_405),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_413),
.A2(n_255),
.B1(n_308),
.B2(n_202),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_415),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_R g470 ( 
.A(n_436),
.B(n_333),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_404),
.B(n_362),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_385),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_405),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_416),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_405),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_384),
.A2(n_381),
.B1(n_296),
.B2(n_301),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_409),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_415),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_415),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_419),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_409),
.B(n_350),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_406),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_418),
.B(n_363),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_418),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_385),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_R g486 ( 
.A(n_440),
.B(n_364),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_419),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_419),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_406),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_411),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_385),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_426),
.B(n_369),
.Y(n_492)
);

INVx5_ASAP7_75t_L g493 ( 
.A(n_425),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g494 ( 
.A(n_423),
.B(n_378),
.C(n_354),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_418),
.B(n_371),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_418),
.B(n_372),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_418),
.B(n_374),
.Y(n_497)
);

INVxp33_ASAP7_75t_L g498 ( 
.A(n_411),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_406),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_425),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_406),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_436),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_400),
.A2(n_295),
.B1(n_305),
.B2(n_287),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_431),
.Y(n_504)
);

NAND2xp33_ASAP7_75t_R g505 ( 
.A(n_437),
.B(n_162),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_416),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_416),
.B(n_341),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_425),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_392),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_422),
.Y(n_510)
);

OR2x6_ASAP7_75t_L g511 ( 
.A(n_437),
.B(n_156),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_400),
.A2(n_280),
.B1(n_306),
.B2(n_281),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_431),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_422),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_423),
.B(n_350),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_431),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_431),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_422),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_442),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_400),
.A2(n_330),
.B1(n_358),
.B2(n_244),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_385),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_442),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_424),
.B(n_361),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_442),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_L g525 ( 
.A(n_424),
.B(n_428),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_428),
.B(n_294),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_382),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_416),
.B(n_161),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_421),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_392),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_434),
.B(n_439),
.Y(n_531)
);

OR2x6_ASAP7_75t_L g532 ( 
.A(n_437),
.B(n_163),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_417),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_421),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_392),
.Y(n_535)
);

OR2x6_ASAP7_75t_L g536 ( 
.A(n_400),
.B(n_170),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_392),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_385),
.Y(n_538)
);

INVx6_ASAP7_75t_L g539 ( 
.A(n_421),
.Y(n_539)
);

OAI22xp33_ASAP7_75t_SL g540 ( 
.A1(n_434),
.A2(n_439),
.B1(n_413),
.B2(n_417),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_382),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_443),
.B(n_351),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_383),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_L g544 ( 
.A1(n_443),
.A2(n_232),
.B1(n_309),
.B2(n_217),
.Y(n_544)
);

AND3x2_ASAP7_75t_L g545 ( 
.A(n_423),
.B(n_289),
.C(n_175),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_383),
.Y(n_546)
);

BUFx6f_ASAP7_75t_SL g547 ( 
.A(n_400),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_387),
.Y(n_548)
);

AOI21x1_ASAP7_75t_L g549 ( 
.A1(n_412),
.A2(n_187),
.B(n_173),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_387),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_421),
.B(n_171),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_395),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_395),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_396),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_407),
.B(n_223),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_396),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_397),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_397),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_408),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_421),
.B(n_171),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_408),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_443),
.B(n_351),
.Y(n_562)
);

NAND3xp33_ASAP7_75t_L g563 ( 
.A(n_429),
.B(n_354),
.C(n_353),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_443),
.B(n_328),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_443),
.B(n_193),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_407),
.B(n_225),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_407),
.B(n_234),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_410),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_410),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_414),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_420),
.B(n_193),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_414),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_R g573 ( 
.A(n_441),
.B(n_356),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_407),
.B(n_380),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_427),
.Y(n_575)
);

INVx5_ASAP7_75t_L g576 ( 
.A(n_425),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_427),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_432),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_432),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_385),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_407),
.B(n_238),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_386),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_425),
.Y(n_583)
);

OAI21xp33_ASAP7_75t_SL g584 ( 
.A1(n_429),
.A2(n_379),
.B(n_377),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_429),
.B(n_190),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_386),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_386),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_420),
.B(n_193),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_433),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_412),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_433),
.B(n_164),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_425),
.B(n_209),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_435),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_435),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_530),
.Y(n_595)
);

A2O1A1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_584),
.A2(n_441),
.B(n_379),
.C(n_377),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_449),
.B(n_477),
.Y(n_597)
);

O2A1O1Ixp33_ASAP7_75t_L g598 ( 
.A1(n_584),
.A2(n_368),
.B(n_438),
.C(n_373),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_515),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_530),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_449),
.B(n_425),
.Y(n_601)
);

NAND2xp33_ASAP7_75t_L g602 ( 
.A(n_531),
.B(n_244),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_477),
.B(n_531),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_585),
.A2(n_525),
.B1(n_462),
.B2(n_452),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_590),
.B(n_425),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_527),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_486),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_535),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_451),
.B(n_430),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_515),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_509),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_535),
.Y(n_612)
);

INVxp33_ASAP7_75t_L g613 ( 
.A(n_523),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_590),
.B(n_430),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_483),
.B(n_430),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_526),
.B(n_430),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_536),
.B(n_194),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_452),
.B(n_430),
.Y(n_618)
);

NAND2xp33_ASAP7_75t_L g619 ( 
.A(n_529),
.B(n_534),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_527),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_466),
.B(n_164),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_459),
.B(n_484),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_539),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_495),
.B(n_430),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_471),
.B(n_167),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_537),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_537),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_459),
.B(n_430),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_496),
.B(n_430),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_529),
.B(n_244),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_546),
.Y(n_631)
);

NOR3xp33_ASAP7_75t_L g632 ( 
.A(n_571),
.B(n_353),
.C(n_375),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_448),
.B(n_355),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_585),
.A2(n_226),
.B1(n_291),
.B2(n_285),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_497),
.B(n_438),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_546),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_542),
.B(n_388),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_550),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_509),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_562),
.B(n_388),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_550),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_541),
.Y(n_642)
);

O2A1O1Ixp5_ASAP7_75t_L g643 ( 
.A1(n_585),
.A2(n_220),
.B(n_206),
.C(n_284),
.Y(n_643)
);

NOR2xp67_ASAP7_75t_L g644 ( 
.A(n_534),
.B(n_247),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_541),
.Y(n_645)
);

NAND2x1p5_ASAP7_75t_L g646 ( 
.A(n_453),
.B(n_208),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_502),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_502),
.B(n_355),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_564),
.A2(n_267),
.B1(n_261),
.B2(n_257),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_509),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_543),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_470),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_585),
.A2(n_246),
.B1(n_263),
.B2(n_260),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_553),
.Y(n_654)
);

INVxp67_ASAP7_75t_SL g655 ( 
.A(n_485),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_543),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_481),
.B(n_553),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_481),
.B(n_388),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_574),
.B(n_167),
.Y(n_659)
);

O2A1O1Ixp33_ASAP7_75t_L g660 ( 
.A1(n_540),
.A2(n_367),
.B(n_357),
.C(n_359),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_462),
.B(n_224),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_540),
.B(n_228),
.Y(n_662)
);

A2O1A1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_563),
.A2(n_366),
.B(n_375),
.C(n_373),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_556),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_556),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_545),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_557),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_557),
.B(n_388),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_548),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_548),
.B(n_229),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_552),
.B(n_251),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_492),
.B(n_169),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_558),
.B(n_393),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_558),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_SL g675 ( 
.A(n_528),
.B(n_209),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_511),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_511),
.A2(n_209),
.B1(n_398),
.B2(n_393),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_511),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_476),
.B(n_272),
.C(n_188),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_552),
.B(n_252),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_561),
.B(n_393),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_554),
.B(n_254),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_554),
.Y(n_683)
);

O2A1O1Ixp5_ASAP7_75t_L g684 ( 
.A1(n_561),
.A2(n_399),
.B(n_398),
.C(n_357),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_559),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_572),
.B(n_398),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_539),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_559),
.B(n_256),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_568),
.Y(n_689)
);

O2A1O1Ixp5_ASAP7_75t_L g690 ( 
.A1(n_572),
.A2(n_399),
.B(n_367),
.C(n_366),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_568),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_577),
.B(n_399),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_569),
.B(n_258),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_577),
.B(n_386),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_569),
.B(n_269),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_458),
.B(n_169),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_547),
.A2(n_277),
.B1(n_274),
.B2(n_180),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_458),
.B(n_172),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_578),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_578),
.B(n_579),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_579),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_570),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_589),
.B(n_386),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_520),
.B(n_359),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_457),
.B(n_172),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_511),
.B(n_179),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_511),
.A2(n_177),
.B1(n_178),
.B2(n_233),
.Y(n_707)
);

NAND2x1_ASAP7_75t_L g708 ( 
.A(n_539),
.B(n_386),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_589),
.B(n_386),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_593),
.B(n_386),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_593),
.B(n_389),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_547),
.A2(n_293),
.B1(n_180),
.B2(n_283),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_570),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_594),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_575),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_594),
.B(n_389),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_532),
.B(n_283),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_575),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_519),
.B(n_286),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_591),
.B(n_389),
.Y(n_720)
);

OAI22xp33_ASAP7_75t_SL g721 ( 
.A1(n_588),
.A2(n_551),
.B1(n_560),
.B2(n_468),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_555),
.B(n_566),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_519),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_567),
.B(n_389),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_573),
.B(n_360),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_522),
.B(n_286),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_581),
.B(n_389),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_532),
.B(n_507),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_536),
.B(n_360),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_460),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_464),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_464),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_532),
.A2(n_178),
.B1(n_233),
.B2(n_297),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_465),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_522),
.B(n_290),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_454),
.B(n_455),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_532),
.A2(n_297),
.B1(n_299),
.B2(n_307),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_465),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_469),
.Y(n_739)
);

NAND2x1p5_ASAP7_75t_L g740 ( 
.A(n_453),
.B(n_389),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_454),
.B(n_389),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_447),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_454),
.B(n_455),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_469),
.B(n_290),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_447),
.Y(n_745)
);

A2O1A1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_563),
.A2(n_299),
.B(n_347),
.C(n_348),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_450),
.Y(n_747)
);

NOR3xp33_ASAP7_75t_L g748 ( 
.A(n_544),
.B(n_204),
.C(n_198),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_450),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_478),
.B(n_292),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_455),
.B(n_389),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_536),
.B(n_347),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_478),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_479),
.B(n_292),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_468),
.B(n_304),
.Y(n_755)
);

NOR2x1p5_ASAP7_75t_L g756 ( 
.A(n_494),
.B(n_215),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_479),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_480),
.B(n_293),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_480),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_472),
.B(n_491),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_487),
.Y(n_761)
);

O2A1O1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_592),
.A2(n_348),
.B(n_304),
.C(n_300),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_487),
.B(n_300),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_547),
.A2(n_270),
.B1(n_245),
.B2(n_282),
.Y(n_764)
);

OAI21xp33_ASAP7_75t_SL g765 ( 
.A1(n_604),
.A2(n_597),
.B(n_603),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_721),
.B(n_474),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_647),
.Y(n_767)
);

NOR2x2_ASAP7_75t_L g768 ( 
.A(n_755),
.B(n_498),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_674),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_599),
.B(n_536),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_674),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_614),
.B(n_488),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_610),
.B(n_536),
.Y(n_773)
);

INVx5_ASAP7_75t_L g774 ( 
.A(n_623),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_606),
.Y(n_775)
);

INVx4_ASAP7_75t_L g776 ( 
.A(n_611),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_606),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_607),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_621),
.B(n_488),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_R g780 ( 
.A(n_607),
.B(n_490),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_620),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_659),
.A2(n_505),
.B1(n_533),
.B2(n_565),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_648),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_613),
.A2(n_539),
.B1(n_506),
.B2(n_474),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_625),
.B(n_510),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_620),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_633),
.B(n_490),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_729),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_657),
.B(n_510),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_725),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_642),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_642),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_613),
.B(n_514),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_696),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_662),
.A2(n_602),
.B1(n_609),
.B2(n_661),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_652),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_645),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_662),
.A2(n_494),
.B1(n_503),
.B2(n_512),
.Y(n_798)
);

AOI21xp33_ASAP7_75t_L g799 ( 
.A1(n_672),
.A2(n_506),
.B(n_249),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_631),
.B(n_514),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_636),
.B(n_518),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_729),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_638),
.B(n_518),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_597),
.B(n_605),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_729),
.B(n_583),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_641),
.B(n_524),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_722),
.B(n_623),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_645),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_698),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_602),
.A2(n_524),
.B1(n_482),
.B2(n_513),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_611),
.Y(n_811)
);

AND2x4_ASAP7_75t_SL g812 ( 
.A(n_611),
.B(n_485),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_623),
.B(n_485),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_611),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_651),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_654),
.B(n_456),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_651),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_656),
.Y(n_818)
);

OR2x6_ASAP7_75t_L g819 ( 
.A(n_676),
.B(n_549),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_687),
.B(n_485),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_639),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_678),
.B(n_583),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_664),
.B(n_456),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_656),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_669),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_661),
.A2(n_516),
.B1(n_489),
.B2(n_475),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_649),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_605),
.B(n_583),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_669),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_665),
.B(n_461),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_704),
.A2(n_489),
.B1(n_461),
.B2(n_463),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_687),
.B(n_728),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_752),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_639),
.A2(n_587),
.B1(n_586),
.B2(n_472),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_683),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_683),
.Y(n_836)
);

INVx5_ASAP7_75t_L g837 ( 
.A(n_687),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_706),
.A2(n_500),
.B1(n_508),
.B2(n_491),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_R g839 ( 
.A(n_619),
.B(n_549),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_667),
.B(n_500),
.Y(n_840)
);

INVx4_ASAP7_75t_L g841 ( 
.A(n_639),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_699),
.B(n_701),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_685),
.Y(n_843)
);

INVx6_ASAP7_75t_L g844 ( 
.A(n_752),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_685),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_714),
.B(n_463),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_689),
.Y(n_847)
);

NOR2x2_ASAP7_75t_L g848 ( 
.A(n_675),
.B(n_218),
.Y(n_848)
);

AND2x6_ASAP7_75t_L g849 ( 
.A(n_650),
.B(n_467),
.Y(n_849)
);

AND2x2_ASAP7_75t_SL g850 ( 
.A(n_619),
.B(n_500),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_689),
.A2(n_516),
.B1(n_499),
.B2(n_475),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_691),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_650),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_752),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_635),
.B(n_467),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_700),
.B(n_473),
.Y(n_856)
);

BUFx8_ASAP7_75t_L g857 ( 
.A(n_666),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_691),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_702),
.Y(n_859)
);

BUFx4f_ASAP7_75t_L g860 ( 
.A(n_646),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_702),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_622),
.B(n_650),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_713),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_756),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_705),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_744),
.B(n_500),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_SL g867 ( 
.A1(n_707),
.A2(n_259),
.B1(n_264),
.B2(n_268),
.Y(n_867)
);

AND2x6_ASAP7_75t_SL g868 ( 
.A(n_717),
.B(n_271),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_713),
.A2(n_715),
.B1(n_608),
.B2(n_595),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_715),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_744),
.B(n_508),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_723),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_750),
.B(n_508),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_655),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_616),
.B(n_485),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_600),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_612),
.A2(n_501),
.B1(n_473),
.B2(n_482),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_601),
.B(n_582),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_626),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_627),
.A2(n_504),
.B1(n_499),
.B2(n_501),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_658),
.B(n_513),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_724),
.A2(n_580),
.B(n_582),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_718),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_617),
.B(n_587),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_617),
.B(n_587),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_750),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_723),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_596),
.B(n_504),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_596),
.B(n_517),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_646),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_730),
.B(n_517),
.Y(n_891)
);

AO22x1_ASAP7_75t_L g892 ( 
.A1(n_748),
.A2(n_276),
.B1(n_275),
.B2(n_521),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_617),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_731),
.A2(n_521),
.B1(n_472),
.B2(n_538),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_742),
.Y(n_895)
);

NOR2x1p5_ASAP7_75t_L g896 ( 
.A(n_679),
.B(n_586),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_745),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_732),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_734),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_738),
.B(n_521),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_754),
.B(n_538),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_745),
.Y(n_902)
);

AND2x6_ASAP7_75t_L g903 ( 
.A(n_629),
.B(n_538),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_747),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_739),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_618),
.B(n_582),
.Y(n_906)
);

NAND2xp33_ASAP7_75t_L g907 ( 
.A(n_740),
.B(n_582),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_753),
.B(n_582),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_757),
.B(n_580),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_632),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_749),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_759),
.Y(n_912)
);

NAND2xp33_ASAP7_75t_SL g913 ( 
.A(n_733),
.B(n_580),
.Y(n_913)
);

CKINVDCx6p67_ASAP7_75t_R g914 ( 
.A(n_680),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_749),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_761),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_754),
.B(n_758),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_680),
.A2(n_580),
.B1(n_576),
.B2(n_493),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_668),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_758),
.B(n_580),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_737),
.B(n_1),
.Y(n_921)
);

O2A1O1Ixp5_ASAP7_75t_L g922 ( 
.A1(n_615),
.A2(n_576),
.B(n_493),
.C(n_151),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_694),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_703),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_682),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_763),
.B(n_719),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_764),
.B(n_88),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_634),
.A2(n_394),
.B1(n_391),
.B2(n_576),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_763),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_637),
.B(n_576),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_712),
.B(n_719),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_628),
.B(n_576),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_682),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_709),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_740),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_726),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_710),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_653),
.A2(n_394),
.B1(n_391),
.B2(n_576),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_711),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_720),
.B(n_615),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_716),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_624),
.B(n_493),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_673),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_708),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_726),
.B(n_84),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_681),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_697),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_735),
.B(n_3),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_735),
.B(n_3),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_SL g950 ( 
.A(n_778),
.B(n_644),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_774),
.A2(n_837),
.B(n_807),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_876),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_865),
.B(n_677),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_795),
.A2(n_782),
.B1(n_804),
.B2(n_785),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_794),
.B(n_688),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_882),
.A2(n_741),
.B(n_751),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_776),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_833),
.B(n_688),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_SL g959 ( 
.A1(n_947),
.A2(n_760),
.B1(n_743),
.B2(n_736),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_767),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_795),
.A2(n_640),
.B1(n_624),
.B2(n_727),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_778),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_879),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_765),
.A2(n_692),
.B(n_686),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_804),
.A2(n_695),
.B1(n_693),
.B2(n_746),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_917),
.A2(n_762),
.B(n_660),
.C(n_695),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_779),
.A2(n_693),
.B1(n_746),
.B2(n_663),
.Y(n_967)
);

AND2x2_ASAP7_75t_SL g968 ( 
.A(n_927),
.B(n_860),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_809),
.B(n_598),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_827),
.A2(n_663),
.B1(n_671),
.B2(n_670),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_796),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_917),
.A2(n_926),
.B1(n_927),
.B2(n_931),
.Y(n_972)
);

NAND2x1p5_ASAP7_75t_L g973 ( 
.A(n_774),
.B(n_670),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_774),
.A2(n_630),
.B(n_671),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_837),
.A2(n_643),
.B(n_684),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_833),
.B(n_78),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_837),
.A2(n_807),
.B(n_862),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_943),
.B(n_493),
.Y(n_978)
);

AOI22x1_ASAP7_75t_L g979 ( 
.A1(n_896),
.A2(n_690),
.B1(n_394),
.B2(n_391),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_828),
.A2(n_493),
.B(n_99),
.Y(n_980)
);

NOR3xp33_ASAP7_75t_L g981 ( 
.A(n_787),
.B(n_4),
.C(n_5),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_926),
.A2(n_394),
.B(n_391),
.C(n_11),
.Y(n_982)
);

NOR2xp67_ASAP7_75t_L g983 ( 
.A(n_790),
.B(n_148),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_946),
.B(n_919),
.Y(n_984)
);

INVx5_ASAP7_75t_L g985 ( 
.A(n_935),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_783),
.B(n_886),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_936),
.B(n_6),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_814),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_789),
.B(n_394),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_837),
.A2(n_394),
.B(n_391),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_899),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_R g992 ( 
.A(n_913),
.B(n_147),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_940),
.A2(n_391),
.B(n_394),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_915),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_940),
.A2(n_391),
.B(n_394),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_802),
.A2(n_391),
.B1(n_129),
.B2(n_122),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_923),
.B(n_113),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_929),
.A2(n_8),
.B(n_11),
.C(n_12),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_925),
.A2(n_933),
.B(n_828),
.C(n_873),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_910),
.A2(n_8),
.B(n_13),
.C(n_15),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_924),
.B(n_91),
.Y(n_1001)
);

INVxp67_ASAP7_75t_SL g1002 ( 
.A(n_814),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_788),
.Y(n_1003)
);

CKINVDCx11_ASAP7_75t_R g1004 ( 
.A(n_868),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_866),
.A2(n_18),
.B(n_22),
.C(n_23),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_788),
.B(n_18),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_915),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_866),
.A2(n_25),
.B(n_26),
.C(n_28),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_860),
.B(n_77),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_844),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_844),
.A2(n_76),
.B1(n_73),
.B2(n_69),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_805),
.Y(n_1012)
);

HAxp5_ASAP7_75t_L g1013 ( 
.A(n_768),
.B(n_25),
.CON(n_1013),
.SN(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_844),
.A2(n_68),
.B1(n_66),
.B2(n_65),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_793),
.B(n_26),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_SL g1016 ( 
.A(n_890),
.B(n_28),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_872),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_934),
.B(n_31),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_780),
.Y(n_1019)
);

NAND2x1p5_ASAP7_75t_L g1020 ( 
.A(n_776),
.B(n_35),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_937),
.B(n_35),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_864),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_871),
.A2(n_37),
.B(n_39),
.C(n_41),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_905),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_769),
.B(n_44),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_893),
.B(n_45),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_914),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_907),
.A2(n_49),
.B(n_50),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_854),
.A2(n_50),
.B1(n_832),
.B2(n_871),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_941),
.B(n_855),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_772),
.B(n_842),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_856),
.B(n_939),
.Y(n_1032)
);

O2A1O1Ixp5_ASAP7_75t_L g1033 ( 
.A1(n_766),
.A2(n_799),
.B(n_832),
.C(n_922),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_805),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_887),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_939),
.B(n_912),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_854),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_935),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_916),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_857),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_775),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_777),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_945),
.A2(n_770),
.B1(n_773),
.B2(n_771),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_781),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_780),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_841),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_873),
.A2(n_901),
.B(n_945),
.C(n_840),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_R g1048 ( 
.A(n_811),
.B(n_890),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_791),
.B(n_817),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_898),
.B(n_921),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_875),
.A2(n_881),
.B(n_841),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_792),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_770),
.A2(n_773),
.B1(n_884),
.B2(n_885),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_887),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_848),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_935),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_949),
.A2(n_766),
.B(n_948),
.C(n_883),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_898),
.B(n_867),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_798),
.B(n_884),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_R g1060 ( 
.A(n_811),
.B(n_857),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_875),
.A2(n_853),
.B(n_930),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_885),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_791),
.B(n_817),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_798),
.B(n_892),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_840),
.A2(n_853),
.B1(n_869),
.B2(n_874),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_822),
.A2(n_901),
.B1(n_819),
.B2(n_797),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_850),
.A2(n_878),
.B(n_888),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_821),
.B(n_822),
.Y(n_1068)
);

INVxp67_ASAP7_75t_L g1069 ( 
.A(n_920),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_819),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_800),
.A2(n_806),
.B(n_803),
.C(n_801),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_935),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_812),
.A2(n_820),
.B(n_813),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_869),
.A2(n_850),
.B1(n_894),
.B2(n_821),
.Y(n_1074)
);

NAND2x1p5_ASAP7_75t_L g1075 ( 
.A(n_897),
.B(n_904),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_889),
.A2(n_846),
.B(n_830),
.C(n_823),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_816),
.A2(n_784),
.B(n_891),
.C(n_942),
.Y(n_1077)
);

AO21x1_ASAP7_75t_L g1078 ( 
.A1(n_942),
.A2(n_932),
.B(n_878),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_834),
.A2(n_906),
.B(n_900),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_897),
.B(n_911),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_904),
.B(n_911),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_824),
.B(n_870),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_812),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_808),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_815),
.A2(n_852),
.B(n_835),
.C(n_836),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_906),
.A2(n_820),
.B(n_813),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_819),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_786),
.B(n_861),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_824),
.B(n_829),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_858),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_972),
.B(n_863),
.Y(n_1091)
);

BUFx12f_ASAP7_75t_L g1092 ( 
.A(n_1004),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_993),
.A2(n_932),
.B(n_909),
.Y(n_1093)
);

O2A1O1Ixp5_ASAP7_75t_L g1094 ( 
.A1(n_980),
.A2(n_944),
.B(n_908),
.C(n_825),
.Y(n_1094)
);

NOR2x1_ASAP7_75t_L g1095 ( 
.A(n_962),
.B(n_859),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1031),
.B(n_829),
.Y(n_1096)
);

AO21x2_ASAP7_75t_L g1097 ( 
.A1(n_964),
.A2(n_839),
.B(n_838),
.Y(n_1097)
);

NOR2xp67_ASAP7_75t_L g1098 ( 
.A(n_1022),
.B(n_818),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_952),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1031),
.B(n_870),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_971),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_968),
.B(n_839),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_960),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_955),
.B(n_847),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_1012),
.B(n_843),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1013),
.B(n_845),
.Y(n_1106)
);

AOI31xp67_ASAP7_75t_L g1107 ( 
.A1(n_969),
.A2(n_902),
.A3(n_895),
.B(n_918),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_984),
.B(n_831),
.Y(n_1108)
);

INVx3_ASAP7_75t_SL g1109 ( 
.A(n_1040),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1019),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_SL g1111 ( 
.A1(n_1047),
.A2(n_849),
.B(n_903),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_1078),
.A2(n_903),
.A3(n_849),
.B(n_810),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_984),
.B(n_1030),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_993),
.A2(n_810),
.B(n_877),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1030),
.B(n_831),
.Y(n_1115)
);

AOI211x1_ASAP7_75t_L g1116 ( 
.A1(n_953),
.A2(n_894),
.B(n_880),
.C(n_877),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_995),
.A2(n_880),
.B(n_826),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1050),
.B(n_903),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_963),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_954),
.B(n_903),
.Y(n_1120)
);

AO31x2_ASAP7_75t_L g1121 ( 
.A1(n_965),
.A2(n_1067),
.A3(n_967),
.B(n_966),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1071),
.A2(n_928),
.B(n_938),
.Y(n_1122)
);

O2A1O1Ixp5_ASAP7_75t_L g1123 ( 
.A1(n_1033),
.A2(n_903),
.B(n_849),
.C(n_826),
.Y(n_1123)
);

OAI21xp33_ASAP7_75t_L g1124 ( 
.A1(n_1016),
.A2(n_851),
.B(n_928),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_951),
.A2(n_938),
.B(n_851),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_1045),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1058),
.A2(n_849),
.B1(n_1055),
.B2(n_959),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_986),
.B(n_849),
.Y(n_1128)
);

BUFx10_ASAP7_75t_L g1129 ( 
.A(n_1025),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_995),
.A2(n_956),
.B(n_951),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1032),
.B(n_1015),
.Y(n_1131)
);

AOI211x1_ASAP7_75t_L g1132 ( 
.A1(n_991),
.A2(n_1039),
.B(n_1024),
.C(n_1021),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1032),
.B(n_1036),
.Y(n_1133)
);

INVx4_ASAP7_75t_L g1134 ( 
.A(n_985),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_977),
.A2(n_1076),
.B(n_1065),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1012),
.B(n_1034),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1067),
.A2(n_999),
.B(n_1051),
.Y(n_1137)
);

AO31x2_ASAP7_75t_L g1138 ( 
.A1(n_1061),
.A2(n_1074),
.A3(n_982),
.B(n_1029),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_977),
.A2(n_974),
.B(n_1051),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1041),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1042),
.Y(n_1141)
);

OA21x2_ASAP7_75t_L g1142 ( 
.A1(n_1079),
.A2(n_1061),
.B(n_1086),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_974),
.A2(n_1077),
.B(n_1073),
.Y(n_1143)
);

BUFx12f_ASAP7_75t_L g1144 ( 
.A(n_1010),
.Y(n_1144)
);

AOI211x1_ASAP7_75t_L g1145 ( 
.A1(n_1018),
.A2(n_1021),
.B(n_1036),
.C(n_1028),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_950),
.B(n_1043),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_987),
.B(n_1026),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_1060),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1003),
.B(n_1037),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1062),
.B(n_1090),
.Y(n_1150)
);

AOI221x1_ASAP7_75t_L g1151 ( 
.A1(n_1005),
.A2(n_1023),
.B1(n_1008),
.B2(n_981),
.C(n_1064),
.Y(n_1151)
);

NOR4xp25_ASAP7_75t_L g1152 ( 
.A(n_1000),
.B(n_998),
.C(n_1057),
.D(n_970),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1059),
.B(n_1069),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1086),
.A2(n_989),
.B(n_975),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1018),
.A2(n_1009),
.B(n_1001),
.C(n_997),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1088),
.B(n_1063),
.Y(n_1156)
);

OAI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1027),
.A2(n_1053),
.B1(n_996),
.B2(n_983),
.Y(n_1157)
);

CKINVDCx8_ASAP7_75t_R g1158 ( 
.A(n_988),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1049),
.B(n_1063),
.Y(n_1159)
);

AO32x2_ASAP7_75t_L g1160 ( 
.A1(n_1011),
.A2(n_1014),
.A3(n_1066),
.B1(n_979),
.B2(n_1087),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_988),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_988),
.Y(n_1162)
);

BUFx10_ASAP7_75t_L g1163 ( 
.A(n_976),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_994),
.Y(n_1164)
);

O2A1O1Ixp5_ASAP7_75t_SL g1165 ( 
.A1(n_1044),
.A2(n_1052),
.B(n_1084),
.C(n_1082),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_985),
.A2(n_1001),
.B1(n_997),
.B2(n_976),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1007),
.Y(n_1167)
);

AO31x2_ASAP7_75t_L g1168 ( 
.A1(n_1070),
.A2(n_978),
.A3(n_1049),
.B(n_1017),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1068),
.B(n_1035),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_990),
.A2(n_1085),
.B(n_1089),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1034),
.B(n_1010),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_1048),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_990),
.A2(n_978),
.B(n_973),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1054),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1080),
.A2(n_1081),
.B(n_958),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_973),
.A2(n_1046),
.B(n_1075),
.Y(n_1176)
);

AO21x2_ASAP7_75t_L g1177 ( 
.A1(n_992),
.A2(n_958),
.B(n_1002),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1010),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1046),
.A2(n_1075),
.B(n_957),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1006),
.B(n_1034),
.Y(n_1180)
);

AOI21xp33_ASAP7_75t_L g1181 ( 
.A1(n_1020),
.A2(n_1038),
.B(n_1056),
.Y(n_1181)
);

OR2x6_ASAP7_75t_SL g1182 ( 
.A(n_1020),
.B(n_985),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_957),
.A2(n_985),
.B(n_1083),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_1038),
.A2(n_1056),
.A3(n_1072),
.B(n_1078),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1072),
.B(n_1038),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1056),
.B(n_1072),
.Y(n_1186)
);

INVx5_ASAP7_75t_L g1187 ( 
.A(n_985),
.Y(n_1187)
);

AO21x1_ASAP7_75t_L g1188 ( 
.A1(n_954),
.A2(n_965),
.B(n_980),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_961),
.A2(n_837),
.B(n_774),
.Y(n_1189)
);

BUFx12f_ASAP7_75t_L g1190 ( 
.A(n_1004),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_993),
.A2(n_995),
.B(n_956),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_962),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_962),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_962),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1031),
.B(n_984),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_972),
.B(n_613),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_993),
.A2(n_995),
.B(n_956),
.Y(n_1197)
);

AOI211x1_ASAP7_75t_L g1198 ( 
.A1(n_969),
.A2(n_953),
.B(n_984),
.C(n_571),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_993),
.A2(n_995),
.B(n_956),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_960),
.B(n_787),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1031),
.B(n_984),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1031),
.B(n_984),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_993),
.A2(n_995),
.B(n_956),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_962),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1047),
.A2(n_1067),
.B(n_954),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_961),
.A2(n_837),
.B(n_774),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_SL g1207 ( 
.A1(n_972),
.A2(n_498),
.B(n_755),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_993),
.A2(n_995),
.B(n_956),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1031),
.B(n_984),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1031),
.B(n_984),
.Y(n_1210)
);

AO21x2_ASAP7_75t_L g1211 ( 
.A1(n_980),
.A2(n_964),
.B(n_1047),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_960),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1078),
.A2(n_961),
.A3(n_1047),
.B(n_954),
.Y(n_1213)
);

NOR4xp25_ASAP7_75t_L g1214 ( 
.A(n_1000),
.B(n_1008),
.C(n_1023),
.D(n_1005),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1031),
.B(n_984),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_968),
.A2(n_827),
.B1(n_312),
.B2(n_328),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1038),
.Y(n_1217)
);

O2A1O1Ixp5_ASAP7_75t_SL g1218 ( 
.A1(n_965),
.A2(n_766),
.B(n_662),
.C(n_954),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_972),
.A2(n_968),
.B1(n_984),
.B2(n_1031),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1013),
.B(n_783),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_968),
.A2(n_827),
.B1(n_312),
.B2(n_328),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_961),
.A2(n_837),
.B(n_774),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_972),
.A2(n_1047),
.B(n_917),
.C(n_926),
.Y(n_1223)
);

NAND3x1_ASAP7_75t_L g1224 ( 
.A(n_1027),
.B(n_468),
.C(n_755),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1038),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1038),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1047),
.A2(n_1067),
.B(n_954),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_972),
.A2(n_1047),
.B(n_917),
.C(n_926),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_961),
.A2(n_837),
.B(n_774),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1130),
.A2(n_1197),
.B(n_1191),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1199),
.A2(n_1208),
.B(n_1203),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1188),
.A2(n_1196),
.B1(n_1211),
.B2(n_1205),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_1187),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1099),
.Y(n_1234)
);

O2A1O1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1207),
.A2(n_1228),
.B(n_1223),
.C(n_1146),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1119),
.Y(n_1236)
);

CKINVDCx20_ASAP7_75t_R g1237 ( 
.A(n_1192),
.Y(n_1237)
);

AOI221xp5_ASAP7_75t_L g1238 ( 
.A1(n_1152),
.A2(n_1214),
.B1(n_1207),
.B2(n_1219),
.C(n_1157),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1224),
.A2(n_1221),
.B1(n_1216),
.B2(n_1219),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1143),
.A2(n_1154),
.B(n_1093),
.Y(n_1240)
);

AOI21xp33_ASAP7_75t_L g1241 ( 
.A1(n_1155),
.A2(n_1131),
.B(n_1104),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_SL g1242 ( 
.A(n_1158),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1173),
.A2(n_1170),
.B(n_1137),
.Y(n_1243)
);

AO21x2_ASAP7_75t_L g1244 ( 
.A1(n_1227),
.A2(n_1229),
.B(n_1222),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1195),
.B(n_1201),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1211),
.A2(n_1227),
.B1(n_1195),
.B2(n_1215),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_1101),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1189),
.A2(n_1206),
.B(n_1123),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1201),
.B(n_1202),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1187),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1147),
.B(n_1220),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1218),
.A2(n_1117),
.B(n_1114),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1202),
.A2(n_1215),
.B1(n_1210),
.B2(n_1209),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1140),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1200),
.B(n_1153),
.Y(n_1255)
);

BUFx4f_ASAP7_75t_SL g1256 ( 
.A(n_1144),
.Y(n_1256)
);

NAND2x1p5_ASAP7_75t_L g1257 ( 
.A(n_1134),
.B(n_1102),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1142),
.A2(n_1176),
.B(n_1111),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1142),
.A2(n_1094),
.B(n_1120),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1103),
.Y(n_1260)
);

AO21x2_ASAP7_75t_L g1261 ( 
.A1(n_1097),
.A2(n_1166),
.B(n_1122),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1152),
.A2(n_1091),
.B(n_1166),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1151),
.A2(n_1125),
.A3(n_1118),
.B(n_1096),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1165),
.A2(n_1179),
.B(n_1175),
.Y(n_1264)
);

AO21x2_ASAP7_75t_L g1265 ( 
.A1(n_1177),
.A2(n_1153),
.B(n_1214),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1141),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1209),
.B(n_1210),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1113),
.B(n_1212),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1167),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1113),
.A2(n_1115),
.B(n_1096),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1175),
.A2(n_1159),
.B(n_1183),
.Y(n_1271)
);

AO32x2_ASAP7_75t_L g1272 ( 
.A1(n_1198),
.A2(n_1121),
.A3(n_1213),
.B1(n_1145),
.B2(n_1138),
.Y(n_1272)
);

OAI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1127),
.A2(n_1133),
.B1(n_1108),
.B2(n_1100),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1149),
.B(n_1106),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1108),
.A2(n_1128),
.B(n_1169),
.Y(n_1275)
);

AO21x2_ASAP7_75t_L g1276 ( 
.A1(n_1177),
.A2(n_1181),
.B(n_1183),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1150),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1124),
.A2(n_1180),
.B(n_1156),
.C(n_1121),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1110),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1164),
.A2(n_1174),
.B(n_1095),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1134),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1107),
.A2(n_1225),
.B(n_1185),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1129),
.A2(n_1163),
.B1(n_1105),
.B2(n_1181),
.Y(n_1283)
);

NOR2x1_ASAP7_75t_SL g1284 ( 
.A(n_1217),
.B(n_1226),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1098),
.A2(n_1171),
.B(n_1162),
.Y(n_1285)
);

AND2x2_ASAP7_75t_SL g1286 ( 
.A(n_1121),
.B(n_1182),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1186),
.B(n_1225),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1132),
.A2(n_1126),
.B1(n_1116),
.B2(n_1172),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1112),
.A2(n_1213),
.B(n_1138),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1194),
.Y(n_1290)
);

OR2x2_ASAP7_75t_L g1291 ( 
.A(n_1161),
.B(n_1204),
.Y(n_1291)
);

NAND2x1p5_ASAP7_75t_L g1292 ( 
.A(n_1186),
.B(n_1178),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1112),
.A2(n_1184),
.B(n_1168),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1193),
.A2(n_1129),
.B(n_1160),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1184),
.A2(n_1160),
.B(n_1163),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1184),
.A2(n_1160),
.B(n_1217),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1217),
.A2(n_1226),
.B(n_1148),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_1109),
.Y(n_1298)
);

CKINVDCx6p67_ASAP7_75t_R g1299 ( 
.A(n_1092),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1226),
.Y(n_1300)
);

INVx4_ASAP7_75t_L g1301 ( 
.A(n_1190),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_SL g1302 ( 
.A(n_1192),
.B(n_607),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1147),
.B(n_1013),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1136),
.B(n_976),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1224),
.A2(n_312),
.B1(n_328),
.B2(n_317),
.Y(n_1305)
);

NAND3xp33_ASAP7_75t_L g1306 ( 
.A(n_1207),
.B(n_625),
.C(n_621),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1224),
.A2(n_312),
.B1(n_328),
.B2(n_317),
.Y(n_1307)
);

NOR2xp67_ASAP7_75t_L g1308 ( 
.A(n_1212),
.B(n_607),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1147),
.B(n_1013),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1130),
.A2(n_1197),
.B(n_1191),
.Y(n_1310)
);

NAND3xp33_ASAP7_75t_L g1311 ( 
.A(n_1207),
.B(n_625),
.C(n_621),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1130),
.A2(n_1197),
.B(n_1191),
.Y(n_1312)
);

AO32x2_ASAP7_75t_L g1313 ( 
.A1(n_1219),
.A2(n_954),
.A3(n_965),
.B1(n_1166),
.B2(n_1029),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1212),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1099),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1195),
.B(n_1201),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1130),
.A2(n_1197),
.B(n_1191),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1195),
.B(n_1201),
.Y(n_1318)
);

AO221x2_ASAP7_75t_L g1319 ( 
.A1(n_1207),
.A2(n_1205),
.B1(n_1227),
.B2(n_1219),
.C(n_954),
.Y(n_1319)
);

OR2x6_ASAP7_75t_L g1320 ( 
.A(n_1111),
.B(n_1198),
.Y(n_1320)
);

AOI21xp33_ASAP7_75t_L g1321 ( 
.A1(n_1207),
.A2(n_659),
.B(n_613),
.Y(n_1321)
);

INVxp67_ASAP7_75t_L g1322 ( 
.A(n_1212),
.Y(n_1322)
);

INVx6_ASAP7_75t_L g1323 ( 
.A(n_1187),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1099),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1212),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1130),
.A2(n_1197),
.B(n_1191),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1187),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1195),
.B(n_1201),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1195),
.B(n_1201),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_SL g1330 ( 
.A1(n_1155),
.A2(n_1057),
.B(n_1219),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1130),
.A2(n_1197),
.B(n_1191),
.Y(n_1331)
);

CKINVDCx8_ASAP7_75t_R g1332 ( 
.A(n_1192),
.Y(n_1332)
);

NOR4xp25_ASAP7_75t_L g1333 ( 
.A(n_1224),
.B(n_1207),
.C(n_1000),
.D(n_1008),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1099),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1195),
.A2(n_972),
.B1(n_968),
.B2(n_1201),
.Y(n_1335)
);

A2O1A1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1122),
.A2(n_972),
.B(n_1124),
.C(n_1047),
.Y(n_1336)
);

AO21x2_ASAP7_75t_L g1337 ( 
.A1(n_1143),
.A2(n_1139),
.B(n_1135),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1158),
.Y(n_1338)
);

BUFx4f_ASAP7_75t_L g1339 ( 
.A(n_1144),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1195),
.B(n_1201),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1101),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1212),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1195),
.B(n_1201),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1147),
.B(n_1013),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1195),
.B(n_1201),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1099),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1187),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1147),
.B(n_1013),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1130),
.A2(n_1197),
.B(n_1191),
.Y(n_1349)
);

BUFx10_ASAP7_75t_L g1350 ( 
.A(n_1192),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1340),
.B(n_1343),
.Y(n_1351)
);

NOR2xp67_ASAP7_75t_L g1352 ( 
.A(n_1255),
.B(n_1322),
.Y(n_1352)
);

NOR2x1_ASAP7_75t_SL g1353 ( 
.A(n_1276),
.B(n_1320),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1268),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1350),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1306),
.A2(n_1311),
.B(n_1239),
.C(n_1235),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1251),
.B(n_1303),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1253),
.A2(n_1345),
.B1(n_1318),
.B2(n_1267),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1253),
.B(n_1249),
.Y(n_1359)
);

AND2x6_ASAP7_75t_L g1360 ( 
.A(n_1250),
.B(n_1327),
.Y(n_1360)
);

AOI221xp5_ASAP7_75t_L g1361 ( 
.A1(n_1321),
.A2(n_1333),
.B1(n_1238),
.B2(n_1241),
.C(n_1262),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1259),
.A2(n_1248),
.B(n_1243),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1316),
.B(n_1328),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1234),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1329),
.B(n_1245),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1274),
.B(n_1319),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1245),
.B(n_1277),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1319),
.B(n_1314),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1325),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1270),
.B(n_1275),
.Y(n_1370)
);

OA21x2_ASAP7_75t_L g1371 ( 
.A1(n_1259),
.A2(n_1248),
.B(n_1243),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1336),
.A2(n_1330),
.B(n_1288),
.C(n_1294),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1319),
.B(n_1342),
.Y(n_1373)
);

AOI221x1_ASAP7_75t_SL g1374 ( 
.A1(n_1273),
.A2(n_1335),
.B1(n_1308),
.B2(n_1324),
.C(n_1254),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1278),
.B(n_1247),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_SL g1376 ( 
.A1(n_1232),
.A2(n_1285),
.B(n_1283),
.C(n_1281),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1246),
.B(n_1273),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1336),
.A2(n_1246),
.B1(n_1232),
.B2(n_1286),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1309),
.B(n_1344),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1278),
.B(n_1341),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1260),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1236),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_SL g1383 ( 
.A1(n_1250),
.A2(n_1327),
.B(n_1304),
.Y(n_1383)
);

OA22x2_ASAP7_75t_L g1384 ( 
.A1(n_1305),
.A2(n_1307),
.B1(n_1320),
.B2(n_1266),
.Y(n_1384)
);

NOR2xp67_ASAP7_75t_L g1385 ( 
.A(n_1291),
.B(n_1269),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1315),
.B(n_1334),
.Y(n_1386)
);

NAND2x1p5_ASAP7_75t_L g1387 ( 
.A(n_1271),
.B(n_1250),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_SL g1388 ( 
.A1(n_1250),
.A2(n_1327),
.B(n_1304),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1237),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1327),
.A2(n_1347),
.B(n_1233),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1286),
.A2(n_1242),
.B1(n_1346),
.B2(n_1283),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1271),
.A2(n_1339),
.B(n_1295),
.C(n_1264),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_SL g1393 ( 
.A1(n_1237),
.A2(n_1332),
.B1(n_1301),
.B2(n_1338),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1287),
.B(n_1300),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1265),
.B(n_1263),
.Y(n_1395)
);

NOR2x1_ASAP7_75t_SL g1396 ( 
.A(n_1276),
.B(n_1320),
.Y(n_1396)
);

O2A1O1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1257),
.A2(n_1320),
.B(n_1302),
.C(n_1261),
.Y(n_1397)
);

OA22x2_ASAP7_75t_L g1398 ( 
.A1(n_1297),
.A2(n_1296),
.B1(n_1295),
.B2(n_1233),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1265),
.Y(n_1399)
);

OA21x2_ASAP7_75t_L g1400 ( 
.A1(n_1252),
.A2(n_1293),
.B(n_1264),
.Y(n_1400)
);

O2A1O1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1257),
.A2(n_1298),
.B(n_1290),
.C(n_1244),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1292),
.B(n_1297),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1292),
.B(n_1279),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_SL g1404 ( 
.A1(n_1347),
.A2(n_1284),
.B(n_1337),
.Y(n_1404)
);

O2A1O1Ixp5_ASAP7_75t_L g1405 ( 
.A1(n_1339),
.A2(n_1313),
.B(n_1301),
.C(n_1272),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1332),
.A2(n_1323),
.B1(n_1256),
.B2(n_1313),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1280),
.B(n_1350),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1280),
.B(n_1272),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1256),
.B(n_1299),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1323),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1282),
.B(n_1296),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_SL g1412 ( 
.A1(n_1323),
.A2(n_1282),
.B(n_1258),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1289),
.B(n_1252),
.Y(n_1413)
);

BUFx8_ASAP7_75t_SL g1414 ( 
.A(n_1289),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1258),
.B(n_1240),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1230),
.B(n_1310),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1312),
.A2(n_1317),
.B(n_1326),
.C(n_1331),
.Y(n_1417)
);

OA22x2_ASAP7_75t_L g1418 ( 
.A1(n_1331),
.A2(n_1231),
.B1(n_1349),
.B2(n_1239),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1349),
.Y(n_1419)
);

A2O1A1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1306),
.A2(n_1311),
.B(n_1239),
.C(n_1235),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1350),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1321),
.A2(n_721),
.B(n_1207),
.C(n_1306),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1260),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1253),
.A2(n_1224),
.B1(n_968),
.B2(n_972),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1251),
.B(n_1348),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1253),
.A2(n_1224),
.B1(n_968),
.B2(n_972),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1251),
.B(n_1348),
.Y(n_1427)
);

A2O1A1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1306),
.A2(n_1311),
.B(n_1239),
.C(n_1235),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1251),
.B(n_1348),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1411),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1399),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1353),
.B(n_1396),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1364),
.Y(n_1433)
);

OAI211xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1361),
.A2(n_1420),
.B(n_1428),
.C(n_1356),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1366),
.B(n_1351),
.Y(n_1435)
);

INVx4_ASAP7_75t_L g1436 ( 
.A(n_1360),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1418),
.A2(n_1371),
.B(n_1362),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1419),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1387),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1398),
.Y(n_1440)
);

INVxp67_ASAP7_75t_R g1441 ( 
.A(n_1393),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1370),
.B(n_1358),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1402),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1398),
.Y(n_1444)
);

OR2x6_ASAP7_75t_L g1445 ( 
.A(n_1412),
.B(n_1397),
.Y(n_1445)
);

OR2x6_ASAP7_75t_L g1446 ( 
.A(n_1387),
.B(n_1378),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1414),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1370),
.A2(n_1378),
.B(n_1404),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1418),
.A2(n_1371),
.B(n_1362),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1369),
.Y(n_1450)
);

OR2x6_ASAP7_75t_L g1451 ( 
.A(n_1401),
.B(n_1407),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1358),
.B(n_1359),
.Y(n_1452)
);

OA21x2_ASAP7_75t_L g1453 ( 
.A1(n_1392),
.A2(n_1405),
.B(n_1417),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1416),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1354),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1382),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1389),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1395),
.B(n_1368),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1400),
.Y(n_1459)
);

OR2x6_ASAP7_75t_L g1460 ( 
.A(n_1383),
.B(n_1388),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1373),
.B(n_1380),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1413),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1375),
.B(n_1408),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1386),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1415),
.Y(n_1465)
);

AO21x2_ASAP7_75t_L g1466 ( 
.A1(n_1377),
.A2(n_1376),
.B(n_1406),
.Y(n_1466)
);

OR2x6_ASAP7_75t_L g1467 ( 
.A(n_1377),
.B(n_1372),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1357),
.B(n_1429),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1425),
.B(n_1427),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1365),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1352),
.Y(n_1471)
);

INVxp67_ASAP7_75t_SL g1472 ( 
.A(n_1367),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1381),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1359),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1423),
.B(n_1363),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1465),
.Y(n_1476)
);

INVx4_ASAP7_75t_L g1477 ( 
.A(n_1436),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1465),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1465),
.B(n_1394),
.Y(n_1479)
);

INVx8_ASAP7_75t_L g1480 ( 
.A(n_1460),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1462),
.B(n_1379),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1458),
.B(n_1391),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1462),
.B(n_1384),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1432),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1438),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1438),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1430),
.B(n_1385),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1433),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1459),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1440),
.B(n_1384),
.Y(n_1490)
);

OR2x6_ASAP7_75t_L g1491 ( 
.A(n_1432),
.B(n_1422),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1440),
.B(n_1391),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1474),
.B(n_1374),
.Y(n_1493)
);

INVx5_ASAP7_75t_L g1494 ( 
.A(n_1446),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1431),
.Y(n_1495)
);

NOR2x1_ASAP7_75t_L g1496 ( 
.A(n_1451),
.B(n_1390),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1444),
.B(n_1426),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1460),
.A2(n_1426),
.B(n_1424),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1454),
.B(n_1437),
.Y(n_1499)
);

OAI211xp5_ASAP7_75t_L g1500 ( 
.A1(n_1493),
.A2(n_1434),
.B(n_1448),
.C(n_1452),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1481),
.B(n_1443),
.Y(n_1501)
);

NOR4xp25_ASAP7_75t_SL g1502 ( 
.A(n_1496),
.B(n_1447),
.C(n_1434),
.D(n_1439),
.Y(n_1502)
);

INVx5_ASAP7_75t_L g1503 ( 
.A(n_1480),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1490),
.A2(n_1467),
.B1(n_1466),
.B2(n_1452),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1485),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1484),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1485),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1485),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1481),
.B(n_1443),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_L g1510 ( 
.A(n_1493),
.B(n_1448),
.C(n_1442),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1489),
.Y(n_1511)
);

OAI221xp5_ASAP7_75t_L g1512 ( 
.A1(n_1496),
.A2(n_1374),
.B1(n_1442),
.B2(n_1467),
.C(n_1471),
.Y(n_1512)
);

AOI221xp5_ASAP7_75t_L g1513 ( 
.A1(n_1498),
.A2(n_1474),
.B1(n_1472),
.B2(n_1475),
.C(n_1455),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1481),
.B(n_1443),
.Y(n_1514)
);

AND2x6_ASAP7_75t_SL g1515 ( 
.A(n_1491),
.B(n_1409),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1476),
.B(n_1435),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1495),
.B(n_1458),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1486),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1497),
.B(n_1472),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1476),
.B(n_1435),
.Y(n_1520)
);

NAND2xp33_ASAP7_75t_SL g1521 ( 
.A(n_1477),
.B(n_1447),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1476),
.B(n_1454),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1495),
.B(n_1463),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1496),
.A2(n_1467),
.B1(n_1441),
.B2(n_1460),
.Y(n_1524)
);

OAI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1491),
.A2(n_1467),
.B1(n_1441),
.B2(n_1446),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1478),
.B(n_1463),
.Y(n_1526)
);

INVxp67_ASAP7_75t_L g1527 ( 
.A(n_1490),
.Y(n_1527)
);

OAI221xp5_ASAP7_75t_L g1528 ( 
.A1(n_1491),
.A2(n_1445),
.B1(n_1451),
.B2(n_1461),
.C(n_1355),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1478),
.B(n_1454),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1479),
.B(n_1421),
.Y(n_1530)
);

AOI221xp5_ASAP7_75t_L g1531 ( 
.A1(n_1497),
.A2(n_1450),
.B1(n_1466),
.B2(n_1456),
.C(n_1464),
.Y(n_1531)
);

OAI221xp5_ASAP7_75t_L g1532 ( 
.A1(n_1491),
.A2(n_1445),
.B1(n_1451),
.B2(n_1461),
.C(n_1460),
.Y(n_1532)
);

OAI211xp5_ASAP7_75t_L g1533 ( 
.A1(n_1482),
.A2(n_1453),
.B(n_1456),
.C(n_1470),
.Y(n_1533)
);

AO21x2_ASAP7_75t_L g1534 ( 
.A1(n_1489),
.A2(n_1437),
.B(n_1449),
.Y(n_1534)
);

AOI21xp33_ASAP7_75t_L g1535 ( 
.A1(n_1500),
.A2(n_1466),
.B(n_1451),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1517),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1505),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1505),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1511),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1519),
.B(n_1488),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1507),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1506),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1516),
.B(n_1484),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1510),
.B(n_1531),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1507),
.Y(n_1545)
);

NOR3xp33_ASAP7_75t_L g1546 ( 
.A(n_1510),
.B(n_1473),
.C(n_1403),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1503),
.B(n_1484),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1530),
.B(n_1457),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1508),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1508),
.Y(n_1550)
);

NAND3xp33_ASAP7_75t_SL g1551 ( 
.A(n_1502),
.B(n_1482),
.C(n_1363),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1517),
.B(n_1482),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1523),
.B(n_1478),
.Y(n_1553)
);

AO21x2_ASAP7_75t_L g1554 ( 
.A1(n_1533),
.A2(n_1534),
.B(n_1525),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1503),
.B(n_1484),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1521),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1515),
.Y(n_1557)
);

NAND2x1p5_ASAP7_75t_L g1558 ( 
.A(n_1503),
.B(n_1494),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1522),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1523),
.Y(n_1560)
);

INVx4_ASAP7_75t_L g1561 ( 
.A(n_1503),
.Y(n_1561)
);

BUFx8_ASAP7_75t_L g1562 ( 
.A(n_1516),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1527),
.B(n_1488),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1526),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1513),
.B(n_1487),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1544),
.B(n_1520),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1556),
.B(n_1520),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1556),
.B(n_1522),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1557),
.B(n_1529),
.Y(n_1569)
);

CKINVDCx16_ASAP7_75t_R g1570 ( 
.A(n_1557),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1543),
.B(n_1529),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1544),
.B(n_1504),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1537),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1537),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1538),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1536),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1552),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1561),
.B(n_1503),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1546),
.B(n_1483),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1535),
.B(n_1483),
.Y(n_1580)
);

NOR3xp33_ASAP7_75t_L g1581 ( 
.A(n_1535),
.B(n_1512),
.C(n_1532),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1548),
.B(n_1468),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1552),
.B(n_1526),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1547),
.B(n_1501),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1539),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1560),
.B(n_1483),
.Y(n_1586)
);

NOR3xp33_ASAP7_75t_SL g1587 ( 
.A(n_1551),
.B(n_1528),
.C(n_1524),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1564),
.B(n_1518),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1538),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1541),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1541),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1545),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1547),
.B(n_1509),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1565),
.B(n_1509),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1540),
.B(n_1564),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1563),
.B(n_1540),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1545),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1549),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1547),
.B(n_1514),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1547),
.B(n_1514),
.Y(n_1600)
);

AND2x6_ASAP7_75t_SL g1601 ( 
.A(n_1555),
.B(n_1491),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1549),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1562),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1550),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1562),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1561),
.B(n_1503),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1570),
.B(n_1562),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1566),
.B(n_1563),
.Y(n_1608)
);

AOI32xp33_ASAP7_75t_L g1609 ( 
.A1(n_1581),
.A2(n_1555),
.A3(n_1561),
.B1(n_1559),
.B2(n_1492),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1566),
.B(n_1553),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1573),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1573),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1570),
.B(n_1555),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1576),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1585),
.Y(n_1615)
);

INVx4_ASAP7_75t_L g1616 ( 
.A(n_1603),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1572),
.B(n_1562),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1574),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1569),
.B(n_1468),
.Y(n_1619)
);

INVxp67_ASAP7_75t_SL g1620 ( 
.A(n_1605),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1574),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1585),
.Y(n_1622)
);

NAND2x1p5_ASAP7_75t_L g1623 ( 
.A(n_1578),
.B(n_1561),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1575),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1575),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_SL g1626 ( 
.A(n_1569),
.B(n_1551),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1579),
.B(n_1469),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1589),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1577),
.B(n_1469),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1589),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1590),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1585),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1590),
.Y(n_1633)
);

NAND2xp67_ASAP7_75t_SL g1634 ( 
.A(n_1567),
.B(n_1499),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1596),
.B(n_1553),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1571),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1571),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1591),
.Y(n_1638)
);

NAND2x1p5_ASAP7_75t_L g1639 ( 
.A(n_1578),
.B(n_1555),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1596),
.B(n_1550),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1594),
.B(n_1559),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1613),
.B(n_1567),
.Y(n_1642)
);

INVxp67_ASAP7_75t_SL g1643 ( 
.A(n_1613),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1612),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1610),
.B(n_1583),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1607),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1612),
.Y(n_1647)
);

INVxp67_ASAP7_75t_SL g1648 ( 
.A(n_1639),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1638),
.Y(n_1649)
);

INVxp33_ASAP7_75t_L g1650 ( 
.A(n_1617),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1639),
.Y(n_1651)
);

CKINVDCx16_ASAP7_75t_R g1652 ( 
.A(n_1616),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1638),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1611),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1614),
.Y(n_1655)
);

CKINVDCx16_ASAP7_75t_R g1656 ( 
.A(n_1616),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1610),
.B(n_1608),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1639),
.A2(n_1558),
.B(n_1542),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1620),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1609),
.A2(n_1587),
.B1(n_1580),
.B2(n_1558),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1618),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1621),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1616),
.B(n_1582),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1626),
.A2(n_1554),
.B1(n_1606),
.B2(n_1578),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1636),
.A2(n_1554),
.B1(n_1606),
.B2(n_1578),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1608),
.B(n_1583),
.Y(n_1666)
);

OAI21xp33_ASAP7_75t_L g1667 ( 
.A1(n_1643),
.A2(n_1637),
.B(n_1636),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1664),
.B(n_1623),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1659),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1642),
.B(n_1652),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1647),
.Y(n_1671)
);

NAND3xp33_ASAP7_75t_SL g1672 ( 
.A(n_1646),
.B(n_1623),
.C(n_1641),
.Y(n_1672)
);

AOI211xp5_ASAP7_75t_L g1673 ( 
.A1(n_1660),
.A2(n_1606),
.B(n_1624),
.C(n_1631),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1642),
.A2(n_1637),
.B1(n_1554),
.B2(n_1606),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1651),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1647),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1656),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1657),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1648),
.B(n_1663),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1655),
.A2(n_1554),
.B1(n_1568),
.B2(n_1584),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1649),
.Y(n_1681)
);

O2A1O1Ixp33_ASAP7_75t_L g1682 ( 
.A1(n_1650),
.A2(n_1623),
.B(n_1625),
.C(n_1628),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1665),
.A2(n_1595),
.B(n_1619),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1657),
.B(n_1627),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1651),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_SL g1686 ( 
.A(n_1682),
.B(n_1645),
.C(n_1666),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1677),
.B(n_1654),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1669),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_SL g1689 ( 
.A(n_1670),
.B(n_1651),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1679),
.B(n_1584),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1678),
.B(n_1654),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1669),
.Y(n_1692)
);

BUFx3_ASAP7_75t_L g1693 ( 
.A(n_1675),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1685),
.B(n_1661),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1671),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1680),
.B(n_1645),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1686),
.A2(n_1672),
.B(n_1668),
.Y(n_1697)
);

AOI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1696),
.A2(n_1672),
.B1(n_1668),
.B2(n_1667),
.C(n_1673),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1696),
.A2(n_1683),
.B(n_1674),
.Y(n_1699)
);

AOI21xp33_ASAP7_75t_L g1700 ( 
.A1(n_1689),
.A2(n_1684),
.B(n_1666),
.Y(n_1700)
);

OAI211xp5_ASAP7_75t_L g1701 ( 
.A1(n_1691),
.A2(n_1681),
.B(n_1676),
.C(n_1662),
.Y(n_1701)
);

AOI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1688),
.A2(n_1692),
.B1(n_1687),
.B2(n_1694),
.C(n_1690),
.Y(n_1702)
);

AOI311xp33_ASAP7_75t_L g1703 ( 
.A1(n_1693),
.A2(n_1662),
.A3(n_1661),
.B(n_1649),
.C(n_1653),
.Y(n_1703)
);

OAI21xp33_ASAP7_75t_L g1704 ( 
.A1(n_1693),
.A2(n_1644),
.B(n_1635),
.Y(n_1704)
);

OAI221xp5_ASAP7_75t_SL g1705 ( 
.A1(n_1695),
.A2(n_1635),
.B1(n_1630),
.B2(n_1633),
.C(n_1640),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1695),
.B(n_1629),
.Y(n_1706)
);

OA211x2_ASAP7_75t_L g1707 ( 
.A1(n_1689),
.A2(n_1586),
.B(n_1601),
.C(n_1634),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1704),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1700),
.B(n_1593),
.Y(n_1709)
);

OAI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1699),
.A2(n_1558),
.B1(n_1640),
.B2(n_1632),
.C(n_1615),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1698),
.A2(n_1568),
.B1(n_1658),
.B2(n_1600),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_SL g1712 ( 
.A(n_1705),
.B(n_1410),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1709),
.Y(n_1713)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1714 ( 
.A1(n_1710),
.A2(n_1697),
.B(n_1701),
.C(n_1706),
.D(n_1707),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1708),
.Y(n_1715)
);

AOI21xp33_ASAP7_75t_L g1716 ( 
.A1(n_1712),
.A2(n_1702),
.B(n_1658),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1711),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1709),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1713),
.Y(n_1719)
);

NAND3xp33_ASAP7_75t_SL g1720 ( 
.A(n_1717),
.B(n_1703),
.C(n_1632),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1713),
.Y(n_1721)
);

CKINVDCx16_ASAP7_75t_R g1722 ( 
.A(n_1715),
.Y(n_1722)
);

NAND2x1_ASAP7_75t_L g1723 ( 
.A(n_1718),
.B(n_1615),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1723),
.Y(n_1724)
);

AND3x4_ASAP7_75t_L g1725 ( 
.A(n_1722),
.B(n_1714),
.C(n_1716),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1721),
.B(n_1622),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1725),
.A2(n_1719),
.B1(n_1622),
.B2(n_1598),
.Y(n_1727)
);

INVx1_ASAP7_75t_SL g1728 ( 
.A(n_1727),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1728),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1729),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1730),
.A2(n_1724),
.B1(n_1726),
.B2(n_1720),
.Y(n_1731)
);

NAND2x1_ASAP7_75t_L g1732 ( 
.A(n_1731),
.B(n_1591),
.Y(n_1732)
);

OA22x2_ASAP7_75t_L g1733 ( 
.A1(n_1732),
.A2(n_1597),
.B1(n_1604),
.B2(n_1598),
.Y(n_1733)
);

AOI21xp33_ASAP7_75t_L g1734 ( 
.A1(n_1733),
.A2(n_1604),
.B(n_1592),
.Y(n_1734)
);

AOI22x1_ASAP7_75t_L g1735 ( 
.A1(n_1734),
.A2(n_1597),
.B1(n_1602),
.B2(n_1592),
.Y(n_1735)
);

AOI21xp33_ASAP7_75t_L g1736 ( 
.A1(n_1734),
.A2(n_1602),
.B(n_1588),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1735),
.A2(n_1588),
.B1(n_1593),
.B2(n_1599),
.Y(n_1737)
);

AOI211xp5_ASAP7_75t_L g1738 ( 
.A1(n_1737),
.A2(n_1736),
.B(n_1599),
.C(n_1600),
.Y(n_1738)
);


endmodule