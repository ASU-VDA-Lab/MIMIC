module fake_jpeg_27312_n_277 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_277);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVxp67_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_24),
.B1(n_26),
.B2(n_18),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_39),
.B(n_49),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_24),
.B1(n_26),
.B2(n_17),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_34),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_30),
.A2(n_17),
.B1(n_26),
.B2(n_24),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx2_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_53),
.A2(n_62),
.B(n_63),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_33),
.B1(n_36),
.B2(n_29),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_57),
.B1(n_45),
.B2(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_61),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_33),
.B1(n_36),
.B2(n_35),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_31),
.Y(n_61)
);

OR2x2_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_21),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_43),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_69),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_27),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_15),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_20),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_37),
.B1(n_42),
.B2(n_40),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_78),
.B1(n_80),
.B2(n_91),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_42),
.B1(n_36),
.B2(n_45),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_83),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_45),
.B1(n_35),
.B2(n_25),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_81),
.A2(n_90),
.B1(n_93),
.B2(n_58),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_20),
.Y(n_106)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_55),
.B(n_25),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_94),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_56),
.Y(n_109)
);

MAJx2_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_14),
.C(n_11),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_88),
.A2(n_96),
.B(n_85),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_22),
.B1(n_21),
.B2(n_19),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_53),
.A2(n_25),
.B1(n_22),
.B2(n_21),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_22),
.B1(n_19),
.B2(n_16),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_16),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_62),
.A2(n_16),
.B(n_19),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_69),
.B(n_70),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_62),
.A2(n_0),
.B(n_1),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_105),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_82),
.C(n_77),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_100),
.B(n_106),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_104),
.B(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_71),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_107),
.B(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_115),
.Y(n_125)
);

AO22x1_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_63),
.B1(n_72),
.B2(n_65),
.Y(n_110)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_83),
.A2(n_58),
.B1(n_67),
.B2(n_72),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_117),
.B1(n_119),
.B2(n_102),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_59),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_80),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_86),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_124),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_99),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_122),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g123 ( 
.A(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_146),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_96),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_92),
.B1(n_74),
.B2(n_89),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_133),
.A2(n_137),
.B(n_143),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_78),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_139),
.B(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_88),
.C(n_95),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_147),
.Y(n_160)
);

OR2x6_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_95),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_101),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_144),
.B(n_145),
.Y(n_176)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_88),
.C(n_81),
.Y(n_147)
);

AOI22x1_ASAP7_75t_L g148 ( 
.A1(n_114),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_148),
.A2(n_120),
.B1(n_115),
.B2(n_116),
.Y(n_151)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_66),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_151),
.A2(n_138),
.B1(n_148),
.B2(n_143),
.Y(n_182)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_153),
.Y(n_185)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_110),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_158),
.B(n_129),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_108),
.B(n_103),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_98),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_168),
.Y(n_190)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_166),
.Y(n_196)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_169),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_98),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_174),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_97),
.Y(n_177)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_74),
.C(n_14),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_155),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_121),
.C(n_124),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_183),
.C(n_195),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_174),
.A2(n_138),
.B1(n_136),
.B2(n_127),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_153),
.B1(n_178),
.B2(n_177),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_182),
.A2(n_193),
.B1(n_197),
.B2(n_191),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_143),
.C(n_148),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_189),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_187),
.B(n_188),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_164),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_151),
.A2(n_74),
.B1(n_66),
.B2(n_97),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_173),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_158),
.B(n_59),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_SL g211 ( 
.A(n_198),
.B(n_172),
.C(n_56),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_56),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_41),
.C(n_1),
.Y(n_214)
);

XNOR2x2_ASAP7_75t_SL g201 ( 
.A(n_159),
.B(n_8),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_15),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_185),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_204),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_184),
.B(n_150),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_203),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_190),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_209),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_179),
.A2(n_161),
.B1(n_168),
.B2(n_157),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_206),
.A2(n_211),
.B1(n_213),
.B2(n_198),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_161),
.B1(n_157),
.B2(n_171),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_216),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_187),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_11),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_215),
.A2(n_201),
.B(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_190),
.Y(n_217)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_191),
.Y(n_237)
);

O2A1O1Ixp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_194),
.B(n_188),
.C(n_183),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_221),
.B(n_223),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_226),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_180),
.C(n_195),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_207),
.C(n_212),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_182),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_226),
.C(n_228),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_240),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_212),
.C(n_196),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_230),
.C(n_220),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_218),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_239),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_219),
.B(n_204),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_215),
.B1(n_193),
.B2(n_214),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_244),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_229),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_12),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_248),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_222),
.C(n_10),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_254),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_234),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_251),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_238),
.A2(n_10),
.B(n_9),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_253),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_10),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_239),
.Y(n_255)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

O2A1O1Ixp33_ASAP7_75t_R g259 ( 
.A1(n_249),
.A2(n_242),
.B(n_9),
.C(n_8),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_251),
.Y(n_264)
);

NOR3xp33_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_8),
.C(n_6),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_261),
.B(n_255),
.Y(n_266)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

NOR2x1_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_250),
.Y(n_263)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

AOI21x1_ASAP7_75t_L g271 ( 
.A1(n_264),
.A2(n_267),
.B(n_5),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_246),
.C(n_248),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_266),
.C(n_256),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_258),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_269),
.A2(n_267),
.B(n_268),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_271),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_270),
.C(n_6),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_273),
.C(n_6),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_275),
.A2(n_7),
.B(n_258),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_7),
.B(n_204),
.Y(n_277)
);


endmodule