module real_jpeg_2993_n_7 (n_5, n_4, n_39, n_0, n_40, n_43, n_1, n_41, n_2, n_6, n_42, n_44, n_3, n_7);

input n_5;
input n_4;
input n_39;
input n_0;
input n_40;
input n_43;
input n_1;
input n_41;
input n_2;
input n_6;
input n_42;
input n_44;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_36;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AND2x2_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_9),
.Y(n_8)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

AO22x1_ASAP7_75t_L g14 ( 
.A1(n_4),
.A2(n_15),
.B1(n_19),
.B2(n_30),
.Y(n_14)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_14),
.C(n_31),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_6),
.A2(n_21),
.B(n_25),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_12),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_11),
.Y(n_9)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_33),
.C(n_34),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_17),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_18),
.Y(n_37)
);

NAND3xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_28),
.C(n_29),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_28),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_25),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_39),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_40),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_41),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_42),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_43),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_44),
.Y(n_36)
);


endmodule