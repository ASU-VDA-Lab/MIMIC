module fake_jpeg_1681_n_382 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_382);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_382;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_43),
.B(n_47),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_27),
.B(n_2),
.CON(n_56),
.SN(n_56)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_63),
.Y(n_88)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_2),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_58),
.B(n_73),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

OR2x4_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_12),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_26),
.B(n_12),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_26),
.B(n_13),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_34),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_71),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_23),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_78),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_32),
.B(n_2),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_20),
.B(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_75),
.B(n_28),
.Y(n_87)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_34),
.Y(n_79)
);

INVx6_ASAP7_75t_SL g121 ( 
.A(n_79),
.Y(n_121)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_31),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_80),
.Y(n_106)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

NAND3xp33_ASAP7_75t_L g149 ( 
.A(n_87),
.B(n_105),
.C(n_110),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_63),
.A2(n_75),
.B1(n_77),
.B2(n_70),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_89),
.A2(n_90),
.B1(n_94),
.B2(n_96),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_15),
.B1(n_39),
.B2(n_33),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_41),
.B1(n_15),
.B2(n_28),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_93),
.A2(n_115),
.B1(n_117),
.B2(n_130),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_15),
.B1(n_39),
.B2(n_33),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_46),
.A2(n_39),
.B1(n_33),
.B2(n_23),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_54),
.A2(n_23),
.B1(n_36),
.B2(n_76),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_99),
.A2(n_120),
.B1(n_129),
.B2(n_85),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_55),
.B(n_41),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_L g110 ( 
.A1(n_73),
.A2(n_40),
.B(n_38),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_67),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_123),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_42),
.A2(n_38),
.B1(n_35),
.B2(n_30),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_51),
.B(n_29),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_50),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_48),
.A2(n_35),
.B1(n_30),
.B2(n_29),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_61),
.A2(n_25),
.B1(n_37),
.B2(n_31),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_53),
.B(n_25),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_56),
.A2(n_13),
.B(n_11),
.C(n_5),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_13),
.B(n_4),
.C(n_5),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_61),
.A2(n_31),
.B1(n_4),
.B2(n_5),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_52),
.A2(n_60),
.B1(n_74),
.B2(n_68),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_132),
.Y(n_186)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_88),
.A2(n_125),
.B1(n_116),
.B2(n_57),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_135),
.A2(n_140),
.B1(n_151),
.B2(n_154),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_82),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_138),
.Y(n_193)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_139),
.B(n_142),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_88),
.A2(n_105),
.B1(n_114),
.B2(n_98),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_107),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_121),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_143),
.B(n_159),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_147),
.B(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_87),
.B(n_80),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_146),
.B(n_148),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_80),
.Y(n_148)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_103),
.A2(n_49),
.B1(n_62),
.B2(n_59),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_121),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_164),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_113),
.C(n_83),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_163),
.C(n_174),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_113),
.A2(n_81),
.B1(n_72),
.B2(n_31),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_3),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_106),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_158),
.B(n_160),
.Y(n_220)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_111),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_106),
.B(n_5),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_161),
.B(n_166),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_107),
.B(n_6),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_147),
.Y(n_207)
);

AND2x6_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_6),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_44),
.B1(n_8),
.B2(n_9),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_165),
.A2(n_172),
.B(n_132),
.C(n_171),
.Y(n_218)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_85),
.Y(n_167)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_107),
.B(n_7),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_169),
.Y(n_188)
);

AOI32xp33_ASAP7_75t_L g170 ( 
.A1(n_131),
.A2(n_7),
.A3(n_8),
.B1(n_102),
.B2(n_127),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_165),
.Y(n_197)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

CKINVDCx6p67_ASAP7_75t_R g172 ( 
.A(n_128),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_86),
.Y(n_173)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_179),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_95),
.A2(n_7),
.B1(n_124),
.B2(n_101),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_175),
.A2(n_176),
.B1(n_173),
.B2(n_150),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_91),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_92),
.A2(n_7),
.B1(n_119),
.B2(n_102),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_177),
.A2(n_162),
.B(n_141),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_128),
.A2(n_97),
.B(n_118),
.C(n_109),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_178),
.B(n_180),
.Y(n_213)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_101),
.Y(n_179)
);

AO22x1_ASAP7_75t_L g180 ( 
.A1(n_118),
.A2(n_109),
.B1(n_124),
.B2(n_104),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_95),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_182),
.B(n_205),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_134),
.A2(n_91),
.B1(n_104),
.B2(n_144),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_189),
.A2(n_191),
.B1(n_201),
.B2(n_202),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_146),
.A2(n_137),
.B1(n_148),
.B2(n_168),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_197),
.A2(n_215),
.B1(n_192),
.B2(n_195),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_185),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_133),
.B1(n_145),
.B2(n_180),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_151),
.B1(n_154),
.B2(n_178),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_149),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_207),
.B(n_192),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_172),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_211),
.B(n_190),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_167),
.A2(n_172),
.B(n_164),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_SL g240 ( 
.A1(n_218),
.A2(n_209),
.B(n_213),
.C(n_219),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_156),
.A2(n_141),
.B1(n_162),
.B2(n_136),
.Y(n_219)
);

AO21x2_ASAP7_75t_L g235 ( 
.A1(n_219),
.A2(n_221),
.B(n_213),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_221),
.Y(n_256)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_223),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_224),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_225),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_217),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_226),
.B(n_227),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_200),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_182),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_234),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_217),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_233),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_197),
.A2(n_209),
.B(n_207),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_230),
.A2(n_244),
.B(n_186),
.Y(n_257)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_231),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_232),
.B(n_184),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_214),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_185),
.B(n_198),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_235),
.A2(n_184),
.B1(n_256),
.B2(n_240),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_183),
.B(n_206),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_241),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_220),
.B(n_206),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_246),
.Y(n_271)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_199),
.Y(n_238)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_238),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

OA21x2_ASAP7_75t_L g282 ( 
.A1(n_240),
.A2(n_235),
.B(n_243),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_183),
.B(n_211),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_196),
.B(n_197),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_247),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_218),
.A2(n_214),
.B(n_212),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_245),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_208),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_212),
.A2(n_188),
.B1(n_205),
.B2(n_195),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_248),
.A2(n_251),
.B1(n_234),
.B2(n_242),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_216),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_249),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_208),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_252),
.Y(n_268)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_199),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_253),
.A2(n_254),
.B1(n_186),
.B2(n_210),
.Y(n_266)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_204),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_255),
.B(n_242),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_257),
.B(n_266),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_259),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_230),
.A2(n_194),
.B(n_187),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_270),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_256),
.A2(n_194),
.B(n_187),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_232),
.B(n_215),
.C(n_187),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_274),
.C(n_283),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_222),
.A2(n_184),
.B1(n_244),
.B2(n_235),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_275),
.A2(n_277),
.B1(n_281),
.B2(n_285),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_222),
.A2(n_235),
.B1(n_241),
.B2(n_228),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_278),
.A2(n_269),
.B1(n_257),
.B2(n_282),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_225),
.A2(n_248),
.B(n_240),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_240),
.Y(n_300)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_236),
.B(n_250),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_229),
.B(n_246),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_239),
.C(n_274),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_287),
.B(n_283),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_271),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_288),
.A2(n_304),
.B1(n_309),
.B2(n_307),
.Y(n_330)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_263),
.B(n_231),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_296),
.Y(n_314)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_292),
.Y(n_326)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_293),
.Y(n_328)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_262),
.Y(n_294)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_294),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_235),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_302),
.C(n_261),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_258),
.B(n_238),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_286),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_298),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_300),
.A2(n_301),
.B(n_310),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_245),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_265),
.B(n_254),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_273),
.Y(n_318)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_280),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_307),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_268),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_308),
.A2(n_261),
.B1(n_264),
.B2(n_270),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_265),
.B(n_284),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_268),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_259),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_319),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_301),
.A2(n_279),
.B(n_272),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_316),
.A2(n_317),
.B(n_299),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_297),
.A2(n_282),
.B(n_272),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_299),
.C(n_292),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_321),
.B(n_327),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_323),
.A2(n_324),
.B1(n_325),
.B2(n_322),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_289),
.A2(n_264),
.B1(n_286),
.B2(n_266),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_289),
.A2(n_260),
.B1(n_280),
.B2(n_310),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_295),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_329),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_303),
.B(n_305),
.Y(n_329)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_330),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_314),
.Y(n_331)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_331),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_293),
.Y(n_332)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_332),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_315),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_333),
.B(n_339),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_323),
.A2(n_302),
.B1(n_297),
.B2(n_299),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_334),
.A2(n_324),
.B1(n_320),
.B2(n_325),
.Y(n_356)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_335),
.Y(n_351)
);

XNOR2x1_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_316),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_329),
.B(n_294),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_328),
.B(n_290),
.Y(n_340)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_340),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_320),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_341),
.B(n_345),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_297),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_344),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_318),
.B(n_319),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_346),
.B(n_317),
.C(n_312),
.Y(n_358)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_343),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_353),
.B(n_357),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_355),
.B(n_342),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_356),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_346),
.B(n_313),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_358),
.B(n_352),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_336),
.C(n_338),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_359),
.B(n_360),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_354),
.A2(n_334),
.B(n_313),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_357),
.A2(n_349),
.B(n_348),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_361),
.A2(n_350),
.B1(n_351),
.B2(n_356),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_362),
.B(n_363),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_347),
.B(n_336),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_366),
.A2(n_352),
.B1(n_313),
.B2(n_326),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_367),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_359),
.B(n_338),
.C(n_344),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_371),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_364),
.A2(n_351),
.B1(n_365),
.B2(n_363),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_372),
.B(n_364),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_374),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_368),
.B(n_369),
.C(n_370),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_376),
.B(n_370),
.Y(n_378)
);

A2O1A1O1Ixp25_ASAP7_75t_L g379 ( 
.A1(n_378),
.A2(n_375),
.B(n_373),
.C(n_371),
.D(n_337),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_377),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_380),
.A2(n_322),
.B1(n_306),
.B2(n_355),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_298),
.Y(n_382)
);


endmodule