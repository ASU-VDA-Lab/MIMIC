module fake_jpeg_21329_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_42),
.Y(n_59)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_48),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_18),
.B1(n_21),
.B2(n_26),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_62),
.B1(n_36),
.B2(n_23),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_27),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_51),
.B(n_27),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_21),
.B1(n_26),
.B2(n_16),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_37),
.B1(n_18),
.B2(n_21),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_26),
.B1(n_22),
.B2(n_20),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_66),
.A2(n_39),
.B1(n_44),
.B2(n_37),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_77),
.Y(n_109)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

NAND2x1_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_39),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_74),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_75),
.A2(n_92),
.B1(n_93),
.B2(n_99),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_83),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_80),
.A2(n_102),
.B1(n_52),
.B2(n_43),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_31),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_64),
.A2(n_39),
.B1(n_22),
.B2(n_34),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_84),
.A2(n_104),
.B1(n_75),
.B2(n_78),
.Y(n_111)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_88),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_89),
.B(n_100),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_53),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_91),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_63),
.Y(n_94)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_94),
.Y(n_124)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

FAx1_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_45),
.CI(n_43),
.CON(n_97),
.SN(n_97)
);

FAx1_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_107),
.CI(n_108),
.CON(n_112),
.SN(n_112)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_31),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_49),
.A2(n_22),
.B1(n_34),
.B2(n_32),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_56),
.A2(n_32),
.B1(n_20),
.B2(n_23),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_111),
.A2(n_117),
.B1(n_126),
.B2(n_133),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_61),
.C(n_45),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_95),
.C(n_88),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_78),
.A2(n_52),
.B1(n_45),
.B2(n_43),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_120),
.A2(n_86),
.B1(n_29),
.B2(n_99),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_80),
.A2(n_25),
.B1(n_24),
.B2(n_19),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_129),
.B1(n_132),
.B2(n_135),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_97),
.A2(n_43),
.B1(n_41),
.B2(n_40),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_25),
.B1(n_24),
.B2(n_19),
.Y(n_129)
);

AO21x2_ASAP7_75t_SL g130 ( 
.A1(n_74),
.A2(n_41),
.B(n_40),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_81),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_70),
.A2(n_25),
.B1(n_24),
.B2(n_19),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_41),
.B1(n_40),
.B2(n_29),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_41),
.B1(n_10),
.B2(n_11),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_139),
.A2(n_146),
.B(n_169),
.Y(n_199)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_140),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_111),
.A2(n_68),
.B1(n_71),
.B2(n_105),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_141),
.A2(n_164),
.B1(n_118),
.B2(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

BUFx8_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_148),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_138),
.A2(n_76),
.B(n_84),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_87),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_150),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_86),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_138),
.A2(n_96),
.B1(n_98),
.B2(n_87),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_149),
.B(n_122),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_91),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_115),
.B(n_124),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_165),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_115),
.B(n_15),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_159),
.B(n_12),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_69),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_155),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_82),
.Y(n_156)
);

AO22x1_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_114),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_72),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_14),
.C(n_15),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_129),
.A2(n_73),
.B1(n_103),
.B2(n_68),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_162),
.B1(n_163),
.B2(n_130),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_109),
.A2(n_29),
.B(n_17),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_135),
.B(n_131),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_125),
.B1(n_126),
.B2(n_134),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_130),
.A2(n_29),
.B1(n_28),
.B2(n_17),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_110),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_137),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_128),
.B1(n_127),
.B2(n_27),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_130),
.A2(n_133),
.B(n_117),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_170),
.B(n_176),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_172),
.A2(n_179),
.B(n_180),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_173),
.A2(n_183),
.B1(n_142),
.B2(n_144),
.Y(n_218)
);

XOR2x2_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_132),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_137),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_198),
.B1(n_201),
.B2(n_142),
.Y(n_214)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_118),
.B1(n_116),
.B2(n_128),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_123),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_150),
.Y(n_206)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_186),
.B(n_188),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_187),
.A2(n_0),
.B(n_1),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_143),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_147),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_190),
.B(n_196),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_191),
.A2(n_161),
.B1(n_140),
.B2(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_193),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_127),
.C(n_28),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_146),
.C(n_156),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_149),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_127),
.B1(n_31),
.B2(n_28),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_144),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_153),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_154),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_204),
.B(n_228),
.C(n_202),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_205),
.B(n_215),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_206),
.B(n_194),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_207),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_192),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_158),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_213),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_154),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_214),
.A2(n_226),
.B1(n_231),
.B2(n_178),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_193),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_164),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_216),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_218),
.A2(n_189),
.B1(n_175),
.B2(n_174),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_196),
.A2(n_144),
.B1(n_152),
.B2(n_2),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_220),
.A2(n_222),
.B(n_227),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_199),
.A2(n_0),
.B(n_1),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_223),
.A2(n_229),
.B(n_230),
.Y(n_235)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_178),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_224),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_180),
.A2(n_179),
.B1(n_173),
.B2(n_197),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_174),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_3),
.C(n_4),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_199),
.A2(n_9),
.B(n_4),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_180),
.A2(n_9),
.B(n_4),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_197),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_232),
.A2(n_234),
.B1(n_226),
.B2(n_225),
.Y(n_260)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_183),
.B1(n_185),
.B2(n_175),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_237),
.Y(n_268)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_238),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_217),
.A2(n_172),
.B(n_176),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_241),
.A2(n_244),
.B(n_222),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_245),
.Y(n_273)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_243),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_229),
.A2(n_176),
.B(n_182),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_177),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_177),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_251),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_195),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_252),
.B1(n_210),
.B2(n_230),
.Y(n_258)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_209),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_228),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_211),
.C(n_204),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_256),
.C(n_262),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_225),
.C(n_217),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_263),
.Y(n_279)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_264),
.B1(n_270),
.B2(n_259),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_241),
.B(n_220),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_234),
.A2(n_214),
.B1(n_209),
.B2(n_231),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_242),
.C(n_245),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_223),
.B(n_203),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_224),
.C(n_227),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_269),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_232),
.A2(n_202),
.B1(n_7),
.B2(n_8),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_235),
.B(n_6),
.Y(n_274)
);

NOR2xp67_ASAP7_75t_SL g278 ( 
.A(n_274),
.B(n_235),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_238),
.Y(n_276)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_278),
.A2(n_285),
.B1(n_287),
.B2(n_288),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_283),
.Y(n_295)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

INVxp33_ASAP7_75t_SL g284 ( 
.A(n_272),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_284),
.A2(n_236),
.B(n_254),
.Y(n_302)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_246),
.B1(n_243),
.B2(n_237),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_261),
.B1(n_252),
.B2(n_233),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_277),
.B(n_250),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_296),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_284),
.A2(n_246),
.B1(n_274),
.B2(n_254),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_276),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_256),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_279),
.Y(n_310)
);

FAx1_ASAP7_75t_SL g296 ( 
.A(n_279),
.B(n_260),
.CI(n_263),
.CON(n_296),
.SN(n_296)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_299),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_266),
.C(n_255),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_275),
.A2(n_257),
.B(n_267),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_300),
.A2(n_275),
.B(n_240),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_262),
.C(n_273),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_302),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_286),
.C(n_273),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_309),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_305),
.A2(n_292),
.B1(n_297),
.B2(n_296),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_311),
.B(n_302),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_282),
.B1(n_247),
.B2(n_289),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_301),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_240),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_314),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_294),
.Y(n_314)
);

OAI21x1_ASAP7_75t_L g318 ( 
.A1(n_315),
.A2(n_307),
.B(n_311),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_317),
.B(n_6),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_296),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_318),
.B(n_321),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_304),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_319),
.A2(n_312),
.B(n_313),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_322),
.Y(n_324)
);

OAI311xp33_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_320),
.A3(n_323),
.B1(n_8),
.C1(n_6),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_7),
.C(n_8),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_8),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);


endmodule