module fake_jpeg_10412_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_28),
.Y(n_53)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_8),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_40),
.Y(n_47)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_8),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_16),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_57),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_28),
.B1(n_26),
.B2(n_23),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_52),
.B1(n_55),
.B2(n_18),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_32),
.A2(n_28),
.B1(n_23),
.B2(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_55),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_25),
.B(n_15),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_29),
.C(n_17),
.Y(n_82)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_60),
.B(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_65),
.Y(n_84)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_42),
.B1(n_35),
.B2(n_27),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_70),
.B(n_76),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

NAND2x1_ASAP7_75t_SL g70 ( 
.A(n_58),
.B(n_39),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_77),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_43),
.A2(n_42),
.B1(n_35),
.B2(n_39),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_41),
.B1(n_58),
.B2(n_45),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_47),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_30),
.B1(n_29),
.B2(n_18),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_53),
.B(n_17),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_25),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_0),
.Y(n_81)
);

HAxp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_82),
.CON(n_97),
.SN(n_97)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_27),
.B1(n_21),
.B2(n_33),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_57),
.B1(n_41),
.B2(n_46),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_79),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_105),
.C(n_71),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_95),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_56),
.B1(n_46),
.B2(n_33),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_94),
.B1(n_65),
.B2(n_86),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_90),
.B(n_103),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_47),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_91),
.B(n_101),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_80),
.B(n_67),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_68),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_100),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_66),
.A2(n_41),
.B1(n_37),
.B2(n_44),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_67),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_41),
.B1(n_37),
.B2(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_19),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_37),
.B1(n_19),
.B2(n_15),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_1),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_24),
.C(n_22),
.Y(n_105)
);

XOR2x1_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_81),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_121),
.B(n_91),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_110),
.A2(n_115),
.B(n_119),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_84),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_89),
.B1(n_99),
.B2(n_96),
.Y(n_136)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_117),
.C(n_120),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_70),
.C(n_72),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_84),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_72),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_77),
.B(n_72),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_124),
.B(n_100),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_72),
.B1(n_68),
.B2(n_64),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_125),
.A2(n_64),
.B1(n_68),
.B2(n_95),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_129),
.B(n_138),
.Y(n_150)
);

AOI21x1_ASAP7_75t_SL g130 ( 
.A1(n_117),
.A2(n_86),
.B(n_93),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_131),
.B(n_137),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_106),
.C(n_108),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_135),
.C(n_114),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_105),
.C(n_98),
.Y(n_135)
);

AOI221xp5_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_143),
.B1(n_144),
.B2(n_125),
.C(n_113),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_102),
.B(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_126),
.B(n_105),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_126),
.B(n_11),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_147),
.A2(n_160),
.B1(n_164),
.B2(n_143),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_112),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_149),
.C(n_151),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_121),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_123),
.C(n_124),
.Y(n_152)
);

OAI322xp33_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_24),
.A3(n_10),
.B1(n_14),
.B2(n_4),
.C1(n_6),
.C2(n_7),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_135),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_153),
.B(n_156),
.Y(n_167)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_123),
.C(n_115),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_163),
.B(n_145),
.Y(n_165)
);

INVxp67_ASAP7_75t_SL g159 ( 
.A(n_128),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_109),
.B1(n_117),
.B2(n_119),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_107),
.C(n_75),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_130),
.A2(n_138),
.B1(n_133),
.B2(n_128),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_156),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_130),
.B(n_137),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_168),
.A2(n_170),
.B1(n_172),
.B2(n_174),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_145),
.B(n_140),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_133),
.B1(n_139),
.B2(n_132),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_132),
.B1(n_136),
.B2(n_141),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_161),
.A2(n_107),
.B1(n_146),
.B2(n_144),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_176),
.B(n_179),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_158),
.A2(n_87),
.B1(n_69),
.B2(n_24),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_162),
.A2(n_87),
.B1(n_10),
.B2(n_11),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_155),
.A2(n_10),
.B(n_14),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_150),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_180),
.B(n_168),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_183),
.C(n_185),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_184),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_151),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_153),
.C(n_148),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_189),
.C(n_185),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_155),
.C(n_162),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_175),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_154),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_187),
.C(n_188),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_177),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_199),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_4),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_SL g195 ( 
.A(n_189),
.B(n_171),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_195),
.A2(n_196),
.B(n_171),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_200),
.C(n_191),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_178),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_202),
.B(n_194),
.Y(n_213)
);

AOI31xp33_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_180),
.A3(n_11),
.B(n_12),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_203),
.A2(n_9),
.B(n_13),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_87),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_205),
.Y(n_210)
);

NAND4xp25_ASAP7_75t_SL g205 ( 
.A(n_198),
.B(n_69),
.C(n_2),
.D(n_3),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_9),
.Y(n_209)
);

INVxp33_ASAP7_75t_SL g208 ( 
.A(n_205),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_208),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_211),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_212),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_201),
.C(n_204),
.Y(n_215)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_215),
.A2(n_1),
.B(n_2),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_210),
.B1(n_4),
.B2(n_7),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_220),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_214),
.A2(n_12),
.B(n_13),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_219),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_221),
.A2(n_2),
.B1(n_217),
.B2(n_222),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_223),
.B(n_2),
.Y(n_224)
);


endmodule