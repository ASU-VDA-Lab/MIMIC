module fake_jpeg_19603_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_42),
.Y(n_53)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_43),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_26),
.Y(n_77)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_63),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_61),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_20),
.B1(n_33),
.B2(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_20),
.Y(n_63)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_68),
.Y(n_95)
);

CKINVDCx12_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_33),
.B1(n_39),
.B2(n_23),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_69),
.Y(n_113)
);

HAxp5_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_20),
.CON(n_71),
.SN(n_71)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_71),
.A2(n_16),
.B(n_21),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_72),
.B(n_77),
.Y(n_109)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_81),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_74),
.Y(n_107)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_54),
.Y(n_76)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_80),
.B(n_82),
.Y(n_119)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_88),
.Y(n_93)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_16),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_48),
.B(n_40),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_37),
.C(n_45),
.Y(n_112)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_45),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_96),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_45),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_48),
.B1(n_33),
.B2(n_44),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_97),
.A2(n_101),
.B1(n_108),
.B2(n_92),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_78),
.B1(n_48),
.B2(n_84),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_29),
.B(n_21),
.Y(n_103)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_103),
.A2(n_104),
.A3(n_25),
.B1(n_28),
.B2(n_26),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_31),
.B1(n_23),
.B2(n_19),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_52),
.B1(n_58),
.B2(n_31),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_115),
.C(n_120),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_37),
.C(n_45),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_37),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_122),
.B(n_24),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_89),
.B1(n_83),
.B2(n_87),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_128),
.B1(n_129),
.B2(n_134),
.Y(n_152)
);

AO22x1_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_87),
.B1(n_91),
.B2(n_54),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_76),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_127),
.B(n_130),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_93),
.A2(n_86),
.B1(n_75),
.B2(n_62),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_37),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_30),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_132),
.B(n_138),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_93),
.A2(n_62),
.B1(n_55),
.B2(n_30),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_94),
.A2(n_79),
.B1(n_12),
.B2(n_13),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_136),
.A2(n_104),
.B1(n_119),
.B2(n_99),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_102),
.A2(n_28),
.B1(n_25),
.B2(n_27),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_100),
.B1(n_102),
.B2(n_117),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_118),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_148),
.B(n_120),
.Y(n_170)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

CKINVDCx12_ASAP7_75t_R g147 ( 
.A(n_95),
.Y(n_147)
);

INVxp33_ASAP7_75t_SL g150 ( 
.A(n_147),
.Y(n_150)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_154),
.A2(n_160),
.B1(n_179),
.B2(n_24),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_135),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_155),
.B(n_168),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_112),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_161),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_139),
.B1(n_143),
.B2(n_136),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_122),
.Y(n_161)
);

NAND2x1p5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_120),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_170),
.B(n_24),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_133),
.B1(n_111),
.B2(n_123),
.Y(n_197)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_126),
.A2(n_107),
.B(n_121),
.C(n_98),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_172),
.Y(n_203)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_107),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_137),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_174),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_98),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_103),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_175),
.B(n_131),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_137),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_79),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_124),
.A2(n_117),
.B1(n_99),
.B2(n_110),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_177),
.A2(n_125),
.B1(n_110),
.B2(n_111),
.Y(n_195)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_126),
.A2(n_131),
.B1(n_141),
.B2(n_144),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_180),
.B(n_198),
.C(n_165),
.Y(n_226)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_190),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_151),
.B(n_163),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_184),
.A2(n_189),
.B(n_206),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_149),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_199),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_125),
.B(n_133),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx6_ASAP7_75t_SL g191 ( 
.A(n_150),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_192),
.Y(n_230)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

OR2x2_ASAP7_75t_SL g193 ( 
.A(n_156),
.B(n_28),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_SL g218 ( 
.A1(n_193),
.A2(n_208),
.B(n_177),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_158),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_168),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_197),
.B1(n_176),
.B2(n_173),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_175),
.B(n_26),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_196),
.B(n_205),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_26),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_178),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_201),
.B(n_207),
.Y(n_225)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_154),
.B(n_26),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_153),
.A2(n_27),
.B(n_25),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_162),
.Y(n_207)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_79),
.B1(n_10),
.B2(n_11),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_210),
.A2(n_152),
.B1(n_167),
.B2(n_165),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_162),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_24),
.Y(n_235)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_179),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_223),
.Y(n_249)
);

AOI21xp33_ASAP7_75t_L g217 ( 
.A1(n_199),
.A2(n_161),
.B(n_153),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_217),
.A2(n_206),
.B(n_210),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_218),
.A2(n_219),
.B1(n_189),
.B2(n_234),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g221 ( 
.A(n_194),
.Y(n_221)
);

BUFx24_ASAP7_75t_SL g242 ( 
.A(n_221),
.Y(n_242)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_228),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_188),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_182),
.A2(n_172),
.B1(n_152),
.B2(n_156),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_227),
.A2(n_182),
.B1(n_208),
.B2(n_203),
.Y(n_238)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_171),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_229),
.Y(n_243)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_231),
.Y(n_246)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_232),
.B(n_235),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_195),
.B1(n_209),
.B2(n_181),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_191),
.B(n_24),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_237),
.B(n_0),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_238),
.A2(n_250),
.B1(n_233),
.B2(n_215),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_198),
.C(n_186),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_257),
.C(n_222),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_241),
.A2(n_219),
.B1(n_220),
.B2(n_234),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_245),
.A2(n_213),
.B1(n_214),
.B2(n_224),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_227),
.B(n_184),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_255),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_180),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_253),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_216),
.A2(n_202),
.B1(n_200),
.B2(n_188),
.Y(n_251)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_236),
.B(n_183),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_254),
.B(n_258),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_185),
.C(n_181),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_229),
.B(n_185),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_258),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_262),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_265),
.A2(n_271),
.B1(n_272),
.B2(n_246),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_225),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_266),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_267),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_230),
.C(n_231),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_22),
.C(n_32),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_256),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_275),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_238),
.A2(n_223),
.B1(n_10),
.B2(n_11),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_9),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_273),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_241),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_6),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_276),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_274),
.B(n_242),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_277),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_278),
.A2(n_259),
.B1(n_265),
.B2(n_264),
.Y(n_298)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_246),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_286),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_239),
.Y(n_286)
);

OA21x2_ASAP7_75t_SL g288 ( 
.A1(n_260),
.A2(n_253),
.B(n_248),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_289),
.B(n_6),
.Y(n_293)
);

OA21x2_ASAP7_75t_SL g289 ( 
.A1(n_269),
.A2(n_6),
.B(n_12),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_290),
.B(n_291),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_0),
.Y(n_291)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_268),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_297),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_280),
.B(n_261),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_298),
.A2(n_279),
.B1(n_11),
.B2(n_5),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_264),
.C(n_270),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_300),
.C(n_283),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_270),
.C(n_27),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_290),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_302),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_287),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_32),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_278),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_306),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_282),
.C(n_291),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_310),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_304),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_279),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_312),
.B(n_313),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_32),
.C(n_5),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_314),
.B(n_0),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_308),
.A2(n_292),
.B(n_295),
.Y(n_315)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_315),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_318),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_311),
.B(n_303),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_310),
.A2(n_300),
.B(n_2),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_1),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_309),
.B(n_312),
.Y(n_324)
);

OAI21x1_ASAP7_75t_L g327 ( 
.A1(n_324),
.A2(n_320),
.B(n_316),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_2),
.Y(n_326)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_327),
.C(n_323),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_322),
.C(n_305),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_3),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_3),
.B(n_4),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_3),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_3),
.B(n_4),
.Y(n_333)
);


endmodule