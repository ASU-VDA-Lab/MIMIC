module fake_netlist_6_3049_n_2146 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2146);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2146;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1794;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g220 ( 
.A(n_70),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_123),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_36),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_160),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_0),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_89),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_51),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_94),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_29),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_159),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_105),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_46),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_201),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_5),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_109),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_57),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_68),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_208),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_212),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_59),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_129),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_43),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_192),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_126),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_80),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_8),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_48),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_72),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_79),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_43),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_187),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_172),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_62),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_93),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_60),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_60),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_155),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_147),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_36),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_97),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_132),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_218),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_138),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_14),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_114),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_78),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_113),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_16),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_25),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_15),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_90),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_135),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_115),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_170),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_5),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_195),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_108),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_102),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_110),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_158),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_207),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_168),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_139),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_78),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_178),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_157),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_206),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_119),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_1),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_156),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_76),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_118),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_104),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_169),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_1),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_3),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_72),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_112),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_100),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_29),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_40),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_6),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_65),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_26),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_210),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_26),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_203),
.Y(n_308)
);

BUFx8_ASAP7_75t_SL g309 ( 
.A(n_95),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_39),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_27),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_197),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_163),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_202),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_96),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_47),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_4),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_47),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_88),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_17),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_186),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_133),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_140),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_39),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_32),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_13),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_134),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_33),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_33),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_16),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_161),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_41),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_86),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_66),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_38),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_83),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_185),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_51),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_28),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_49),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_213),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_106),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_180),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_70),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_98),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_44),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_188),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_53),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_107),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_66),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_6),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_209),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_116),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_211),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_62),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_120),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_141),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_103),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_81),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_121),
.Y(n_360)
);

BUFx2_ASAP7_75t_SL g361 ( 
.A(n_184),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_171),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_143),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_125),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_167),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_217),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_7),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_189),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_136),
.Y(n_369)
);

INVxp33_ASAP7_75t_SL g370 ( 
.A(n_193),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_24),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_151),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_19),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_154),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_124),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_130),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_87),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_199),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_85),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_131),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_183),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_214),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_10),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_71),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_44),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_3),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_38),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_55),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_57),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_67),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_69),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_216),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_127),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_21),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_58),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_14),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_25),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_164),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_82),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_194),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_0),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_59),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_71),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_111),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_10),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_219),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_64),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_7),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_61),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_12),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_144),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_165),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_149),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_182),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_148),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_176),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_173),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_11),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_18),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_41),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_35),
.Y(n_421)
);

INVxp33_ASAP7_75t_L g422 ( 
.A(n_37),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_49),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_91),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_31),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_19),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_50),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_137),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_11),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_152),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_34),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_290),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_240),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_227),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_290),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_309),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_290),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_278),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_290),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_290),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_288),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_282),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_315),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_280),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_393),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_284),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_287),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_294),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_232),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_325),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_325),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_295),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_300),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_325),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_306),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_325),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_325),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_308),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_321),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_333),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_272),
.B(n_2),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_326),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_326),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_326),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_326),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_322),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_326),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_336),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_342),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_343),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_347),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_240),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_349),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_354),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_260),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_385),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_356),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_359),
.B(n_2),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_385),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_224),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_360),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_385),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_385),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_224),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_388),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_362),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_228),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_365),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_388),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_366),
.Y(n_491)
);

BUFx6f_ASAP7_75t_SL g492 ( 
.A(n_235),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_L g493 ( 
.A(n_276),
.B(n_4),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_285),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_260),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_292),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_297),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_401),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_298),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_401),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_301),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_370),
.B(n_8),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_316),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_279),
.B(n_9),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_316),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_330),
.Y(n_506)
);

INVx4_ASAP7_75t_R g507 ( 
.A(n_235),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_220),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_302),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_221),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_330),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_226),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_237),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_228),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_305),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_311),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_248),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_250),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_274),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_256),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_318),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_221),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_320),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_265),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_303),
.Y(n_525)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_257),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_223),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_304),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_307),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_310),
.Y(n_530)
);

INVxp33_ASAP7_75t_L g531 ( 
.A(n_422),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_317),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_274),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_332),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_293),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_223),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_334),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_335),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_293),
.Y(n_539)
);

INVxp33_ASAP7_75t_SL g540 ( 
.A(n_234),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_340),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_225),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_344),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_346),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_348),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_367),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_383),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_225),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_350),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_234),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_494),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_452),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_458),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_468),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_470),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_456),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_519),
.B(n_299),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_432),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_456),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_434),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_438),
.B(n_299),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_435),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_496),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_473),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_435),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_437),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_437),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_442),
.B(n_313),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_482),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_439),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_533),
.B(n_313),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_439),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_440),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_440),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_535),
.B(n_296),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_450),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_487),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_450),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_443),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_451),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_535),
.B(n_279),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_451),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_454),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_480),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_454),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_539),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_457),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_510),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_457),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_446),
.B(n_291),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_531),
.A2(n_236),
.B1(n_246),
.B2(n_242),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_539),
.B(n_291),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_488),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_462),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_436),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_462),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_522),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_527),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_463),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_L g600 ( 
.A(n_461),
.B(n_431),
.C(n_242),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_441),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_463),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_536),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_542),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_548),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_464),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_447),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_504),
.B(n_252),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_464),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_465),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_465),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_503),
.B(n_296),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_448),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_453),
.B(n_455),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_497),
.B(n_312),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_467),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_467),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_476),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_514),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_476),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_479),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_479),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_481),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_481),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_483),
.Y(n_625)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_491),
.B(n_329),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_483),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_459),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_460),
.Y(n_629)
);

INVx5_ASAP7_75t_L g630 ( 
.A(n_475),
.Y(n_630)
);

AND3x2_ASAP7_75t_L g631 ( 
.A(n_478),
.B(n_264),
.C(n_249),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_484),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_484),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_469),
.B(n_312),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_499),
.B(n_353),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_503),
.B(n_387),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_501),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_471),
.B(n_353),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_505),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_509),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_486),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_445),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_570),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_639),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_570),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_556),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_556),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_558),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_615),
.B(n_474),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_586),
.Y(n_650)
);

BUFx10_ASAP7_75t_L g651 ( 
.A(n_607),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_607),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_570),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_570),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_SL g655 ( 
.A(n_575),
.B(n_338),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_635),
.B(n_477),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_586),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_562),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_630),
.B(n_557),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_590),
.B(n_489),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_559),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_559),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_SL g663 ( 
.A(n_613),
.B(n_628),
.Y(n_663)
);

OR2x6_ASAP7_75t_L g664 ( 
.A(n_614),
.B(n_361),
.Y(n_664)
);

BUFx10_ASAP7_75t_L g665 ( 
.A(n_613),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_570),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_630),
.B(n_502),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_557),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_608),
.A2(n_444),
.B1(n_466),
.B2(n_449),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_557),
.B(n_515),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_566),
.Y(n_671)
);

OAI22xp33_ASAP7_75t_SL g672 ( 
.A1(n_634),
.A2(n_638),
.B1(n_568),
.B2(n_561),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_565),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_571),
.B(n_516),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_630),
.B(n_249),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_567),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_582),
.Y(n_677)
);

INVxp33_ASAP7_75t_L g678 ( 
.A(n_575),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_571),
.B(n_521),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_585),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_576),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_576),
.Y(n_682)
);

BUFx10_ASAP7_75t_L g683 ( 
.A(n_628),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_596),
.Y(n_684)
);

OAI22xp33_ASAP7_75t_L g685 ( 
.A1(n_600),
.A2(n_339),
.B1(n_403),
.B2(n_222),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_599),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_565),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_606),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_609),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_630),
.Y(n_690)
);

INVx5_ASAP7_75t_L g691 ( 
.A(n_608),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_588),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_576),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_571),
.B(n_523),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_610),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_616),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_630),
.B(n_485),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_587),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_630),
.B(n_540),
.Y(n_699)
);

INVx4_ASAP7_75t_L g700 ( 
.A(n_576),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_620),
.Y(n_701)
);

OR2x6_ASAP7_75t_L g702 ( 
.A(n_563),
.B(n_493),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_584),
.A2(n_541),
.B1(n_543),
.B2(n_538),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_L g704 ( 
.A1(n_593),
.A2(n_506),
.B1(n_472),
.B2(n_355),
.Y(n_704)
);

OR2x6_ASAP7_75t_L g705 ( 
.A(n_563),
.B(n_640),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_587),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_621),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_636),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_622),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_632),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_619),
.B(n_544),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_572),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_629),
.B(n_545),
.Y(n_713)
);

NAND3xp33_ASAP7_75t_L g714 ( 
.A(n_591),
.B(n_549),
.C(n_550),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_576),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_594),
.Y(n_716)
);

BUFx6f_ASAP7_75t_SL g717 ( 
.A(n_595),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_572),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_573),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_608),
.B(n_364),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_573),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_581),
.B(n_592),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_608),
.A2(n_364),
.B1(n_395),
.B2(n_391),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_SL g724 ( 
.A(n_629),
.B(n_640),
.Y(n_724)
);

AO22x2_ASAP7_75t_L g725 ( 
.A1(n_581),
.A2(n_283),
.B1(n_314),
.B2(n_264),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_574),
.Y(n_726)
);

AND2x2_ASAP7_75t_SL g727 ( 
.A(n_581),
.B(n_283),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_578),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_608),
.B(n_275),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_580),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_608),
.B(n_345),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_551),
.B(n_492),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_592),
.B(n_245),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_578),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_589),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_594),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_589),
.Y(n_737)
);

OR2x6_ASAP7_75t_L g738 ( 
.A(n_637),
.B(n_508),
.Y(n_738)
);

AND2x2_ASAP7_75t_SL g739 ( 
.A(n_592),
.B(n_314),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_602),
.B(n_281),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_641),
.B(n_357),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_580),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_636),
.B(n_512),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_612),
.B(n_505),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_641),
.B(n_357),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_631),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_580),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_611),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_641),
.B(n_374),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_611),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_612),
.B(n_492),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_580),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_602),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_602),
.B(n_374),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_617),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_617),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_579),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_641),
.B(n_492),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_580),
.B(n_583),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_583),
.B(n_229),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_583),
.B(n_230),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_641),
.Y(n_762)
);

INVx4_ASAP7_75t_SL g763 ( 
.A(n_583),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_583),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_618),
.B(n_511),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_623),
.B(n_526),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_623),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_618),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_624),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_624),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_627),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_623),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_627),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_623),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_623),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_625),
.Y(n_776)
);

NOR2x1p5_ASAP7_75t_L g777 ( 
.A(n_579),
.B(n_236),
.Y(n_777)
);

BUFx10_ASAP7_75t_L g778 ( 
.A(n_552),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_625),
.B(n_231),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_625),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_625),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_625),
.B(n_633),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_633),
.B(n_243),
.Y(n_783)
);

AND2x6_ASAP7_75t_L g784 ( 
.A(n_633),
.B(n_252),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_633),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_633),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_588),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_553),
.Y(n_788)
);

NOR2x1p5_ASAP7_75t_L g789 ( 
.A(n_553),
.B(n_246),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_595),
.B(n_252),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_595),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_554),
.B(n_475),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_554),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_555),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_555),
.B(n_495),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_564),
.B(n_495),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_727),
.B(n_252),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_765),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_727),
.B(n_252),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_668),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_650),
.B(n_512),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_739),
.B(n_251),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_739),
.B(n_253),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_678),
.B(n_233),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_678),
.A2(n_381),
.B(n_380),
.C(n_378),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_646),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_670),
.Y(n_807)
);

NAND3xp33_ASAP7_75t_SL g808 ( 
.A(n_669),
.B(n_598),
.C(n_597),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_647),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_647),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_674),
.B(n_233),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_672),
.B(n_289),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_708),
.B(n_564),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_729),
.A2(n_262),
.B(n_258),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_708),
.A2(n_397),
.B(n_418),
.C(n_419),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_660),
.B(n_263),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_691),
.B(n_289),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_661),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_691),
.B(n_289),
.Y(n_819)
);

NOR3xp33_ASAP7_75t_L g820 ( 
.A(n_792),
.B(n_796),
.C(n_795),
.Y(n_820)
);

NOR2xp67_ASAP7_75t_L g821 ( 
.A(n_791),
.B(n_569),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_679),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_722),
.B(n_569),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_722),
.A2(n_668),
.B1(n_664),
.B2(n_694),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_664),
.A2(n_377),
.B1(n_239),
.B2(n_241),
.Y(n_825)
);

NAND2x1_ASAP7_75t_L g826 ( 
.A(n_643),
.B(n_507),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_743),
.A2(n_323),
.B(n_369),
.C(n_368),
.Y(n_827)
);

INVxp33_ASAP7_75t_L g828 ( 
.A(n_711),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_788),
.Y(n_829)
);

BUFx4f_ASAP7_75t_L g830 ( 
.A(n_705),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_691),
.B(n_731),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_649),
.B(n_266),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_744),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_656),
.B(n_712),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_664),
.A2(n_238),
.B1(n_239),
.B2(n_241),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_788),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_714),
.B(n_644),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_765),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_659),
.A2(n_277),
.B(n_273),
.Y(n_839)
);

BUFx5_ASAP7_75t_L g840 ( 
.A(n_784),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_744),
.A2(n_407),
.B(n_420),
.C(n_427),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_718),
.B(n_286),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_719),
.B(n_319),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_721),
.B(n_331),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_723),
.A2(n_425),
.B1(n_394),
.B2(n_373),
.Y(n_845)
);

NOR3xp33_ASAP7_75t_L g846 ( 
.A(n_685),
.B(n_598),
.C(n_597),
.Y(n_846)
);

OAI21xp33_ASAP7_75t_L g847 ( 
.A1(n_743),
.A2(n_433),
.B(n_517),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_726),
.Y(n_848)
);

OR2x6_ASAP7_75t_L g849 ( 
.A(n_705),
.B(n_547),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_691),
.B(n_289),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_691),
.B(n_327),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_743),
.B(n_577),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_728),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_664),
.A2(n_268),
.B1(n_238),
.B2(n_244),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_661),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_734),
.B(n_358),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_713),
.B(n_577),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_735),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_737),
.Y(n_859)
);

BUFx5_ASAP7_75t_L g860 ( 
.A(n_784),
.Y(n_860)
);

NAND2xp33_ASAP7_75t_L g861 ( 
.A(n_690),
.B(n_327),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_659),
.B(n_327),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_648),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_766),
.B(n_244),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_650),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_658),
.B(n_363),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_662),
.Y(n_867)
);

AND2x2_ASAP7_75t_SL g868 ( 
.A(n_720),
.B(n_327),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_671),
.B(n_372),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_676),
.B(n_376),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_725),
.A2(n_327),
.B1(n_337),
.B2(n_341),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_703),
.B(n_255),
.Y(n_872)
);

OR2x6_ASAP7_75t_L g873 ( 
.A(n_705),
.B(n_794),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_677),
.B(n_411),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_680),
.B(n_412),
.Y(n_875)
);

OAI22xp33_ASAP7_75t_L g876 ( 
.A1(n_733),
.A2(n_409),
.B1(n_254),
.B2(n_267),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_684),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_692),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_657),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_657),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_686),
.B(n_417),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_725),
.A2(n_337),
.B1(n_341),
.B2(n_352),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_725),
.A2(n_337),
.B1(n_341),
.B2(n_352),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_667),
.A2(n_428),
.B1(n_259),
.B2(n_261),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_688),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_689),
.B(n_337),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_738),
.B(n_705),
.Y(n_887)
);

NOR2x1p5_ASAP7_75t_L g888 ( 
.A(n_791),
.B(n_603),
.Y(n_888)
);

OR2x6_ASAP7_75t_L g889 ( 
.A(n_794),
.B(n_511),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_695),
.B(n_337),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_696),
.B(n_341),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_701),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_707),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_709),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_673),
.Y(n_895)
);

NAND2xp33_ASAP7_75t_L g896 ( 
.A(n_740),
.B(n_341),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_753),
.B(n_352),
.Y(n_897)
);

NOR3xp33_ASAP7_75t_L g898 ( 
.A(n_704),
.B(n_604),
.C(n_603),
.Y(n_898)
);

NAND2xp33_ASAP7_75t_L g899 ( 
.A(n_710),
.B(n_746),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_697),
.B(n_352),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_673),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_687),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_699),
.B(n_382),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_746),
.B(n_255),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_687),
.Y(n_905)
);

NAND2x1p5_ASAP7_75t_L g906 ( 
.A(n_675),
.B(n_382),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_762),
.B(n_382),
.Y(n_907)
);

O2A1O1Ixp5_ASAP7_75t_L g908 ( 
.A1(n_741),
.A2(n_525),
.B(n_546),
.C(n_537),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_775),
.B(n_382),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_698),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_776),
.B(n_259),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_653),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_738),
.B(n_604),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_655),
.A2(n_513),
.B(n_518),
.C(n_520),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_751),
.B(n_786),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_786),
.B(n_261),
.Y(n_916)
);

NAND2xp33_ASAP7_75t_L g917 ( 
.A(n_784),
.B(n_268),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_698),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_706),
.Y(n_919)
);

NOR2xp67_ASAP7_75t_L g920 ( 
.A(n_732),
.B(n_605),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_757),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_790),
.B(n_375),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_693),
.B(n_375),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_693),
.B(n_377),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_655),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_790),
.A2(n_528),
.B(n_513),
.C(n_518),
.Y(n_926)
);

BUFx12f_ASAP7_75t_SL g927 ( 
.A(n_738),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_738),
.B(n_379),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_681),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_675),
.B(n_392),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_716),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_754),
.A2(n_520),
.B(n_524),
.C(n_525),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_724),
.B(n_392),
.Y(n_933)
);

NAND2xp33_ASAP7_75t_L g934 ( 
.A(n_784),
.B(n_398),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_716),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_725),
.A2(n_247),
.B1(n_254),
.B2(n_267),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_747),
.B(n_772),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_789),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_759),
.B(n_399),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_736),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_736),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_782),
.B(n_400),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_702),
.B(n_404),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_787),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_748),
.Y(n_945)
);

BUFx8_ASAP7_75t_L g946 ( 
.A(n_717),
.Y(n_946)
);

AOI221xp5_ASAP7_75t_L g947 ( 
.A1(n_793),
.A2(n_247),
.B1(n_396),
.B2(n_269),
.C(n_270),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_702),
.A2(n_416),
.B1(n_404),
.B2(n_430),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_702),
.B(n_406),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_750),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_750),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_755),
.A2(n_421),
.B1(n_324),
.B2(n_328),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_755),
.B(n_406),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_756),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_880),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_834),
.B(n_816),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_864),
.B(n_832),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_864),
.B(n_772),
.Y(n_958)
);

AOI21x1_ASAP7_75t_L g959 ( 
.A1(n_831),
.A2(n_781),
.B(n_780),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_812),
.A2(n_799),
.B(n_797),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_837),
.A2(n_758),
.B(n_663),
.C(n_783),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_811),
.B(n_774),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_848),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_811),
.B(n_774),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_850),
.A2(n_645),
.B(n_643),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_802),
.A2(n_702),
.B1(n_601),
.B2(n_560),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_853),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_828),
.B(n_651),
.Y(n_968)
);

O2A1O1Ixp5_ASAP7_75t_L g969 ( 
.A1(n_812),
.A2(n_749),
.B(n_745),
.C(n_760),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_833),
.B(n_651),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_837),
.A2(n_761),
.B(n_779),
.C(n_757),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_937),
.A2(n_666),
.B(n_645),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_912),
.A2(n_700),
.B(n_666),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_803),
.A2(n_642),
.B1(n_605),
.B2(n_777),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_858),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_798),
.B(n_838),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_800),
.B(n_767),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_912),
.A2(n_700),
.B(n_666),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_800),
.B(n_774),
.Y(n_979)
);

BUFx4f_ASAP7_75t_L g980 ( 
.A(n_873),
.Y(n_980)
);

AO21x1_ASAP7_75t_L g981 ( 
.A1(n_797),
.A2(n_749),
.B(n_745),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_859),
.B(n_767),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_836),
.Y(n_983)
);

INVx5_ASAP7_75t_L g984 ( 
.A(n_929),
.Y(n_984)
);

NAND2xp33_ASAP7_75t_L g985 ( 
.A(n_840),
.B(n_653),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_929),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_807),
.B(n_626),
.Y(n_987)
);

AO21x1_ASAP7_75t_L g988 ( 
.A1(n_799),
.A2(n_730),
.B(n_715),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_813),
.B(n_651),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_804),
.B(n_785),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_804),
.B(n_785),
.Y(n_991)
);

CKINVDCx10_ASAP7_75t_R g992 ( 
.A(n_829),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_880),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_915),
.B(n_756),
.Y(n_994)
);

NAND2xp33_ASAP7_75t_SL g995 ( 
.A(n_888),
.B(n_717),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_925),
.A2(n_717),
.B1(n_652),
.B2(n_665),
.Y(n_996)
);

NOR2xp67_ASAP7_75t_L g997 ( 
.A(n_808),
.B(n_768),
.Y(n_997)
);

O2A1O1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_914),
.A2(n_768),
.B(n_773),
.C(n_771),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_822),
.B(n_769),
.Y(n_999)
);

AO21x1_ASAP7_75t_L g1000 ( 
.A1(n_814),
.A2(n_742),
.B(n_771),
.Y(n_1000)
);

OAI321xp33_ASAP7_75t_L g1001 ( 
.A1(n_876),
.A2(n_532),
.A3(n_529),
.B1(n_530),
.B2(n_534),
.C(n_546),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_815),
.A2(n_773),
.B(n_770),
.C(n_769),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_922),
.B(n_770),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_922),
.B(n_654),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_944),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_806),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_878),
.B(n_626),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_918),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_820),
.A2(n_652),
.B1(n_665),
.B2(n_683),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_872),
.A2(n_424),
.B(n_413),
.C(n_414),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_872),
.B(n_787),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_862),
.A2(n_654),
.B(n_764),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_863),
.B(n_877),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_862),
.A2(n_681),
.B(n_764),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_865),
.Y(n_1015)
);

NOR2x1p5_ASAP7_75t_L g1016 ( 
.A(n_921),
.B(n_652),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_900),
.A2(n_903),
.B(n_923),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_857),
.B(n_665),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_924),
.A2(n_681),
.B(n_764),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_841),
.A2(n_537),
.B(n_534),
.C(n_532),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_932),
.A2(n_529),
.B(n_500),
.C(n_498),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_879),
.B(n_763),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_946),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_801),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_885),
.B(n_681),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_845),
.A2(n_386),
.B1(n_384),
.B2(n_371),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_892),
.B(n_682),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_801),
.B(n_763),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_921),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_SL g1030 ( 
.A(n_830),
.B(n_683),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_904),
.A2(n_415),
.B(n_430),
.C(n_424),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_845),
.A2(n_408),
.B1(n_328),
.B2(n_324),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_889),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_932),
.A2(n_500),
.B(n_498),
.C(n_490),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_826),
.A2(n_752),
.B(n_763),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_871),
.A2(n_271),
.B1(n_431),
.B2(n_371),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_899),
.A2(n_763),
.B(n_413),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_916),
.A2(n_414),
.B(n_415),
.Y(n_1038)
);

NOR3xp33_ASAP7_75t_L g1039 ( 
.A(n_933),
.B(n_416),
.C(n_351),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_861),
.A2(n_784),
.B(n_429),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_873),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_893),
.B(n_683),
.Y(n_1042)
);

NOR2xp67_ASAP7_75t_L g1043 ( 
.A(n_938),
.B(n_84),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_894),
.B(n_784),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_824),
.B(n_778),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_907),
.A2(n_384),
.B(n_429),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_895),
.A2(n_386),
.B(n_426),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_904),
.B(n_389),
.Y(n_1048)
);

OAI321xp33_ASAP7_75t_L g1049 ( 
.A1(n_876),
.A2(n_426),
.A3(n_423),
.B1(n_421),
.B2(n_410),
.C(n_409),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_953),
.A2(n_423),
.B(n_410),
.C(n_408),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_943),
.A2(n_949),
.B(n_928),
.C(n_847),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_852),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_901),
.A2(n_389),
.B(n_405),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_943),
.A2(n_405),
.B(n_402),
.C(n_396),
.Y(n_1054)
);

OAI21xp33_ASAP7_75t_L g1055 ( 
.A1(n_950),
.A2(n_402),
.B(n_390),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_842),
.B(n_390),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_873),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_809),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_810),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_902),
.A2(n_153),
.B(n_205),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_821),
.B(n_778),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_953),
.A2(n_9),
.B(n_12),
.C(n_13),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_939),
.A2(n_778),
.B1(n_204),
.B2(n_198),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_905),
.A2(n_919),
.B(n_910),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_843),
.B(n_17),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_931),
.A2(n_940),
.B(n_935),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_941),
.A2(n_196),
.B(n_191),
.Y(n_1067)
);

O2A1O1Ixp5_ASAP7_75t_L g1068 ( 
.A1(n_939),
.A2(n_190),
.B(n_181),
.C(n_179),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_871),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_945),
.A2(n_819),
.B(n_851),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_817),
.A2(n_177),
.B(n_175),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_823),
.B(n_174),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_882),
.A2(n_166),
.B1(n_162),
.B2(n_150),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_817),
.A2(n_146),
.B(n_145),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_889),
.B(n_20),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_948),
.B(n_142),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_819),
.A2(n_128),
.B(n_122),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_933),
.B(n_22),
.Y(n_1078)
);

OAI321xp33_ASAP7_75t_L g1079 ( 
.A1(n_936),
.A2(n_22),
.A3(n_23),
.B1(n_24),
.B2(n_27),
.C(n_28),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_942),
.A2(n_117),
.B(n_101),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_882),
.A2(n_23),
.B1(n_30),
.B2(n_31),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_942),
.A2(n_99),
.B(n_92),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_818),
.A2(n_855),
.B(n_867),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_889),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_844),
.B(n_35),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_949),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_1086)
);

BUFx12f_ASAP7_75t_L g1087 ( 
.A(n_946),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_954),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_951),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_911),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_927),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_856),
.B(n_52),
.Y(n_1092)
);

OR2x6_ASAP7_75t_SL g1093 ( 
.A(n_884),
.B(n_54),
.Y(n_1093)
);

NOR3xp33_ASAP7_75t_L g1094 ( 
.A(n_846),
.B(n_55),
.C(n_56),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_908),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_830),
.B(n_61),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_849),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_911),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_1098)
);

AO22x1_ASAP7_75t_L g1099 ( 
.A1(n_928),
.A2(n_63),
.B1(n_67),
.B2(n_68),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_825),
.B(n_69),
.Y(n_1100)
);

BUFx12f_ASAP7_75t_L g1101 ( 
.A(n_849),
.Y(n_1101)
);

O2A1O1Ixp5_ASAP7_75t_L g1102 ( 
.A1(n_839),
.A2(n_874),
.B(n_866),
.C(n_869),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_926),
.A2(n_854),
.B(n_835),
.C(n_805),
.Y(n_1103)
);

INVxp33_ASAP7_75t_L g1104 ( 
.A(n_913),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_909),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_870),
.A2(n_77),
.B(n_74),
.C(n_75),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_849),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_920),
.B(n_73),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_868),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_887),
.B(n_77),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_875),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_881),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_868),
.B(n_883),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_886),
.A2(n_891),
.B(n_890),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_883),
.A2(n_936),
.B(n_930),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_909),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_950),
.A2(n_952),
.B1(n_947),
.B2(n_930),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_952),
.B(n_827),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_906),
.B(n_840),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_897),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_840),
.B(n_860),
.Y(n_1121)
);

O2A1O1Ixp5_ASAP7_75t_L g1122 ( 
.A1(n_897),
.A2(n_896),
.B(n_906),
.C(n_934),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_840),
.B(n_860),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_840),
.B(n_860),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_840),
.B(n_860),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_898),
.B(n_917),
.Y(n_1126)
);

INVx4_ASAP7_75t_SL g1127 ( 
.A(n_860),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_963),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_1011),
.B(n_956),
.Y(n_1129)
);

O2A1O1Ixp5_ASAP7_75t_L g1130 ( 
.A1(n_1000),
.A2(n_957),
.B(n_1017),
.C(n_960),
.Y(n_1130)
);

INVx5_ASAP7_75t_L g1131 ( 
.A(n_984),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_959),
.A2(n_972),
.B(n_1019),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1111),
.B(n_1112),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1078),
.A2(n_1051),
.B(n_1117),
.C(n_1115),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_1005),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1112),
.B(n_976),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1112),
.B(n_961),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_955),
.B(n_993),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1113),
.A2(n_969),
.B(n_971),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_1028),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1117),
.A2(n_1100),
.B(n_1079),
.C(n_1069),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_999),
.B(n_1048),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1118),
.A2(n_1126),
.B(n_1103),
.C(n_1010),
.Y(n_1143)
);

OAI22x1_ASAP7_75t_L g1144 ( 
.A1(n_1009),
.A2(n_1018),
.B1(n_1110),
.B2(n_996),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1004),
.A2(n_991),
.B(n_990),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_967),
.B(n_975),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_958),
.A2(n_964),
.B(n_962),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_987),
.B(n_1104),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1050),
.A2(n_997),
.B(n_1031),
.C(n_1039),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1013),
.B(n_994),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1079),
.A2(n_1069),
.B(n_1081),
.C(n_1001),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1003),
.B(n_1056),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_985),
.A2(n_965),
.B(n_1102),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1120),
.B(n_1008),
.Y(n_1154)
);

BUFx12f_ASAP7_75t_L g1155 ( 
.A(n_1087),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_989),
.B(n_1052),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1088),
.B(n_1089),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1081),
.A2(n_1001),
.B(n_1049),
.C(n_1109),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_981),
.A2(n_979),
.B(n_1114),
.Y(n_1159)
);

O2A1O1Ixp5_ASAP7_75t_L g1160 ( 
.A1(n_1122),
.A2(n_1092),
.B(n_1065),
.C(n_1085),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_998),
.A2(n_1070),
.B(n_1119),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1006),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_982),
.B(n_1042),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1028),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_1029),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_SL g1166 ( 
.A1(n_1086),
.A2(n_1026),
.B(n_1032),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1007),
.B(n_1075),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1049),
.A2(n_1062),
.B(n_1090),
.C(n_1098),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1058),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1110),
.B(n_1033),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1059),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_984),
.A2(n_1027),
.B(n_1025),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1106),
.A2(n_1095),
.A3(n_1073),
.B(n_1054),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1002),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_986),
.Y(n_1175)
);

NAND3xp33_ASAP7_75t_L g1176 ( 
.A(n_1026),
.B(n_1032),
.C(n_1094),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1015),
.B(n_1024),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_984),
.A2(n_973),
.B(n_978),
.Y(n_1178)
);

AND3x4_ASAP7_75t_L g1179 ( 
.A(n_1043),
.B(n_1022),
.C(n_1093),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_955),
.B(n_993),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_966),
.B(n_974),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_977),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_983),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1015),
.B(n_1024),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_986),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_980),
.A2(n_977),
.B1(n_984),
.B2(n_1045),
.Y(n_1186)
);

NAND2x1p5_ASAP7_75t_L g1187 ( 
.A(n_980),
.B(n_955),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1014),
.A2(n_1035),
.B(n_1012),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1024),
.B(n_968),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_993),
.B(n_1084),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_992),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1041),
.B(n_1057),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1123),
.A2(n_1124),
.B(n_1125),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1063),
.A2(n_1076),
.B(n_1072),
.C(n_1108),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1022),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1015),
.B(n_1055),
.Y(n_1196)
);

OAI22x1_ASAP7_75t_L g1197 ( 
.A1(n_1096),
.A2(n_1097),
.B1(n_1016),
.B2(n_1107),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1046),
.B(n_1038),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1084),
.B(n_1047),
.Y(n_1199)
);

INVx5_ASAP7_75t_L g1200 ( 
.A(n_1084),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1053),
.B(n_1036),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_1101),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1064),
.A2(n_1083),
.B(n_1066),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1020),
.A2(n_1068),
.B(n_1080),
.C(n_1082),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1036),
.B(n_1116),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1105),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1041),
.B(n_1057),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1030),
.B(n_1044),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1041),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1121),
.A2(n_1037),
.B(n_1071),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_970),
.A2(n_1060),
.B(n_1067),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_1057),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1074),
.A2(n_1077),
.B(n_1034),
.Y(n_1213)
);

INVx5_ASAP7_75t_L g1214 ( 
.A(n_1107),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1021),
.A2(n_1040),
.B(n_1061),
.Y(n_1215)
);

AOI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1099),
.A2(n_1127),
.B(n_1030),
.Y(n_1216)
);

NAND2x1p5_ASAP7_75t_L g1217 ( 
.A(n_1127),
.B(n_995),
.Y(n_1217)
);

OAI22x1_ASAP7_75t_L g1218 ( 
.A1(n_1091),
.A2(n_1011),
.B1(n_1100),
.B2(n_626),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1127),
.A2(n_959),
.B(n_972),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1023),
.A2(n_959),
.B(n_972),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_1000),
.A2(n_981),
.A3(n_988),
.B(n_971),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_1005),
.Y(n_1222)
);

NOR2xp67_ASAP7_75t_L g1223 ( 
.A(n_983),
.B(n_791),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_956),
.B(n_957),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1028),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_959),
.A2(n_972),
.B(n_1019),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_956),
.A2(n_1004),
.B(n_957),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_957),
.A2(n_1078),
.B(n_956),
.C(n_1011),
.Y(n_1228)
);

CKINVDCx11_ASAP7_75t_R g1229 ( 
.A(n_1087),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_955),
.B(n_880),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1011),
.B(n_828),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_956),
.B(n_957),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_956),
.B(n_957),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_1087),
.Y(n_1234)
);

NAND2xp33_ASAP7_75t_L g1235 ( 
.A(n_956),
.B(n_957),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_956),
.B(n_957),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1011),
.B(n_828),
.Y(n_1237)
);

AOI21x1_ASAP7_75t_SL g1238 ( 
.A1(n_1118),
.A2(n_1085),
.B(n_1065),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_963),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1011),
.B(n_828),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1005),
.Y(n_1241)
);

INVx4_ASAP7_75t_L g1242 ( 
.A(n_955),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_956),
.A2(n_1004),
.B(n_957),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_956),
.A2(n_1004),
.B(n_957),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_959),
.A2(n_972),
.B(n_1019),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_984),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1028),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1011),
.B(n_828),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_957),
.A2(n_1078),
.B(n_956),
.C(n_1011),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_956),
.B(n_957),
.Y(n_1250)
);

OAI22x1_ASAP7_75t_L g1251 ( 
.A1(n_1011),
.A2(n_1100),
.B1(n_626),
.B2(n_1009),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_956),
.B(n_957),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_959),
.A2(n_972),
.B(n_1019),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_956),
.B(n_957),
.Y(n_1254)
);

AOI211x1_ASAP7_75t_L g1255 ( 
.A1(n_1117),
.A2(n_1115),
.B(n_1069),
.C(n_1081),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1078),
.A2(n_1115),
.B(n_1117),
.C(n_1011),
.Y(n_1256)
);

NAND2x1p5_ASAP7_75t_L g1257 ( 
.A(n_984),
.B(n_1028),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_956),
.B(n_957),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_956),
.B(n_957),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_956),
.A2(n_1004),
.B(n_957),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_956),
.B(n_957),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_960),
.A2(n_957),
.B(n_1113),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1088),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_956),
.B(n_957),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_963),
.Y(n_1265)
);

NOR2xp67_ASAP7_75t_L g1266 ( 
.A(n_983),
.B(n_791),
.Y(n_1266)
);

NOR2x1_ASAP7_75t_SL g1267 ( 
.A(n_984),
.B(n_1069),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_956),
.B(n_957),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_956),
.B(n_957),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_959),
.A2(n_972),
.B(n_1019),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1005),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_992),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_959),
.A2(n_972),
.B(n_1019),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_963),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_956),
.B(n_957),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_959),
.A2(n_972),
.B(n_1019),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_956),
.B(n_957),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_956),
.B(n_957),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_963),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1128),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1190),
.B(n_1138),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1129),
.B(n_1224),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1239),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1240),
.B(n_1167),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1129),
.B(n_1232),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1138),
.B(n_1180),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1181),
.A2(n_1248),
.B1(n_1237),
.B2(n_1231),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1135),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1265),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1236),
.B(n_1250),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_SL g1291 ( 
.A(n_1141),
.B(n_1256),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1252),
.B(n_1254),
.Y(n_1292)
);

NOR2x1_ASAP7_75t_SL g1293 ( 
.A(n_1131),
.B(n_1246),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1180),
.B(n_1230),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1274),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1279),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1258),
.B(n_1278),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1146),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1181),
.A2(n_1176),
.B1(n_1251),
.B2(n_1218),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1259),
.B(n_1261),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1157),
.Y(n_1301)
);

NAND2xp33_ASAP7_75t_L g1302 ( 
.A(n_1228),
.B(n_1249),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1206),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1200),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1264),
.A2(n_1277),
.B1(n_1275),
.B2(n_1268),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1246),
.Y(n_1306)
);

AO21x1_ASAP7_75t_L g1307 ( 
.A1(n_1227),
.A2(n_1244),
.B(n_1243),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1263),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1200),
.Y(n_1309)
);

NOR2xp67_ASAP7_75t_L g1310 ( 
.A(n_1131),
.B(n_1142),
.Y(n_1310)
);

OA21x2_ASAP7_75t_L g1311 ( 
.A1(n_1139),
.A2(n_1130),
.B(n_1159),
.Y(n_1311)
);

OAI21xp33_ASAP7_75t_L g1312 ( 
.A1(n_1256),
.A2(n_1141),
.B(n_1166),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1260),
.A2(n_1153),
.B(n_1235),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1191),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1156),
.B(n_1231),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1237),
.B(n_1248),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1134),
.A2(n_1143),
.B(n_1130),
.Y(n_1317)
);

INVx6_ASAP7_75t_L g1318 ( 
.A(n_1200),
.Y(n_1318)
);

O2A1O1Ixp5_ASAP7_75t_L g1319 ( 
.A1(n_1194),
.A2(n_1160),
.B(n_1168),
.C(n_1151),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1135),
.B(n_1241),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1200),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1230),
.B(n_1192),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_R g1323 ( 
.A(n_1272),
.B(n_1222),
.Y(n_1323)
);

INVx1_ASAP7_75t_SL g1324 ( 
.A(n_1241),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1229),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1233),
.B(n_1269),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1271),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1170),
.B(n_1148),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1165),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1183),
.Y(n_1330)
);

INVx5_ASAP7_75t_L g1331 ( 
.A(n_1246),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1171),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1246),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1148),
.B(n_1136),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1233),
.B(n_1269),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1162),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1131),
.Y(n_1337)
);

INVx5_ASAP7_75t_L g1338 ( 
.A(n_1131),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1169),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1133),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_SL g1341 ( 
.A(n_1151),
.B(n_1158),
.Y(n_1341)
);

NAND2x1p5_ASAP7_75t_L g1342 ( 
.A(n_1242),
.B(n_1214),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1150),
.B(n_1152),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1154),
.B(n_1196),
.Y(n_1344)
);

AND2x6_ASAP7_75t_L g1345 ( 
.A(n_1140),
.B(n_1164),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1260),
.B(n_1163),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1223),
.B(n_1266),
.Y(n_1347)
);

OR2x6_ASAP7_75t_L g1348 ( 
.A(n_1187),
.B(n_1257),
.Y(n_1348)
);

NAND3xp33_ASAP7_75t_L g1349 ( 
.A(n_1255),
.B(n_1168),
.C(n_1158),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1192),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1179),
.B(n_1177),
.Y(n_1351)
);

INVx4_ASAP7_75t_L g1352 ( 
.A(n_1214),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_SL g1353 ( 
.A1(n_1210),
.A2(n_1262),
.B(n_1211),
.C(n_1145),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1175),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1189),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1147),
.A2(n_1159),
.B(n_1178),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1195),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1257),
.Y(n_1358)
);

AOI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1179),
.A2(n_1201),
.B1(n_1144),
.B2(n_1137),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1185),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_SL g1361 ( 
.A(n_1242),
.B(n_1187),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1199),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1149),
.B(n_1137),
.C(n_1160),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1147),
.A2(n_1178),
.B(n_1161),
.Y(n_1364)
);

NOR2xp67_ASAP7_75t_L g1365 ( 
.A(n_1140),
.B(n_1164),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1184),
.B(n_1205),
.Y(n_1366)
);

NAND2x1p5_ASAP7_75t_L g1367 ( 
.A(n_1214),
.B(n_1225),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1193),
.A2(n_1204),
.B(n_1211),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1174),
.A2(n_1193),
.B(n_1204),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1207),
.Y(n_1370)
);

CKINVDCx11_ASAP7_75t_R g1371 ( 
.A(n_1155),
.Y(n_1371)
);

INVxp67_ASAP7_75t_SL g1372 ( 
.A(n_1225),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1207),
.B(n_1247),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1209),
.B(n_1212),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1247),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1186),
.A2(n_1208),
.B1(n_1214),
.B2(n_1198),
.Y(n_1376)
);

OR2x6_ASAP7_75t_L g1377 ( 
.A(n_1202),
.B(n_1217),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1209),
.Y(n_1378)
);

OA21x2_ASAP7_75t_L g1379 ( 
.A1(n_1132),
.A2(n_1276),
.B(n_1273),
.Y(n_1379)
);

NAND2x1p5_ASAP7_75t_L g1380 ( 
.A(n_1182),
.B(n_1220),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1197),
.B(n_1173),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1173),
.Y(n_1382)
);

AND2x6_ASAP7_75t_L g1383 ( 
.A(n_1267),
.B(n_1216),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1217),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1172),
.A2(n_1219),
.B(n_1203),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_1234),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1221),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1173),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1215),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1188),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1213),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1226),
.A2(n_1245),
.B(n_1253),
.C(n_1270),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1238),
.Y(n_1393)
);

NOR2xp67_ASAP7_75t_SL g1394 ( 
.A(n_1221),
.B(n_1131),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1221),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1221),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1129),
.A2(n_1232),
.B1(n_1236),
.B2(n_1224),
.Y(n_1397)
);

OR2x6_ASAP7_75t_L g1398 ( 
.A(n_1187),
.B(n_1133),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1240),
.B(n_1167),
.Y(n_1399)
);

AOI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1129),
.A2(n_1011),
.B1(n_1032),
.B2(n_1026),
.C(n_1117),
.Y(n_1400)
);

BUFx4_ASAP7_75t_SL g1401 ( 
.A(n_1191),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1191),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_1135),
.Y(n_1403)
);

INVx5_ASAP7_75t_L g1404 ( 
.A(n_1246),
.Y(n_1404)
);

AOI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1129),
.A2(n_1166),
.B1(n_1176),
.B2(n_1117),
.Y(n_1405)
);

INVx4_ASAP7_75t_L g1406 ( 
.A(n_1131),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1181),
.A2(n_1176),
.B1(n_1129),
.B2(n_1011),
.Y(n_1407)
);

AO32x1_ASAP7_75t_L g1408 ( 
.A1(n_1174),
.A2(n_1069),
.A3(n_1081),
.B1(n_1117),
.B2(n_1073),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1129),
.B(n_1224),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1139),
.A2(n_1130),
.B(n_1159),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1128),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1246),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1246),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1128),
.Y(n_1414)
);

BUFx2_ASAP7_75t_SL g1415 ( 
.A(n_1200),
.Y(n_1415)
);

INVxp67_ASAP7_75t_L g1416 ( 
.A(n_1135),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1240),
.B(n_724),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1141),
.A2(n_1129),
.B1(n_1151),
.B2(n_1224),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1181),
.A2(n_1176),
.B1(n_1129),
.B2(n_1011),
.Y(n_1419)
);

O2A1O1Ixp33_ASAP7_75t_SL g1420 ( 
.A1(n_1256),
.A2(n_1141),
.B(n_1134),
.C(n_1151),
.Y(n_1420)
);

BUFx2_ASAP7_75t_SL g1421 ( 
.A(n_1200),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1240),
.B(n_1167),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1231),
.B(n_1237),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1190),
.B(n_1138),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1129),
.A2(n_1166),
.B1(n_1176),
.B2(n_1117),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1128),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1129),
.A2(n_1232),
.B1(n_1236),
.B2(n_1224),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_1135),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1240),
.B(n_1167),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1128),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1134),
.A2(n_1256),
.B(n_1143),
.Y(n_1431)
);

INVx5_ASAP7_75t_L g1432 ( 
.A(n_1246),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1200),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1240),
.B(n_1167),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1135),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1129),
.B(n_1224),
.Y(n_1436)
);

NOR2x1_ASAP7_75t_L g1437 ( 
.A(n_1183),
.B(n_921),
.Y(n_1437)
);

OAI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1129),
.A2(n_724),
.B1(n_1011),
.B2(n_1224),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1128),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1318),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1405),
.B(n_1425),
.Y(n_1441)
);

CKINVDCx11_ASAP7_75t_R g1442 ( 
.A(n_1325),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1405),
.B(n_1425),
.Y(n_1443)
);

AO21x2_ASAP7_75t_L g1444 ( 
.A1(n_1385),
.A2(n_1364),
.B(n_1392),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1400),
.A2(n_1419),
.B1(n_1407),
.B2(n_1312),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1312),
.A2(n_1299),
.B1(n_1291),
.B2(n_1287),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1283),
.Y(n_1447)
);

NAND2x1p5_ASAP7_75t_L g1448 ( 
.A(n_1394),
.B(n_1384),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1289),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1318),
.Y(n_1450)
);

OAI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1438),
.A2(n_1427),
.B(n_1397),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1282),
.B(n_1285),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1320),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1338),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1338),
.Y(n_1455)
);

CKINVDCx11_ASAP7_75t_R g1456 ( 
.A(n_1371),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1409),
.B(n_1436),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1292),
.A2(n_1297),
.B1(n_1300),
.B2(n_1343),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1414),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1291),
.A2(n_1341),
.B1(n_1349),
.B2(n_1423),
.Y(n_1460)
);

NAND2x1p5_ASAP7_75t_L g1461 ( 
.A(n_1384),
.B(n_1338),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1305),
.B(n_1334),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1280),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1295),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1296),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1288),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1411),
.Y(n_1467)
);

INVx6_ASAP7_75t_L g1468 ( 
.A(n_1331),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1426),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1341),
.A2(n_1349),
.B1(n_1302),
.B2(n_1417),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1418),
.A2(n_1431),
.B1(n_1344),
.B2(n_1351),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1304),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1304),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1322),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1322),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1430),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1324),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1324),
.Y(n_1478)
);

BUFx2_ASAP7_75t_SL g1479 ( 
.A(n_1331),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1316),
.A2(n_1434),
.B1(n_1284),
.B2(n_1422),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1439),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1382),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_SL g1483 ( 
.A1(n_1418),
.A2(n_1431),
.B1(n_1317),
.B2(n_1355),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1406),
.Y(n_1484)
);

AO21x2_ASAP7_75t_L g1485 ( 
.A1(n_1369),
.A2(n_1353),
.B(n_1317),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1403),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1359),
.A2(n_1429),
.B1(n_1399),
.B2(n_1362),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1336),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1294),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1359),
.B(n_1366),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1339),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1328),
.A2(n_1315),
.B1(n_1290),
.B2(n_1381),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1303),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1326),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1379),
.A2(n_1319),
.B(n_1380),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1355),
.A2(n_1335),
.B1(n_1388),
.B2(n_1363),
.Y(n_1496)
);

CKINVDCx11_ASAP7_75t_R g1497 ( 
.A(n_1386),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1307),
.A2(n_1346),
.B(n_1376),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1308),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1363),
.A2(n_1298),
.B1(n_1329),
.B2(n_1301),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1393),
.Y(n_1501)
);

CKINVDCx20_ASAP7_75t_R g1502 ( 
.A(n_1314),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1393),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_SL g1504 ( 
.A1(n_1340),
.A2(n_1361),
.B1(n_1383),
.B2(n_1330),
.Y(n_1504)
);

CKINVDCx11_ASAP7_75t_R g1505 ( 
.A(n_1401),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1311),
.A2(n_1410),
.B(n_1387),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1354),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_SL g1508 ( 
.A1(n_1361),
.A2(n_1383),
.B1(n_1403),
.B2(n_1428),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1281),
.B(n_1424),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1428),
.A2(n_1398),
.B1(n_1416),
.B2(n_1377),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1309),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1383),
.A2(n_1421),
.B1(n_1415),
.B2(n_1377),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1383),
.A2(n_1377),
.B1(n_1384),
.B2(n_1435),
.Y(n_1513)
);

AOI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1389),
.A2(n_1410),
.B(n_1311),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1360),
.Y(n_1515)
);

NAND2x1p5_ASAP7_75t_L g1516 ( 
.A(n_1352),
.B(n_1310),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1398),
.A2(n_1370),
.B1(n_1437),
.B2(n_1310),
.Y(n_1517)
);

BUFx4f_ASAP7_75t_SL g1518 ( 
.A(n_1350),
.Y(n_1518)
);

INVx3_ASAP7_75t_L g1519 ( 
.A(n_1345),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1345),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1398),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1347),
.B(n_1365),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1332),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1281),
.B(n_1424),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_SL g1525 ( 
.A1(n_1293),
.A2(n_1420),
.B1(n_1323),
.B2(n_1408),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1294),
.B(n_1373),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1378),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_SL g1528 ( 
.A1(n_1395),
.A2(n_1396),
.B(n_1352),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1357),
.B(n_1286),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1372),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1374),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1367),
.A2(n_1337),
.B(n_1342),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1375),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1375),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1286),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1306),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1348),
.B(n_1365),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1327),
.B(n_1350),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1309),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1350),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1345),
.A2(n_1348),
.B1(n_1358),
.B2(n_1391),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1309),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_SL g1543 ( 
.A1(n_1408),
.A2(n_1345),
.B1(n_1433),
.B2(n_1321),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1348),
.B(n_1358),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1402),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1390),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1391),
.A2(n_1390),
.B1(n_1412),
.B2(n_1333),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1412),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_SL g1549 ( 
.A1(n_1408),
.A2(n_1433),
.B1(n_1321),
.B2(n_1404),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1413),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1433),
.A2(n_1331),
.B1(n_1404),
.B2(n_1432),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1432),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1432),
.A2(n_1129),
.B1(n_1011),
.B2(n_1407),
.Y(n_1553)
);

OA21x2_ASAP7_75t_L g1554 ( 
.A1(n_1404),
.A2(n_1356),
.B(n_1368),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1413),
.B(n_1129),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_SL g1556 ( 
.A1(n_1291),
.A2(n_1011),
.B1(n_1181),
.B2(n_1129),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1338),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1407),
.A2(n_1129),
.B1(n_1011),
.B2(n_1419),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1283),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1299),
.A2(n_1011),
.B(n_626),
.Y(n_1560)
);

AOI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1400),
.A2(n_1011),
.B1(n_987),
.B2(n_553),
.Y(n_1561)
);

OAI22xp33_ASAP7_75t_R g1562 ( 
.A1(n_1423),
.A2(n_1011),
.B1(n_1237),
.B2(n_1231),
.Y(n_1562)
);

CKINVDCx11_ASAP7_75t_R g1563 ( 
.A(n_1325),
.Y(n_1563)
);

CKINVDCx11_ASAP7_75t_R g1564 ( 
.A(n_1325),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1318),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1282),
.B(n_1129),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1338),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1288),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1320),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1320),
.Y(n_1570)
);

INVx6_ASAP7_75t_L g1571 ( 
.A(n_1338),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1283),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1283),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1282),
.B(n_1129),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1283),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1281),
.B(n_1424),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1356),
.A2(n_1368),
.B(n_1313),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1338),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1400),
.A2(n_1011),
.B1(n_1181),
.B2(n_1176),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_SL g1580 ( 
.A1(n_1291),
.A2(n_1011),
.B1(n_1181),
.B2(n_1129),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1283),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1320),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1407),
.A2(n_1129),
.B1(n_1011),
.B2(n_1419),
.Y(n_1583)
);

OA21x2_ASAP7_75t_L g1584 ( 
.A1(n_1356),
.A2(n_1368),
.B(n_1313),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1283),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1288),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1338),
.Y(n_1587)
);

AO21x1_ASAP7_75t_SL g1588 ( 
.A1(n_1431),
.A2(n_1359),
.B(n_1312),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1401),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1320),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1423),
.B(n_828),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1283),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1405),
.B(n_1425),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1441),
.B(n_1443),
.Y(n_1594)
);

BUFx12f_ASAP7_75t_L g1595 ( 
.A(n_1505),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1477),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1441),
.B(n_1443),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1477),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1558),
.A2(n_1583),
.B1(n_1579),
.B2(n_1556),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1482),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1482),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1593),
.B(n_1588),
.Y(n_1602)
);

OR2x6_ASAP7_75t_L g1603 ( 
.A(n_1554),
.B(n_1498),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1591),
.B(n_1561),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1506),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1580),
.B(n_1458),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1490),
.B(n_1451),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1478),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1494),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1490),
.B(n_1494),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1486),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1485),
.B(n_1471),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1566),
.B(n_1574),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1546),
.B(n_1537),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1568),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1446),
.A2(n_1460),
.B1(n_1445),
.B2(n_1560),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1521),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1568),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1485),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1485),
.Y(n_1620)
);

NAND2x1p5_ASAP7_75t_L g1621 ( 
.A(n_1554),
.B(n_1519),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1514),
.Y(n_1622)
);

OA21x2_ASAP7_75t_L g1623 ( 
.A1(n_1495),
.A2(n_1528),
.B(n_1462),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1554),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1528),
.Y(n_1625)
);

INVxp67_ASAP7_75t_SL g1626 ( 
.A(n_1453),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1569),
.Y(n_1627)
);

BUFx2_ASAP7_75t_L g1628 ( 
.A(n_1521),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1570),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1582),
.B(n_1590),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1562),
.A2(n_1553),
.B1(n_1470),
.B2(n_1487),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1586),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1463),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1527),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1483),
.B(n_1449),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1562),
.A2(n_1492),
.B1(n_1525),
.B2(n_1504),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1530),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1527),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1464),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1530),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1465),
.Y(n_1641)
);

INVx4_ASAP7_75t_SL g1642 ( 
.A(n_1571),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1537),
.B(n_1544),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1467),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1469),
.Y(n_1645)
);

OAI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1577),
.A2(n_1584),
.B(n_1448),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1510),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1452),
.B(n_1457),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1476),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1448),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1466),
.Y(n_1651)
);

AO21x2_ASAP7_75t_L g1652 ( 
.A1(n_1444),
.A2(n_1522),
.B(n_1501),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1555),
.B(n_1500),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1481),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1480),
.B(n_1531),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1448),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1507),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1515),
.Y(n_1658)
);

AO21x2_ASAP7_75t_L g1659 ( 
.A1(n_1501),
.A2(n_1503),
.B(n_1488),
.Y(n_1659)
);

NAND3xp33_ASAP7_75t_L g1660 ( 
.A(n_1496),
.B(n_1517),
.C(n_1508),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1491),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1519),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1493),
.Y(n_1663)
);

BUFx4f_ASAP7_75t_SL g1664 ( 
.A(n_1502),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1447),
.Y(n_1665)
);

AO21x1_ASAP7_75t_SL g1666 ( 
.A1(n_1541),
.A2(n_1547),
.B(n_1550),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1499),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1459),
.B(n_1559),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1520),
.Y(n_1669)
);

BUFx6f_ASAP7_75t_L g1670 ( 
.A(n_1520),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1592),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1549),
.B(n_1529),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1572),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1573),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1516),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1544),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1575),
.Y(n_1677)
);

BUFx6f_ASAP7_75t_L g1678 ( 
.A(n_1544),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1571),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1581),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1516),
.A2(n_1532),
.B(n_1526),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1585),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1523),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1543),
.Y(n_1684)
);

INVx3_ASAP7_75t_L g1685 ( 
.A(n_1455),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1529),
.B(n_1524),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1533),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1534),
.B(n_1509),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1536),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1571),
.Y(n_1690)
);

AO21x2_ASAP7_75t_L g1691 ( 
.A1(n_1548),
.A2(n_1538),
.B(n_1540),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1454),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1454),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1509),
.B(n_1524),
.Y(n_1694)
);

BUFx3_ASAP7_75t_L g1695 ( 
.A(n_1571),
.Y(n_1695)
);

INVx2_ASAP7_75t_SL g1696 ( 
.A(n_1468),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1576),
.B(n_1474),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1567),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1576),
.B(n_1475),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1567),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1455),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1567),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1576),
.B(n_1474),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1475),
.B(n_1489),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1578),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1578),
.Y(n_1706)
);

NOR2x1_ASAP7_75t_SL g1707 ( 
.A(n_1479),
.B(n_1557),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1600),
.B(n_1513),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1607),
.B(n_1512),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1607),
.B(n_1578),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1605),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1612),
.B(n_1489),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1605),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1637),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1612),
.B(n_1484),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1619),
.B(n_1484),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1627),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1602),
.B(n_1484),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1637),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1610),
.B(n_1535),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1599),
.A2(n_1497),
.B1(n_1442),
.B2(n_1563),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1610),
.B(n_1473),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1594),
.B(n_1473),
.Y(n_1723)
);

NAND2x1p5_ASAP7_75t_L g1724 ( 
.A(n_1624),
.B(n_1557),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1616),
.A2(n_1606),
.B1(n_1604),
.B2(n_1631),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1620),
.B(n_1450),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1650),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1597),
.B(n_1557),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1640),
.B(n_1626),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1633),
.B(n_1473),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1614),
.B(n_1557),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1620),
.B(n_1450),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1630),
.B(n_1601),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1601),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_SL g1735 ( 
.A1(n_1660),
.A2(n_1552),
.B1(n_1479),
.B2(n_1468),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1609),
.B(n_1557),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1630),
.B(n_1565),
.Y(n_1737)
);

BUFx3_ASAP7_75t_L g1738 ( 
.A(n_1650),
.Y(n_1738)
);

OAI31xp33_ASAP7_75t_SL g1739 ( 
.A1(n_1684),
.A2(n_1551),
.A3(n_1552),
.B(n_1456),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1631),
.A2(n_1468),
.B1(n_1461),
.B2(n_1455),
.Y(n_1740)
);

NOR2x1p5_ASAP7_75t_L g1741 ( 
.A(n_1653),
.B(n_1587),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1614),
.B(n_1455),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1628),
.B(n_1565),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1659),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1659),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1628),
.B(n_1461),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1596),
.B(n_1461),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1639),
.B(n_1472),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1639),
.B(n_1472),
.Y(n_1749)
);

INVx2_ASAP7_75t_SL g1750 ( 
.A(n_1617),
.Y(n_1750)
);

OAI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1636),
.A2(n_1440),
.B1(n_1468),
.B2(n_1545),
.C(n_1542),
.Y(n_1751)
);

INVx4_ASAP7_75t_R g1752 ( 
.A(n_1679),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1691),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1641),
.B(n_1511),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1598),
.B(n_1440),
.Y(n_1755)
);

OAI211xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1613),
.A2(n_1442),
.B(n_1564),
.C(n_1563),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1644),
.Y(n_1757)
);

INVx3_ASAP7_75t_SL g1758 ( 
.A(n_1642),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1644),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1652),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1621),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1647),
.A2(n_1497),
.B1(n_1564),
.B2(n_1456),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1645),
.B(n_1472),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1645),
.B(n_1472),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1649),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1603),
.B(n_1472),
.Y(n_1766)
);

OAI21xp33_ASAP7_75t_SL g1767 ( 
.A1(n_1635),
.A2(n_1587),
.B(n_1539),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1649),
.Y(n_1768)
);

INVx3_ASAP7_75t_L g1769 ( 
.A(n_1621),
.Y(n_1769)
);

NOR3xp33_ASAP7_75t_L g1770 ( 
.A(n_1751),
.B(n_1681),
.C(n_1648),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1715),
.B(n_1623),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1729),
.B(n_1629),
.Y(n_1772)
);

NAND3xp33_ASAP7_75t_SL g1773 ( 
.A(n_1725),
.B(n_1655),
.C(n_1704),
.Y(n_1773)
);

OAI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1739),
.A2(n_1651),
.B1(n_1611),
.B2(n_1618),
.C(n_1632),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1729),
.B(n_1615),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1717),
.B(n_1634),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1715),
.B(n_1623),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_L g1778 ( 
.A(n_1735),
.B(n_1635),
.C(n_1706),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1751),
.A2(n_1643),
.B1(n_1684),
.B2(n_1676),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1715),
.B(n_1623),
.Y(n_1780)
);

OAI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1735),
.A2(n_1686),
.B1(n_1704),
.B2(n_1650),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1710),
.B(n_1638),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1712),
.B(n_1621),
.Y(n_1783)
);

NAND3xp33_ASAP7_75t_L g1784 ( 
.A(n_1739),
.B(n_1698),
.C(n_1706),
.Y(n_1784)
);

NOR3xp33_ASAP7_75t_L g1785 ( 
.A(n_1756),
.B(n_1675),
.C(n_1685),
.Y(n_1785)
);

NOR3xp33_ASAP7_75t_L g1786 ( 
.A(n_1756),
.B(n_1675),
.C(n_1685),
.Y(n_1786)
);

AOI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1721),
.A2(n_1611),
.B1(n_1608),
.B2(n_1688),
.C(n_1671),
.Y(n_1787)
);

NAND3xp33_ASAP7_75t_L g1788 ( 
.A(n_1740),
.B(n_1698),
.C(n_1705),
.Y(n_1788)
);

NAND3xp33_ASAP7_75t_L g1789 ( 
.A(n_1740),
.B(n_1693),
.C(n_1705),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1710),
.B(n_1608),
.Y(n_1790)
);

OAI221xp5_ASAP7_75t_SL g1791 ( 
.A1(n_1767),
.A2(n_1603),
.B1(n_1672),
.B2(n_1668),
.C(n_1694),
.Y(n_1791)
);

OAI221xp5_ASAP7_75t_SL g1792 ( 
.A1(n_1767),
.A2(n_1603),
.B1(n_1672),
.B2(n_1668),
.C(n_1694),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1733),
.B(n_1658),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1741),
.A2(n_1643),
.B1(n_1676),
.B2(n_1678),
.Y(n_1794)
);

NAND3xp33_ASAP7_75t_L g1795 ( 
.A(n_1709),
.B(n_1692),
.C(n_1702),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1712),
.B(n_1652),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1709),
.B(n_1675),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1766),
.B(n_1624),
.Y(n_1798)
);

NAND2x1p5_ASAP7_75t_L g1799 ( 
.A(n_1769),
.B(n_1624),
.Y(n_1799)
);

NAND3xp33_ASAP7_75t_L g1800 ( 
.A(n_1760),
.B(n_1702),
.C(n_1693),
.Y(n_1800)
);

AOI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1737),
.A2(n_1688),
.B1(n_1680),
.B2(n_1674),
.C(n_1677),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1733),
.B(n_1658),
.Y(n_1802)
);

NAND3xp33_ASAP7_75t_L g1803 ( 
.A(n_1747),
.B(n_1732),
.C(n_1726),
.Y(n_1803)
);

OAI21xp5_ASAP7_75t_SL g1804 ( 
.A1(n_1762),
.A2(n_1643),
.B(n_1703),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_SL g1805 ( 
.A1(n_1766),
.A2(n_1707),
.B1(n_1656),
.B2(n_1643),
.Y(n_1805)
);

OAI221xp5_ASAP7_75t_SL g1806 ( 
.A1(n_1708),
.A2(n_1603),
.B1(n_1656),
.B2(n_1673),
.C(n_1671),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1734),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1766),
.B(n_1624),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1737),
.B(n_1661),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1722),
.B(n_1603),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1730),
.B(n_1748),
.Y(n_1811)
);

OAI221xp5_ASAP7_75t_SL g1812 ( 
.A1(n_1708),
.A2(n_1656),
.B1(n_1677),
.B2(n_1680),
.C(n_1674),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1716),
.B(n_1723),
.Y(n_1813)
);

NAND3xp33_ASAP7_75t_L g1814 ( 
.A(n_1747),
.B(n_1692),
.C(n_1700),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1741),
.A2(n_1664),
.B1(n_1678),
.B2(n_1679),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_SL g1816 ( 
.A1(n_1728),
.A2(n_1703),
.B(n_1699),
.Y(n_1816)
);

NAND3xp33_ASAP7_75t_L g1817 ( 
.A(n_1726),
.B(n_1700),
.C(n_1625),
.Y(n_1817)
);

OAI21xp33_ASAP7_75t_L g1818 ( 
.A1(n_1728),
.A2(n_1753),
.B(n_1748),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1716),
.B(n_1625),
.Y(n_1819)
);

OAI221xp5_ASAP7_75t_L g1820 ( 
.A1(n_1755),
.A2(n_1675),
.B1(n_1696),
.B2(n_1695),
.C(n_1690),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1755),
.B(n_1678),
.Y(n_1821)
);

OAI21xp5_ASAP7_75t_SL g1822 ( 
.A1(n_1731),
.A2(n_1697),
.B(n_1699),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1731),
.A2(n_1678),
.B1(n_1666),
.B2(n_1595),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1749),
.B(n_1691),
.Y(n_1824)
);

OAI221xp5_ASAP7_75t_SL g1825 ( 
.A1(n_1743),
.A2(n_1673),
.B1(n_1657),
.B2(n_1654),
.C(n_1663),
.Y(n_1825)
);

NAND3xp33_ASAP7_75t_L g1826 ( 
.A(n_1732),
.B(n_1753),
.C(n_1743),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1749),
.B(n_1691),
.Y(n_1827)
);

OA21x2_ASAP7_75t_L g1828 ( 
.A1(n_1744),
.A2(n_1646),
.B(n_1622),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_L g1829 ( 
.A(n_1720),
.B(n_1595),
.Y(n_1829)
);

OAI221xp5_ASAP7_75t_SL g1830 ( 
.A1(n_1746),
.A2(n_1657),
.B1(n_1663),
.B2(n_1667),
.C(n_1683),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1731),
.A2(n_1666),
.B1(n_1697),
.B2(n_1695),
.Y(n_1831)
);

OAI221xp5_ASAP7_75t_SL g1832 ( 
.A1(n_1746),
.A2(n_1667),
.B1(n_1683),
.B2(n_1687),
.C(n_1682),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1731),
.A2(n_1670),
.B1(n_1662),
.B2(n_1669),
.Y(n_1833)
);

NAND2xp33_ASAP7_75t_SL g1834 ( 
.A(n_1758),
.B(n_1589),
.Y(n_1834)
);

OAI21xp5_ASAP7_75t_SL g1835 ( 
.A1(n_1742),
.A2(n_1696),
.B(n_1701),
.Y(n_1835)
);

AOI221xp5_ASAP7_75t_L g1836 ( 
.A1(n_1714),
.A2(n_1687),
.B1(n_1689),
.B2(n_1682),
.C(n_1665),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1807),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1798),
.B(n_1769),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1819),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1798),
.B(n_1761),
.Y(n_1840)
);

INVx3_ASAP7_75t_L g1841 ( 
.A(n_1799),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1808),
.B(n_1813),
.Y(n_1842)
);

INVx3_ASAP7_75t_L g1843 ( 
.A(n_1799),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1819),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1793),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1824),
.B(n_1714),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1828),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1775),
.B(n_1719),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1772),
.B(n_1719),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1802),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1813),
.B(n_1769),
.Y(n_1851)
);

BUFx2_ASAP7_75t_L g1852 ( 
.A(n_1810),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1809),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1827),
.B(n_1753),
.Y(n_1854)
);

AND2x4_ASAP7_75t_L g1855 ( 
.A(n_1810),
.B(n_1769),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1803),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1790),
.B(n_1745),
.Y(n_1857)
);

INVxp67_ASAP7_75t_SL g1858 ( 
.A(n_1797),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1782),
.B(n_1754),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1826),
.Y(n_1860)
);

NOR2xp67_ASAP7_75t_L g1861 ( 
.A(n_1817),
.B(n_1745),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1828),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1828),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1800),
.Y(n_1864)
);

NAND3xp33_ASAP7_75t_L g1865 ( 
.A(n_1770),
.B(n_1736),
.C(n_1665),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1814),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1771),
.B(n_1711),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1771),
.Y(n_1868)
);

INVx1_ASAP7_75t_SL g1869 ( 
.A(n_1776),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1783),
.B(n_1727),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1796),
.B(n_1783),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1777),
.B(n_1711),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1780),
.Y(n_1873)
);

NAND2x1p5_ASAP7_75t_L g1874 ( 
.A(n_1821),
.B(n_1750),
.Y(n_1874)
);

INVx1_ASAP7_75t_SL g1875 ( 
.A(n_1811),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1821),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1818),
.B(n_1750),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1799),
.B(n_1718),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1797),
.B(n_1711),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1795),
.B(n_1713),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1837),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1856),
.B(n_1806),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1852),
.B(n_1727),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1837),
.Y(n_1884)
);

INVx1_ASAP7_75t_SL g1885 ( 
.A(n_1869),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1847),
.Y(n_1886)
);

INVxp33_ASAP7_75t_L g1887 ( 
.A(n_1859),
.Y(n_1887)
);

AOI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1856),
.A2(n_1786),
.B1(n_1785),
.B2(n_1774),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1852),
.B(n_1855),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1846),
.B(n_1864),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1847),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1855),
.B(n_1805),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1855),
.B(n_1835),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1880),
.Y(n_1894)
);

OR2x6_ASAP7_75t_SL g1895 ( 
.A(n_1865),
.B(n_1778),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1880),
.Y(n_1896)
);

INVx2_ASAP7_75t_SL g1897 ( 
.A(n_1878),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1846),
.B(n_1791),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1866),
.B(n_1801),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1855),
.B(n_1727),
.Y(n_1900)
);

OAI33xp33_ASAP7_75t_L g1901 ( 
.A1(n_1864),
.A2(n_1781),
.A3(n_1768),
.B1(n_1757),
.B2(n_1765),
.B3(n_1759),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1839),
.Y(n_1902)
);

INVx1_ASAP7_75t_SL g1903 ( 
.A(n_1849),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1866),
.B(n_1792),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1839),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1854),
.B(n_1830),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1844),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1847),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1838),
.B(n_1738),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1838),
.B(n_1738),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1844),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1848),
.B(n_1829),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1879),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1879),
.Y(n_1914)
);

OAI21xp5_ASAP7_75t_L g1915 ( 
.A1(n_1865),
.A2(n_1804),
.B(n_1784),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1862),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1867),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1862),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1862),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1853),
.B(n_1816),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1867),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1853),
.Y(n_1922)
);

INVx3_ASAP7_75t_L g1923 ( 
.A(n_1874),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1845),
.B(n_1836),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1845),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1850),
.B(n_1763),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1872),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1838),
.B(n_1738),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1854),
.B(n_1825),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1838),
.B(n_1871),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1841),
.B(n_1764),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1863),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1872),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1857),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1881),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1899),
.B(n_1924),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1890),
.B(n_1860),
.Y(n_1937)
);

AOI211xp5_ASAP7_75t_L g1938 ( 
.A1(n_1915),
.A2(n_1861),
.B(n_1773),
.C(n_1787),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1881),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1930),
.B(n_1871),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1884),
.Y(n_1941)
);

INVx3_ASAP7_75t_SL g1942 ( 
.A(n_1885),
.Y(n_1942)
);

OAI21xp33_ASAP7_75t_L g1943 ( 
.A1(n_1888),
.A2(n_1904),
.B(n_1882),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1903),
.B(n_1920),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1884),
.Y(n_1945)
);

OAI32xp33_ASAP7_75t_L g1946 ( 
.A1(n_1895),
.A2(n_1874),
.A3(n_1876),
.B1(n_1857),
.B2(n_1873),
.Y(n_1946)
);

AOI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1892),
.A2(n_1904),
.B1(n_1901),
.B2(n_1882),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1886),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1930),
.B(n_1858),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1889),
.B(n_1842),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1889),
.B(n_1842),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1892),
.B(n_1851),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1893),
.B(n_1861),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1894),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1893),
.B(n_1897),
.Y(n_1955)
);

OR2x2_ASAP7_75t_L g1956 ( 
.A(n_1890),
.B(n_1876),
.Y(n_1956)
);

OAI21xp5_ASAP7_75t_SL g1957 ( 
.A1(n_1895),
.A2(n_1823),
.B(n_1779),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1897),
.B(n_1851),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1929),
.B(n_1868),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1929),
.B(n_1906),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1906),
.B(n_1850),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1894),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1896),
.B(n_1870),
.Y(n_1963)
);

NAND3xp33_ASAP7_75t_SL g1964 ( 
.A(n_1898),
.B(n_1896),
.C(n_1831),
.Y(n_1964)
);

INVx1_ASAP7_75t_SL g1965 ( 
.A(n_1883),
.Y(n_1965)
);

INVx1_ASAP7_75t_SL g1966 ( 
.A(n_1883),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1923),
.B(n_1870),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1900),
.B(n_1870),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1922),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1925),
.Y(n_1970)
);

INVx2_ASAP7_75t_SL g1971 ( 
.A(n_1883),
.Y(n_1971)
);

AOI21xp33_ASAP7_75t_SL g1972 ( 
.A1(n_1898),
.A2(n_1589),
.B(n_1815),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1902),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1934),
.B(n_1868),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1886),
.Y(n_1975)
);

NAND2x1_ASAP7_75t_L g1976 ( 
.A(n_1923),
.B(n_1752),
.Y(n_1976)
);

INVxp67_ASAP7_75t_SL g1977 ( 
.A(n_1923),
.Y(n_1977)
);

BUFx3_ASAP7_75t_L g1978 ( 
.A(n_1934),
.Y(n_1978)
);

AOI22x1_ASAP7_75t_L g1979 ( 
.A1(n_1913),
.A2(n_1874),
.B1(n_1877),
.B2(n_1545),
.Y(n_1979)
);

NOR2x1_ASAP7_75t_R g1980 ( 
.A(n_1931),
.B(n_1505),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_L g1981 ( 
.A(n_1912),
.B(n_1875),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1891),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1902),
.Y(n_1983)
);

INVx1_ASAP7_75t_SL g1984 ( 
.A(n_1909),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1900),
.B(n_1870),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1905),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1909),
.B(n_1840),
.Y(n_1987)
);

NOR2x1_ASAP7_75t_L g1988 ( 
.A(n_1891),
.B(n_1502),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1935),
.Y(n_1989)
);

INVx1_ASAP7_75t_SL g1990 ( 
.A(n_1942),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1939),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1942),
.B(n_1887),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1937),
.B(n_1913),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1941),
.Y(n_1994)
);

INVx1_ASAP7_75t_SL g1995 ( 
.A(n_1937),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_L g1996 ( 
.A(n_1980),
.B(n_1926),
.Y(n_1996)
);

OAI21xp5_ASAP7_75t_SL g1997 ( 
.A1(n_1957),
.A2(n_1789),
.B(n_1788),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1945),
.Y(n_1998)
);

NOR2xp67_ASAP7_75t_L g1999 ( 
.A(n_1971),
.B(n_1914),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1968),
.B(n_1910),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1968),
.B(n_1985),
.Y(n_2001)
);

INVx1_ASAP7_75t_SL g2002 ( 
.A(n_1988),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1973),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1983),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1936),
.B(n_1914),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_1960),
.B(n_1917),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1986),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1978),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1960),
.B(n_1959),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1985),
.B(n_1910),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1952),
.B(n_1928),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1978),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1954),
.Y(n_2013)
);

BUFx3_ASAP7_75t_L g2014 ( 
.A(n_1971),
.Y(n_2014)
);

INVx1_ASAP7_75t_SL g2015 ( 
.A(n_1965),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1947),
.B(n_1933),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1948),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1943),
.B(n_1938),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1962),
.Y(n_2019)
);

INVx1_ASAP7_75t_SL g2020 ( 
.A(n_1966),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1948),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1981),
.B(n_1944),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1975),
.Y(n_2023)
);

INVxp67_ASAP7_75t_L g2024 ( 
.A(n_1981),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1952),
.B(n_1950),
.Y(n_2025)
);

AOI22xp33_ASAP7_75t_L g2026 ( 
.A1(n_1964),
.A2(n_1928),
.B1(n_1834),
.B2(n_1794),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1969),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1975),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_2009),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1990),
.B(n_1961),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_2025),
.B(n_1955),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_2014),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_2025),
.B(n_1955),
.Y(n_2033)
);

OAI322xp33_ASAP7_75t_L g2034 ( 
.A1(n_2018),
.A2(n_1959),
.A3(n_1956),
.B1(n_1970),
.B2(n_1984),
.C1(n_1974),
.C2(n_1977),
.Y(n_2034)
);

HB1xp67_ASAP7_75t_L g2035 ( 
.A(n_2009),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2006),
.Y(n_2036)
);

INVxp33_ASAP7_75t_L g2037 ( 
.A(n_1992),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_2024),
.B(n_1950),
.Y(n_2038)
);

OAI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_1997),
.A2(n_1946),
.B(n_1972),
.Y(n_2039)
);

AOI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1997),
.A2(n_1953),
.B1(n_1963),
.B2(n_1949),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2006),
.Y(n_2041)
);

BUFx2_ASAP7_75t_L g2042 ( 
.A(n_2014),
.Y(n_2042)
);

OR2x2_ASAP7_75t_L g2043 ( 
.A(n_1995),
.B(n_1956),
.Y(n_2043)
);

OAI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_2002),
.A2(n_1979),
.B1(n_1953),
.B2(n_1976),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2008),
.B(n_1951),
.Y(n_2045)
);

AOI22xp5_ASAP7_75t_L g2046 ( 
.A1(n_2016),
.A2(n_1953),
.B1(n_1963),
.B2(n_1949),
.Y(n_2046)
);

OAI221xp5_ASAP7_75t_L g2047 ( 
.A1(n_2026),
.A2(n_1974),
.B1(n_1982),
.B2(n_1834),
.C(n_1820),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_2022),
.B(n_1963),
.Y(n_2048)
);

OAI211xp5_ASAP7_75t_L g2049 ( 
.A1(n_2015),
.A2(n_1982),
.B(n_1951),
.C(n_1958),
.Y(n_2049)
);

OR2x2_ASAP7_75t_L g2050 ( 
.A(n_2015),
.B(n_1940),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1989),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_SL g2052 ( 
.A(n_1999),
.B(n_1967),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1989),
.Y(n_2053)
);

BUFx3_ASAP7_75t_L g2054 ( 
.A(n_2008),
.Y(n_2054)
);

AOI221xp5_ASAP7_75t_SL g2055 ( 
.A1(n_2020),
.A2(n_1958),
.B1(n_1940),
.B2(n_1987),
.C(n_1877),
.Y(n_2055)
);

AOI211x1_ASAP7_75t_L g2056 ( 
.A1(n_2005),
.A2(n_1987),
.B(n_1933),
.C(n_1927),
.Y(n_2056)
);

OAI32xp33_ASAP7_75t_L g2057 ( 
.A1(n_2020),
.A2(n_1863),
.A3(n_1841),
.B1(n_1843),
.B2(n_1921),
.Y(n_2057)
);

NOR4xp25_ASAP7_75t_SL g2058 ( 
.A(n_2013),
.B(n_1812),
.C(n_1832),
.D(n_1907),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2035),
.Y(n_2059)
);

HB1xp67_ASAP7_75t_L g2060 ( 
.A(n_2042),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2043),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2031),
.B(n_2001),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_2050),
.B(n_1993),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2043),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_2039),
.B(n_1999),
.Y(n_2065)
);

OR2x2_ASAP7_75t_L g2066 ( 
.A(n_2030),
.B(n_1993),
.Y(n_2066)
);

INVx2_ASAP7_75t_SL g2067 ( 
.A(n_2032),
.Y(n_2067)
);

NOR2x1_ASAP7_75t_L g2068 ( 
.A(n_2054),
.B(n_2008),
.Y(n_2068)
);

INVxp67_ASAP7_75t_L g2069 ( 
.A(n_2052),
.Y(n_2069)
);

AOI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_2044),
.A2(n_1996),
.B1(n_2012),
.B2(n_2001),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2031),
.B(n_2011),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2029),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2054),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2032),
.B(n_2012),
.Y(n_2074)
);

INVxp67_ASAP7_75t_L g2075 ( 
.A(n_2052),
.Y(n_2075)
);

OR2x2_ASAP7_75t_L g2076 ( 
.A(n_2038),
.B(n_2045),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2033),
.B(n_2037),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_2036),
.B(n_2012),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2033),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2037),
.B(n_2011),
.Y(n_2080)
);

O2A1O1Ixp33_ASAP7_75t_L g2081 ( 
.A1(n_2065),
.A2(n_2034),
.B(n_2057),
.C(n_2053),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_2077),
.B(n_2040),
.Y(n_2082)
);

AOI21xp33_ASAP7_75t_L g2083 ( 
.A1(n_2065),
.A2(n_2041),
.B(n_2049),
.Y(n_2083)
);

AOI21xp33_ASAP7_75t_SL g2084 ( 
.A1(n_2069),
.A2(n_2048),
.B(n_2046),
.Y(n_2084)
);

NOR2x1_ASAP7_75t_L g2085 ( 
.A(n_2068),
.B(n_2014),
.Y(n_2085)
);

NAND3xp33_ASAP7_75t_L g2086 ( 
.A(n_2075),
.B(n_2058),
.C(n_2056),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2060),
.Y(n_2087)
);

OAI211xp5_ASAP7_75t_SL g2088 ( 
.A1(n_2070),
.A2(n_2048),
.B(n_2051),
.C(n_2047),
.Y(n_2088)
);

AOI322xp5_ASAP7_75t_L g2089 ( 
.A1(n_2077),
.A2(n_2055),
.A3(n_2013),
.B1(n_2019),
.B2(n_2027),
.C1(n_1998),
.C2(n_2007),
.Y(n_2089)
);

NAND4xp75_ASAP7_75t_L g2090 ( 
.A(n_2073),
.B(n_2019),
.C(n_2027),
.D(n_1998),
.Y(n_2090)
);

OAI21xp5_ASAP7_75t_L g2091 ( 
.A1(n_2080),
.A2(n_1994),
.B(n_1991),
.Y(n_2091)
);

AOI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_2060),
.A2(n_1994),
.B(n_1991),
.Y(n_2092)
);

OAI21xp5_ASAP7_75t_L g2093 ( 
.A1(n_2061),
.A2(n_2004),
.B(n_2003),
.Y(n_2093)
);

OA21x2_ASAP7_75t_L g2094 ( 
.A1(n_2074),
.A2(n_2021),
.B(n_2017),
.Y(n_2094)
);

OAI32xp33_ASAP7_75t_L g2095 ( 
.A1(n_2066),
.A2(n_2003),
.A3(n_2004),
.B1(n_2007),
.B2(n_2017),
.Y(n_2095)
);

OR2x2_ASAP7_75t_L g2096 ( 
.A(n_2087),
.B(n_2079),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2094),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2094),
.Y(n_2098)
);

NOR3x1_ASAP7_75t_L g2099 ( 
.A(n_2082),
.B(n_2067),
.C(n_2059),
.Y(n_2099)
);

OAI222xp33_ASAP7_75t_R g2100 ( 
.A1(n_2084),
.A2(n_2064),
.B1(n_2072),
.B2(n_2067),
.C1(n_2079),
.C2(n_2076),
.Y(n_2100)
);

NAND3xp33_ASAP7_75t_L g2101 ( 
.A(n_2083),
.B(n_2078),
.C(n_2063),
.Y(n_2101)
);

NAND4xp25_ASAP7_75t_SL g2102 ( 
.A(n_2081),
.B(n_2062),
.C(n_2071),
.D(n_2000),
.Y(n_2102)
);

NAND3xp33_ASAP7_75t_L g2103 ( 
.A(n_2086),
.B(n_2062),
.C(n_2071),
.Y(n_2103)
);

AOI211x1_ASAP7_75t_L g2104 ( 
.A1(n_2091),
.A2(n_2010),
.B(n_2000),
.C(n_1905),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_2085),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_2093),
.B(n_2010),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_2090),
.Y(n_2107)
);

NAND5xp2_ASAP7_75t_L g2108 ( 
.A(n_2089),
.B(n_1822),
.C(n_1833),
.D(n_1724),
.E(n_1917),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2106),
.B(n_2105),
.Y(n_2109)
);

NOR3xp33_ASAP7_75t_L g2110 ( 
.A(n_2103),
.B(n_2088),
.C(n_2092),
.Y(n_2110)
);

NOR3xp33_ASAP7_75t_L g2111 ( 
.A(n_2101),
.B(n_2095),
.C(n_2021),
.Y(n_2111)
);

NOR3x1_ASAP7_75t_L g2112 ( 
.A(n_2096),
.B(n_1927),
.C(n_1921),
.Y(n_2112)
);

NOR4xp25_ASAP7_75t_L g2113 ( 
.A(n_2107),
.B(n_2098),
.C(n_2097),
.D(n_2100),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2106),
.Y(n_2114)
);

NAND3xp33_ASAP7_75t_SL g2115 ( 
.A(n_2099),
.B(n_2021),
.C(n_2017),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2114),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2112),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2109),
.Y(n_2118)
);

NOR2xp33_ASAP7_75t_L g2119 ( 
.A(n_2110),
.B(n_2102),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_2111),
.B(n_2099),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2115),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2113),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2114),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2116),
.B(n_1967),
.Y(n_2124)
);

NOR2xp33_ASAP7_75t_SL g2125 ( 
.A(n_2120),
.B(n_2023),
.Y(n_2125)
);

NOR3xp33_ASAP7_75t_L g2126 ( 
.A(n_2119),
.B(n_2108),
.C(n_2028),
.Y(n_2126)
);

NOR3xp33_ASAP7_75t_L g2127 ( 
.A(n_2122),
.B(n_2028),
.C(n_2023),
.Y(n_2127)
);

OAI221xp5_ASAP7_75t_SL g2128 ( 
.A1(n_2121),
.A2(n_2104),
.B1(n_2028),
.B2(n_2023),
.C(n_1916),
.Y(n_2128)
);

OAI21xp5_ASAP7_75t_L g2129 ( 
.A1(n_2120),
.A2(n_1967),
.B(n_1916),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2123),
.B(n_1931),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_2124),
.B(n_2118),
.Y(n_2131)
);

NAND2x1p5_ASAP7_75t_L g2132 ( 
.A(n_2130),
.B(n_2117),
.Y(n_2132)
);

NOR2xp67_ASAP7_75t_L g2133 ( 
.A(n_2129),
.B(n_1908),
.Y(n_2133)
);

INVx2_ASAP7_75t_SL g2134 ( 
.A(n_2125),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2132),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2134),
.Y(n_2136)
);

XNOR2xp5_ASAP7_75t_L g2137 ( 
.A(n_2135),
.B(n_2131),
.Y(n_2137)
);

OAI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_2137),
.A2(n_2136),
.B1(n_2128),
.B2(n_2133),
.Y(n_2138)
);

AOI21xp33_ASAP7_75t_L g2139 ( 
.A1(n_2137),
.A2(n_2127),
.B(n_2126),
.Y(n_2139)
);

AOI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_2138),
.A2(n_1932),
.B1(n_1908),
.B2(n_1919),
.Y(n_2140)
);

OR2x2_ASAP7_75t_L g2141 ( 
.A(n_2139),
.B(n_1918),
.Y(n_2141)
);

OA21x2_ASAP7_75t_L g2142 ( 
.A1(n_2141),
.A2(n_1919),
.B(n_1918),
.Y(n_2142)
);

NAND3xp33_ASAP7_75t_L g2143 ( 
.A(n_2142),
.B(n_2140),
.C(n_1932),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2143),
.Y(n_2144)
);

OAI221xp5_ASAP7_75t_R g2145 ( 
.A1(n_2144),
.A2(n_1518),
.B1(n_1907),
.B2(n_1911),
.C(n_1863),
.Y(n_2145)
);

AOI211xp5_ASAP7_75t_L g2146 ( 
.A1(n_2145),
.A2(n_1587),
.B(n_1542),
.C(n_1539),
.Y(n_2146)
);


endmodule