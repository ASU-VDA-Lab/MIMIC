module fake_netlist_6_879_n_87 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_19, n_87);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;
input n_19;

output n_87;

wire n_52;
wire n_46;
wire n_21;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_77;
wire n_42;
wire n_24;
wire n_54;
wire n_32;
wire n_66;
wire n_85;
wire n_78;
wire n_84;
wire n_23;
wire n_20;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_80;
wire n_41;
wire n_86;
wire n_71;
wire n_74;
wire n_72;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx6p67_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

NAND2xp33_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_9),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_12),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_6),
.Y(n_39)
);

INVxp67_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_21),
.B1(n_27),
.B2(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_35),
.Y(n_49)
);

NOR2xp67_ASAP7_75t_R g50 ( 
.A(n_46),
.B(n_31),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_37),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_20),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_32),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_30),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_55),
.Y(n_60)
);

AND2x4_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_59),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_51),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_49),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_48),
.Y(n_66)
);

OAI211xp5_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_57),
.B(n_24),
.C(n_33),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_53),
.Y(n_68)
);

INVxp33_ASAP7_75t_SL g69 ( 
.A(n_63),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_SL g70 ( 
.A1(n_66),
.A2(n_28),
.B(n_26),
.Y(n_70)
);

AOI222xp33_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_24),
.B1(n_34),
.B2(n_31),
.C1(n_25),
.C2(n_33),
.Y(n_71)
);

A2O1A1O1Ixp25_ASAP7_75t_L g72 ( 
.A1(n_65),
.A2(n_34),
.B(n_31),
.C(n_25),
.D(n_50),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_23),
.B1(n_25),
.B2(n_31),
.Y(n_73)
);

OAI211xp5_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_68),
.B(n_73),
.C(n_69),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

OAI211xp5_ASAP7_75t_SL g76 ( 
.A1(n_72),
.A2(n_64),
.B(n_66),
.C(n_62),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_66),
.C(n_61),
.Y(n_77)
);

NOR5xp2_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_64),
.C(n_34),
.D(n_66),
.E(n_23),
.Y(n_78)
);

NAND4xp25_ASAP7_75t_SL g79 ( 
.A(n_71),
.B(n_61),
.C(n_23),
.D(n_18),
.Y(n_79)
);

NOR4xp75_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_61),
.C(n_17),
.D(n_14),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_81),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_77),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_81),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_79),
.B(n_61),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_85),
.A2(n_83),
.B1(n_86),
.B2(n_78),
.Y(n_87)
);


endmodule