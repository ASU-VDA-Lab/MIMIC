module fake_jpeg_2050_n_80 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_80);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_80;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_0),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_31),
.B1(n_28),
.B2(n_27),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_22),
.B1(n_26),
.B2(n_24),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_26),
.B1(n_24),
.B2(n_20),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_37),
.B1(n_38),
.B2(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_20),
.B1(n_24),
.B2(n_21),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_36),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_19),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2x1_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_34),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_35),
.B(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_51),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_43),
.B1(n_45),
.B2(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_28),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_52),
.B(n_28),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_49),
.B(n_46),
.Y(n_55)
);

AOI322xp5_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_58),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_59),
.C(n_28),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_0),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_45),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_47),
.B1(n_48),
.B2(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_31),
.B1(n_4),
.B2(n_6),
.Y(n_70)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

OAI21x1_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_66),
.B(n_18),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_50),
.B(n_2),
.C(n_3),
.Y(n_63)
);

AOI221xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_64),
.B1(n_60),
.B2(n_65),
.C(n_5),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_74)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_31),
.B(n_14),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_70),
.B(n_64),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_74),
.B1(n_71),
.B2(n_9),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_76),
.C(n_7),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_72),
.Y(n_76)
);

AOI221xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_13),
.Y(n_80)
);


endmodule