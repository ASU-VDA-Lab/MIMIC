module real_aes_11286_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_920, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_920;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_884;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_889;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_914;
wire n_203;
wire n_536;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g573 ( .A(n_0), .B(n_175), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_1), .A2(n_84), .B1(n_572), .B2(n_592), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g110 ( .A1(n_2), .A2(n_102), .B1(n_111), .B2(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_3), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_4), .B(n_147), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_5), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_6), .A2(n_38), .B1(n_138), .B2(n_547), .Y(n_627) );
NOR2xp67_ASAP7_75t_L g865 ( .A(n_7), .B(n_87), .Y(n_865) );
INVx1_ASAP7_75t_L g910 ( .A(n_7), .Y(n_910) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_8), .B(n_144), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_9), .B(n_126), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_10), .A2(n_63), .B1(n_138), .B2(n_219), .Y(n_548) );
NAND3xp33_ASAP7_75t_L g520 ( .A(n_11), .B(n_138), .C(n_172), .Y(n_520) );
NAND2x1p5_ASAP7_75t_L g187 ( .A(n_12), .B(n_126), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_13), .B(n_249), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_14), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_15), .B(n_516), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_16), .B(n_135), .Y(n_559) );
AND2x2_ASAP7_75t_L g218 ( .A(n_17), .B(n_219), .Y(n_218) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_18), .B(n_139), .C(n_144), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_19), .A2(n_27), .B1(n_144), .B2(n_547), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_20), .B(n_516), .Y(n_528) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_21), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_22), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_23), .B(n_174), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g892 ( .A(n_24), .Y(n_892) );
NAND2xp33_ASAP7_75t_L g182 ( .A(n_25), .B(n_183), .Y(n_182) );
NAND2xp33_ASAP7_75t_L g240 ( .A(n_26), .B(n_183), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g855 ( .A1(n_28), .A2(n_73), .B1(n_856), .B2(n_857), .Y(n_855) );
CKINVDCx5p33_ASAP7_75t_R g857 ( .A(n_28), .Y(n_857) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_29), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_30), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_31), .B(n_609), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_32), .A2(n_52), .B1(n_183), .B2(n_219), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_33), .B(n_139), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_34), .B(n_146), .Y(n_186) );
INVx1_ASAP7_75t_L g864 ( .A(n_35), .Y(n_864) );
NOR3xp33_ASAP7_75t_L g911 ( .A(n_35), .B(n_912), .C(n_915), .Y(n_911) );
OAI21x1_ASAP7_75t_L g128 ( .A1(n_36), .A2(n_66), .B(n_129), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_37), .A2(n_167), .B(n_224), .C(n_226), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_39), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_40), .B(n_138), .Y(n_137) );
NAND2xp33_ASAP7_75t_L g270 ( .A(n_41), .B(n_203), .Y(n_270) );
AND2x6_ASAP7_75t_L g152 ( .A(n_42), .B(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g550 ( .A(n_43), .B(n_155), .Y(n_550) );
NAND2x1p5_ASAP7_75t_L g521 ( .A(n_44), .B(n_155), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_45), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_46), .B(n_225), .Y(n_239) );
NAND2xp33_ASAP7_75t_L g253 ( .A(n_47), .B(n_203), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_48), .B(n_135), .Y(n_530) );
INVx1_ASAP7_75t_L g153 ( .A(n_49), .Y(n_153) );
AOI22x1_ASAP7_75t_SL g876 ( .A1(n_50), .A2(n_62), .B1(n_877), .B2(n_878), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_50), .Y(n_877) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_51), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_53), .B(n_203), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_54), .B(n_155), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_55), .B(n_144), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_56), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_57), .B(n_144), .Y(n_607) );
NAND2x1_ASAP7_75t_L g535 ( .A(n_58), .B(n_155), .Y(n_535) );
AND2x2_ASAP7_75t_L g228 ( .A(n_59), .B(n_174), .Y(n_228) );
AND2x2_ASAP7_75t_L g913 ( .A(n_60), .B(n_914), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_61), .B(n_172), .Y(n_571) );
INVx1_ASAP7_75t_L g878 ( .A(n_62), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_64), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_65), .B(n_601), .Y(n_600) );
HB1xp67_ASAP7_75t_L g883 ( .A(n_65), .Y(n_883) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_67), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_68), .Y(n_604) );
NAND2xp33_ASAP7_75t_L g163 ( .A(n_69), .B(n_135), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_70), .B(n_172), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_71), .A2(n_76), .B1(n_144), .B2(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_72), .B(n_181), .Y(n_269) );
INVx1_ASAP7_75t_L g856 ( .A(n_73), .Y(n_856) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_74), .Y(n_581) );
BUFx10_ASAP7_75t_L g862 ( .A(n_75), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_77), .B(n_134), .Y(n_237) );
INVx1_ASAP7_75t_SL g595 ( .A(n_78), .Y(n_595) );
NAND2xp33_ASAP7_75t_L g171 ( .A(n_79), .B(n_144), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_80), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g867 ( .A(n_81), .Y(n_867) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_82), .B(n_183), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_83), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_85), .Y(n_227) );
OAI22xp33_ASAP7_75t_SL g881 ( .A1(n_86), .A2(n_882), .B1(n_883), .B2(n_884), .Y(n_881) );
INVx1_ASAP7_75t_L g884 ( .A(n_86), .Y(n_884) );
AND2x2_ASAP7_75t_L g909 ( .A(n_87), .B(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g129 ( .A(n_88), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_89), .B(n_172), .Y(n_519) );
BUFx2_ASAP7_75t_L g115 ( .A(n_90), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_90), .B(n_863), .Y(n_870) );
OR2x2_ASAP7_75t_L g888 ( .A(n_90), .B(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g915 ( .A(n_90), .Y(n_915) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_91), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_92), .A2(n_105), .B1(n_907), .B2(n_916), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_93), .B(n_203), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_94), .B(n_155), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_95), .B(n_146), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_96), .Y(n_247) );
INVx1_ASAP7_75t_L g914 ( .A(n_97), .Y(n_914) );
INVx1_ASAP7_75t_L g217 ( .A(n_98), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_99), .Y(n_198) );
AND2x2_ASAP7_75t_L g209 ( .A(n_100), .B(n_126), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_101), .B(n_206), .Y(n_605) );
INVx1_ASAP7_75t_L g112 ( .A(n_102), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_103), .B(n_174), .Y(n_173) );
OR2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_895), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_871), .Y(n_106) );
AOI21xp33_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_854), .B(n_866), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_109), .A2(n_897), .B1(n_900), .B2(n_903), .Y(n_896) );
XNOR2x1_ASAP7_75t_L g109 ( .A(n_110), .B(n_113), .Y(n_109) );
OAI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_116), .B(n_502), .Y(n_113) );
NAND2xp33_ASAP7_75t_L g502 ( .A(n_114), .B(n_503), .Y(n_502) );
BUFx8_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI22x1_ASAP7_75t_L g874 ( .A1(n_116), .A2(n_875), .B1(n_876), .B2(n_879), .Y(n_874) );
INVx3_ASAP7_75t_L g879 ( .A(n_116), .Y(n_879) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_410), .Y(n_116) );
NOR4xp25_ASAP7_75t_L g117 ( .A(n_118), .B(n_307), .C(n_351), .D(n_370), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_292), .Y(n_118) );
AOI222xp33_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_188), .B1(n_229), .B2(n_258), .C1(n_273), .C2(n_282), .Y(n_119) );
AOI221xp5_ASAP7_75t_L g489 ( .A1(n_120), .A2(n_315), .B1(n_435), .B2(n_490), .C(n_492), .Y(n_489) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_157), .Y(n_120) );
BUFx2_ASAP7_75t_L g426 ( .A(n_121), .Y(n_426) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x4_ASAP7_75t_L g326 ( .A(n_122), .B(n_311), .Y(n_326) );
AND2x4_ASAP7_75t_L g404 ( .A(n_122), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g461 ( .A(n_122), .B(n_401), .Y(n_461) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g287 ( .A(n_124), .Y(n_287) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_124), .Y(n_407) );
OAI21x1_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_130), .B(n_154), .Y(n_124) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_125), .A2(n_178), .B(n_187), .Y(n_177) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_125), .A2(n_245), .B(n_254), .Y(n_244) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_125), .A2(n_130), .B(n_154), .Y(n_262) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_125), .A2(n_178), .B(n_187), .Y(n_291) );
BUFx4f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_126), .A2(n_161), .B(n_173), .Y(n_160) );
INVx4_ASAP7_75t_L g192 ( .A(n_126), .Y(n_192) );
INVx3_ASAP7_75t_L g233 ( .A(n_126), .Y(n_233) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_126), .A2(n_161), .B(n_173), .Y(n_285) );
OA21x2_ASAP7_75t_L g317 ( .A1(n_126), .A2(n_161), .B(n_173), .Y(n_317) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_126), .Y(n_613) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g156 ( .A(n_127), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_127), .B(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g175 ( .A(n_128), .Y(n_175) );
OAI21x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_140), .B(n_150), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B(n_137), .C(n_139), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g165 ( .A(n_135), .Y(n_165) );
INVx2_ASAP7_75t_L g249 ( .A(n_135), .Y(n_249) );
INVx1_ASAP7_75t_L g532 ( .A(n_135), .Y(n_532) );
INVx2_ASAP7_75t_L g572 ( .A(n_135), .Y(n_572) );
INVx2_ASAP7_75t_L g579 ( .A(n_135), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_135), .B(n_581), .Y(n_580) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_136), .Y(n_138) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
INVx2_ASAP7_75t_L g147 ( .A(n_136), .Y(n_147) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_136), .Y(n_206) );
INVx1_ASAP7_75t_L g221 ( .A(n_136), .Y(n_221) );
INVx5_ASAP7_75t_L g170 ( .A(n_138), .Y(n_170) );
BUFx12f_ASAP7_75t_L g149 ( .A(n_139), .Y(n_149) );
INVx5_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
INVx5_ASAP7_75t_L g172 ( .A(n_139), .Y(n_172) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_139), .A2(n_562), .B1(n_563), .B2(n_564), .Y(n_561) );
OAI321xp33_ASAP7_75t_L g569 ( .A1(n_139), .A2(n_144), .A3(n_570), .B1(n_571), .B2(n_572), .C(n_573), .Y(n_569) );
O2A1O1Ixp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B(n_145), .C(n_148), .Y(n_140) );
O2A1O1Ixp5_ASAP7_75t_L g184 ( .A1(n_142), .A2(n_148), .B(n_185), .C(n_186), .Y(n_184) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g181 ( .A(n_144), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_144), .B(n_196), .Y(n_195) );
INVx2_ASAP7_75t_SL g225 ( .A(n_144), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g603 ( .A1(n_144), .A2(n_172), .B(n_604), .C(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
INVx2_ASAP7_75t_L g203 ( .A(n_147), .Y(n_203) );
O2A1O1Ixp5_ASAP7_75t_L g246 ( .A1(n_148), .A2(n_247), .B(n_248), .C(n_250), .Y(n_246) );
OA22x2_ASAP7_75t_L g545 ( .A1(n_148), .A2(n_166), .B1(n_546), .B2(n_548), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_148), .A2(n_166), .B1(n_590), .B2(n_591), .Y(n_589) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_149), .Y(n_208) );
BUFx2_ASAP7_75t_L g222 ( .A(n_149), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_149), .A2(n_269), .B(n_270), .Y(n_268) );
AOI21x1_ASAP7_75t_L g529 ( .A1(n_149), .A2(n_530), .B(n_531), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_149), .A2(n_607), .B(n_608), .Y(n_606) );
OAI21x1_ASAP7_75t_L g161 ( .A1(n_150), .A2(n_162), .B(n_168), .Y(n_161) );
OAI21x1_ASAP7_75t_L g178 ( .A1(n_150), .A2(n_179), .B(n_184), .Y(n_178) );
OAI21x1_ASAP7_75t_L g234 ( .A1(n_150), .A2(n_235), .B(n_238), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_150), .A2(n_246), .B(n_251), .Y(n_245) );
AO31x2_ASAP7_75t_L g588 ( .A1(n_150), .A2(n_192), .A3(n_589), .B(n_593), .Y(n_588) );
AND2x2_ASAP7_75t_L g625 ( .A(n_150), .B(n_233), .Y(n_625) );
INVx8_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_151), .A2(n_194), .B(n_200), .Y(n_193) );
NOR2xp67_ASAP7_75t_L g212 ( .A(n_151), .B(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g544 ( .A(n_151), .Y(n_544) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_151), .A2(n_573), .B(n_583), .Y(n_582) );
INVx8_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx2_ASAP7_75t_L g271 ( .A(n_152), .Y(n_271) );
OAI21x1_ASAP7_75t_L g512 ( .A1(n_152), .A2(n_513), .B(n_518), .Y(n_512) );
OAI21x1_ASAP7_75t_L g557 ( .A1(n_152), .A2(n_558), .B(n_561), .Y(n_557) );
INVx1_ASAP7_75t_L g611 ( .A(n_152), .Y(n_611) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g366 ( .A(n_157), .B(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_158), .Y(n_429) );
NAND2x1p5_ASAP7_75t_L g158 ( .A(n_159), .B(n_176), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OR2x2_ASAP7_75t_L g377 ( .A(n_160), .B(n_289), .Y(n_377) );
AND2x2_ASAP7_75t_L g434 ( .A(n_160), .B(n_289), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_160), .B(n_342), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_166), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_166), .A2(n_180), .B(n_182), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_166), .A2(n_252), .B(n_253), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_166), .A2(n_208), .B1(n_627), .B2(n_628), .Y(n_626) );
CKINVDCx6p67_ASAP7_75t_R g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_SL g199 ( .A(n_167), .Y(n_199) );
AOI21x1_ASAP7_75t_L g526 ( .A1(n_167), .A2(n_527), .B(n_528), .Y(n_526) );
AOI21x1_ASAP7_75t_L g558 ( .A1(n_167), .A2(n_559), .B(n_560), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_167), .A2(n_575), .B(n_580), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_171), .B(n_172), .Y(n_168) );
NOR2xp67_ASAP7_75t_L g197 ( .A(n_170), .B(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g241 ( .A(n_172), .Y(n_241) );
AOI21x1_ASAP7_75t_L g265 ( .A1(n_172), .A2(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_L g543 ( .A(n_174), .Y(n_543) );
BUFx5_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_175), .Y(n_583) );
INVx1_ASAP7_75t_L g594 ( .A(n_175), .Y(n_594) );
INVx1_ASAP7_75t_L g259 ( .A(n_176), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_176), .B(n_287), .Y(n_330) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g318 ( .A(n_177), .B(n_295), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_183), .B(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g408 ( .A(n_190), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g453 ( .A(n_190), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_210), .Y(n_190) );
AND2x2_ASAP7_75t_L g299 ( .A(n_191), .B(n_257), .Y(n_299) );
OR2x2_ASAP7_75t_L g306 ( .A(n_191), .B(n_231), .Y(n_306) );
AND2x2_ASAP7_75t_L g459 ( .A(n_191), .B(n_244), .Y(n_459) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_209), .Y(n_191) );
INVx3_ASAP7_75t_L g213 ( .A(n_192), .Y(n_213) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_192), .A2(n_193), .B(n_209), .Y(n_280) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_197), .B(n_199), .Y(n_194) );
OAI21xp33_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_204), .B(n_208), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
NOR2xp33_ASAP7_75t_SL g204 ( .A(n_205), .B(n_207), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_205), .B(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g516 ( .A(n_206), .Y(n_516) );
INVx2_ASAP7_75t_L g547 ( .A(n_206), .Y(n_547) );
INVx2_ASAP7_75t_L g609 ( .A(n_206), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_208), .A2(n_236), .B(n_237), .Y(n_235) );
INVx1_ASAP7_75t_L g257 ( .A(n_210), .Y(n_257) );
AND2x2_ASAP7_75t_L g359 ( .A(n_210), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g438 ( .A(n_210), .Y(n_438) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g277 ( .A(n_211), .Y(n_277) );
AOI21x1_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_214), .B(n_228), .Y(n_211) );
OAI21x1_ASAP7_75t_L g524 ( .A1(n_213), .A2(n_525), .B(n_535), .Y(n_524) );
OAI21x1_ASAP7_75t_L g556 ( .A1(n_213), .A2(n_557), .B(n_565), .Y(n_556) );
OAI21x1_ASAP7_75t_L g618 ( .A1(n_213), .A2(n_557), .B(n_565), .Y(n_618) );
OAI21x1_ASAP7_75t_L g647 ( .A1(n_213), .A2(n_525), .B(n_535), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_223), .Y(n_214) );
OAI21x1_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_218), .B(n_222), .Y(n_215) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g592 ( .A(n_221), .Y(n_592) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_224), .A2(n_519), .B(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_229), .A2(n_372), .B1(n_374), .B2(n_378), .C(n_383), .Y(n_371) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_255), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_230), .B(n_389), .Y(n_388) );
NAND2xp67_ASAP7_75t_L g425 ( .A(n_230), .B(n_299), .Y(n_425) );
AND2x4_ASAP7_75t_L g480 ( .A(n_230), .B(n_359), .Y(n_480) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_243), .Y(n_230) );
INVx1_ASAP7_75t_L g281 ( .A(n_231), .Y(n_281) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_231), .Y(n_302) );
INVx1_ASAP7_75t_L g347 ( .A(n_231), .Y(n_347) );
INVx1_ASAP7_75t_L g396 ( .A(n_231), .Y(n_396) );
AND2x2_ASAP7_75t_L g437 ( .A(n_231), .B(n_438), .Y(n_437) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_234), .B(n_242), .Y(n_231) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_232), .A2(n_264), .B(n_272), .Y(n_263) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_232), .A2(n_264), .B(n_272), .Y(n_297) );
OAI21x1_ASAP7_75t_L g511 ( .A1(n_232), .A2(n_512), .B(n_521), .Y(n_511) );
OAI21x1_ASAP7_75t_L g693 ( .A1(n_232), .A2(n_512), .B(n_521), .Y(n_693) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_241), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_243), .B(n_280), .Y(n_337) );
OR2x2_ASAP7_75t_L g395 ( .A(n_243), .B(n_396), .Y(n_395) );
BUFx3_ASAP7_75t_L g484 ( .A(n_243), .Y(n_484) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g278 ( .A(n_244), .Y(n_278) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AOI22xp33_ASAP7_75t_SL g485 ( .A1(n_255), .A2(n_326), .B1(n_486), .B2(n_487), .Y(n_485) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g444 ( .A(n_256), .B(n_380), .Y(n_444) );
OR2x2_ASAP7_75t_L g488 ( .A(n_256), .B(n_306), .Y(n_488) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_258), .A2(n_293), .B1(n_298), .B2(n_303), .Y(n_292) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
OR2x2_ASAP7_75t_L g470 ( .A(n_259), .B(n_386), .Y(n_470) );
BUFx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g364 ( .A(n_261), .Y(n_364) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx1_ASAP7_75t_L g342 ( .A(n_262), .Y(n_342) );
OR2x2_ASAP7_75t_L g355 ( .A(n_262), .B(n_296), .Y(n_355) );
AND2x2_ASAP7_75t_L g452 ( .A(n_262), .B(n_289), .Y(n_452) );
BUFx2_ASAP7_75t_L g387 ( .A(n_263), .Y(n_387) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_268), .B(n_271), .Y(n_264) );
OAI21x1_ASAP7_75t_L g525 ( .A1(n_271), .A2(n_526), .B(n_529), .Y(n_525) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_279), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_276), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g305 ( .A(n_277), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_277), .B(n_278), .Y(n_333) );
INVxp67_ASAP7_75t_SL g390 ( .A(n_277), .Y(n_390) );
OR2x2_ASAP7_75t_L g301 ( .A(n_278), .B(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g381 ( .A(n_278), .Y(n_381) );
AND2x2_ASAP7_75t_L g431 ( .A(n_278), .B(n_347), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_278), .B(n_382), .Y(n_456) );
OR2x2_ASAP7_75t_L g332 ( .A(n_279), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g349 ( .A(n_280), .Y(n_349) );
INVx2_ASAP7_75t_SL g360 ( .A(n_280), .Y(n_360) );
INVx1_ASAP7_75t_L g416 ( .A(n_281), .Y(n_416) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
OR2x2_ASAP7_75t_L g468 ( .A(n_284), .B(n_343), .Y(n_468) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_SL g314 ( .A(n_285), .Y(n_314) );
INVx1_ASAP7_75t_SL g325 ( .A(n_285), .Y(n_325) );
BUFx2_ASAP7_75t_L g474 ( .A(n_285), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_286), .B(n_479), .Y(n_478) );
NAND2x1_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x4_ASAP7_75t_SL g310 ( .A(n_287), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g367 ( .A(n_287), .Y(n_367) );
BUFx2_ASAP7_75t_L g375 ( .A(n_287), .Y(n_375) );
INVx1_ASAP7_75t_L g423 ( .A(n_288), .Y(n_423) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_289), .B(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g313 ( .A(n_289), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g405 ( .A(n_290), .B(n_296), .Y(n_405) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g401 ( .A(n_291), .B(n_296), .Y(n_401) );
AND2x2_ASAP7_75t_L g350 ( .A(n_293), .B(n_317), .Y(n_350) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g406 ( .A(n_294), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g311 ( .A(n_295), .Y(n_311) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_298), .A2(n_316), .B1(n_413), .B2(n_418), .Y(n_412) );
AND2x4_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g368 ( .A(n_299), .Y(n_368) );
INVx1_ASAP7_75t_L g501 ( .A(n_299), .Y(n_501) );
INVx1_ASAP7_75t_L g447 ( .A(n_300), .Y(n_447) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OAI211xp5_ASAP7_75t_L g307 ( .A1(n_304), .A2(n_308), .B(n_319), .C(n_334), .Y(n_307) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g465 ( .A(n_305), .Y(n_465) );
INVx2_ASAP7_75t_L g382 ( .A(n_306), .Y(n_382) );
INVxp67_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
AO21x1_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_312), .B(n_315), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_310), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g373 ( .A(n_310), .Y(n_373) );
INVx1_ASAP7_75t_L g451 ( .A(n_311), .Y(n_451) );
BUFx2_ASAP7_75t_L g486 ( .A(n_311), .Y(n_486) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NOR2x1_ASAP7_75t_SL g363 ( .A(n_313), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_314), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g394 ( .A(n_314), .Y(n_394) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
OR2x6_ASAP7_75t_SL g354 ( .A(n_316), .B(n_355), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_316), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g322 ( .A(n_317), .Y(n_322) );
INVx2_ASAP7_75t_L g343 ( .A(n_318), .Y(n_343) );
OAI31xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_323), .A3(n_327), .B(n_331), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g483 ( .A(n_322), .B(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NOR2x1p5_ASAP7_75t_L g448 ( .A(n_325), .B(n_403), .Y(n_448) );
INVx2_ASAP7_75t_L g417 ( .A(n_326), .Y(n_417) );
INVxp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g491 ( .A(n_333), .Y(n_491) );
AOI22xp33_ASAP7_75t_SL g334 ( .A1(n_335), .A2(n_338), .B1(n_344), .B2(n_350), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g475 ( .A(n_336), .B(n_346), .Y(n_475) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_339), .A2(n_384), .B(n_388), .Y(n_383) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_343), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_340), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_SL g400 ( .A(n_341), .B(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVx1_ASAP7_75t_L g369 ( .A(n_346), .Y(n_369) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx2_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g436 ( .A(n_349), .B(n_437), .Y(n_436) );
O2A1O1Ixp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_356), .B(n_361), .C(n_369), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVxp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_354), .B(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g493 ( .A(n_355), .B(n_394), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_355), .A2(n_496), .B(n_498), .Y(n_495) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g415 ( .A(n_359), .B(n_416), .Y(n_415) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_360), .Y(n_399) );
AO21x1_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B(n_368), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_364), .A2(n_368), .B1(n_414), .B2(n_417), .Y(n_413) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI21xp5_ASAP7_75t_L g440 ( .A1(n_366), .A2(n_441), .B(n_444), .Y(n_440) );
AND2x2_ASAP7_75t_L g433 ( .A(n_367), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_391), .Y(n_370) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g477 ( .A(n_377), .Y(n_477) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
AND2x4_ASAP7_75t_L g435 ( .A(n_381), .B(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g500 ( .A(n_381), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g479 ( .A(n_387), .Y(n_479) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI32xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_397), .A3(n_400), .B1(n_402), .B2(n_408), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g420 ( .A(n_394), .Y(n_420) );
INVx1_ASAP7_75t_L g409 ( .A(n_395), .Y(n_409) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_398), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OAI21xp33_ASAP7_75t_L g498 ( .A1(n_400), .A2(n_453), .B(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g473 ( .A(n_401), .B(n_474), .Y(n_473) );
NAND2xp33_ASAP7_75t_SL g402 ( .A(n_403), .B(n_406), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NOR4xp75_ASAP7_75t_L g410 ( .A(n_411), .B(n_439), .C(n_481), .D(n_495), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_421), .C(n_432), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g454 ( .A(n_416), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_424), .B(n_426), .C(n_427), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI21xp5_ASAP7_75t_L g427 ( .A1(n_426), .A2(n_428), .B(n_430), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g466 ( .A(n_431), .Y(n_466) );
NAND2x1_ASAP7_75t_L g432 ( .A(n_433), .B(n_435), .Y(n_432) );
AND2x4_ASAP7_75t_L g458 ( .A(n_437), .B(n_459), .Y(n_458) );
NAND4xp75_ASAP7_75t_L g439 ( .A(n_440), .B(n_445), .C(n_462), .D(n_471), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI211x1_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_448), .B(n_449), .C(n_455), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_446), .A2(n_463), .B1(n_467), .B2(n_469), .Y(n_462) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_447), .B(n_493), .C(n_494), .Y(n_492) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_453), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B(n_460), .Y(n_455) );
NOR2xp67_ASAP7_75t_L g497 ( .A(n_457), .B(n_474), .Y(n_497) );
INVx2_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g494 ( .A(n_465), .Y(n_494) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_475), .B(n_476), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B(n_480), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_485), .B(n_489), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVxp67_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_754), .Y(n_503) );
NAND4xp25_ASAP7_75t_L g504 ( .A(n_505), .B(n_674), .C(n_701), .D(n_741), .Y(n_504) );
NOR3xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_631), .C(n_648), .Y(n_505) );
OAI21xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_551), .B(n_584), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_536), .Y(n_507) );
AND2x2_ASAP7_75t_L g742 ( .A(n_508), .B(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_522), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_509), .B(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g586 ( .A(n_510), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_510), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g651 ( .A(n_510), .B(n_597), .Y(n_651) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g663 ( .A(n_511), .B(n_612), .Y(n_663) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_517), .Y(n_513) );
INVxp67_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx2_ASAP7_75t_L g660 ( .A(n_522), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_522), .B(n_616), .Y(n_808) );
INVx1_ASAP7_75t_L g814 ( .A(n_522), .Y(n_814) );
OR2x2_ASAP7_75t_L g852 ( .A(n_522), .B(n_616), .Y(n_852) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_523), .Y(n_671) );
OR2x2_ASAP7_75t_L g803 ( .A(n_523), .B(n_623), .Y(n_803) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g620 ( .A(n_524), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g563 ( .A(n_532), .Y(n_563) );
INVx4_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2x1p5_ASAP7_75t_L g853 ( .A(n_537), .B(n_805), .Y(n_853) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g732 ( .A(n_540), .B(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g743 ( .A(n_540), .B(n_719), .Y(n_743) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g677 ( .A(n_541), .Y(n_677) );
INVxp67_ASAP7_75t_SL g695 ( .A(n_541), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_541), .B(n_588), .Y(n_707) );
INVx1_ASAP7_75t_L g748 ( .A(n_541), .Y(n_748) );
HB1xp67_ASAP7_75t_L g838 ( .A(n_541), .Y(n_838) );
OAI21x1_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_545), .B(n_549), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
OA21x2_ASAP7_75t_L g612 ( .A1(n_545), .A2(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVxp67_ASAP7_75t_L g614 ( .A(n_550), .Y(n_614) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g761 ( .A(n_553), .B(n_671), .Y(n_761) );
INVx4_ASAP7_75t_L g815 ( .A(n_553), .Y(n_815) );
AND2x4_ASAP7_75t_L g553 ( .A(n_554), .B(n_566), .Y(n_553) );
AND2x2_ASAP7_75t_L g725 ( .A(n_554), .B(n_654), .Y(n_725) );
AND2x2_ASAP7_75t_L g735 ( .A(n_554), .B(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g653 ( .A(n_555), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_555), .B(n_640), .Y(n_764) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g680 ( .A(n_556), .Y(n_680) );
AND2x2_ASAP7_75t_L g752 ( .A(n_556), .B(n_641), .Y(n_752) );
BUFx2_ASAP7_75t_L g744 ( .A(n_566), .Y(n_744) );
AND2x2_ASAP7_75t_L g760 ( .A(n_566), .B(n_659), .Y(n_760) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g673 ( .A(n_567), .B(n_640), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_567), .B(n_620), .Y(n_730) );
AND2x2_ASAP7_75t_L g825 ( .A(n_567), .B(n_647), .Y(n_825) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g641 ( .A(n_568), .Y(n_641) );
AND2x2_ASAP7_75t_L g654 ( .A(n_568), .B(n_623), .Y(n_654) );
OAI21x1_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_574), .B(n_582), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_615), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_585), .B(n_824), .Y(n_830) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_596), .Y(n_585) );
INVx2_ASAP7_75t_L g697 ( .A(n_586), .Y(n_697) );
INVx1_ASAP7_75t_L g665 ( .A(n_587), .Y(n_665) );
AND2x4_ASAP7_75t_L g719 ( .A(n_587), .B(n_635), .Y(n_719) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g656 ( .A(n_588), .Y(n_656) );
INVx1_ASAP7_75t_L g668 ( .A(n_588), .Y(n_668) );
AND2x2_ASAP7_75t_L g714 ( .A(n_588), .B(n_612), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx1_ASAP7_75t_L g601 ( .A(n_594), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_594), .B(n_630), .Y(n_629) );
AND2x4_ASAP7_75t_L g721 ( .A(n_596), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_612), .Y(n_596) );
AND2x2_ASAP7_75t_L g667 ( .A(n_597), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g710 ( .A(n_597), .Y(n_710) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g733 ( .A(n_598), .B(n_693), .Y(n_733) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g635 ( .A(n_599), .Y(n_635) );
AND2x2_ASAP7_75t_L g692 ( .A(n_599), .B(n_693), .Y(n_692) );
NAND2x1p5_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
OAI21x1_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_606), .B(n_610), .Y(n_602) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_619), .Y(n_615) );
OR2x2_ASAP7_75t_L g818 ( .A(n_616), .B(n_641), .Y(n_818) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_SL g643 ( .A(n_617), .Y(n_643) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g659 ( .A(n_618), .Y(n_659) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVxp67_ASAP7_75t_SL g771 ( .A(n_620), .Y(n_771) );
BUFx2_ASAP7_75t_L g796 ( .A(n_620), .Y(n_796) );
AND2x2_ASAP7_75t_L g782 ( .A(n_621), .B(n_645), .Y(n_782) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_622), .B(n_659), .Y(n_658) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_622), .Y(n_751) );
AND2x2_ASAP7_75t_L g780 ( .A(n_622), .B(n_646), .Y(n_780) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_623), .Y(n_729) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g640 ( .A(n_624), .Y(n_640) );
AOI21x1_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B(n_629), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_636), .Y(n_631) );
INVxp67_ASAP7_75t_SL g689 ( .A(n_632), .Y(n_689) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_633), .B(n_714), .Y(n_753) );
AND2x2_ASAP7_75t_L g809 ( .A(n_633), .B(n_714), .Y(n_809) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g664 ( .A(n_635), .B(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_642), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g786 ( .A(n_639), .B(n_787), .Y(n_786) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_640), .Y(n_737) );
AND2x2_ASAP7_75t_L g679 ( .A(n_641), .B(n_680), .Y(n_679) );
INVxp67_ASAP7_75t_SL g700 ( .A(n_641), .Y(n_700) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
AND2x4_ASAP7_75t_L g781 ( .A(n_643), .B(n_782), .Y(n_781) );
AND2x2_ASAP7_75t_L g678 ( .A(n_644), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g688 ( .A(n_644), .Y(n_688) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g650 ( .A(n_645), .B(n_651), .Y(n_650) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_645), .Y(n_759) );
AND2x2_ASAP7_75t_L g773 ( .A(n_645), .B(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI322xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_652), .A3(n_655), .B1(n_657), .B2(n_661), .C1(n_666), .C2(n_669), .Y(n_648) );
OAI322xp33_ASAP7_75t_L g810 ( .A1(n_649), .A2(n_811), .A3(n_812), .B1(n_813), .B2(n_816), .C1(n_819), .C2(n_920), .Y(n_810) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g790 ( .A(n_651), .B(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_653), .Y(n_702) );
AND2x2_ASAP7_75t_L g795 ( .A(n_654), .B(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g844 ( .A(n_654), .Y(n_844) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2x1_ASAP7_75t_L g767 ( .A(n_656), .B(n_768), .Y(n_767) );
OR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_658), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g788 ( .A(n_659), .Y(n_788) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
AND2x2_ASAP7_75t_L g739 ( .A(n_663), .B(n_740), .Y(n_739) );
INVxp67_ASAP7_75t_L g723 ( .A(n_665), .Y(n_723) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g675 ( .A(n_667), .B(n_676), .Y(n_675) );
NOR2xp67_ASAP7_75t_L g740 ( .A(n_668), .B(n_710), .Y(n_740) );
INVx1_ASAP7_75t_L g849 ( .A(n_668), .Y(n_849) );
OR2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_670), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_672), .A2(n_746), .B1(n_749), .B2(n_753), .Y(n_745) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AND2x4_ASAP7_75t_L g687 ( .A(n_673), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g833 ( .A(n_673), .B(n_788), .Y(n_833) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_678), .B1(n_681), .B2(n_689), .C(n_690), .Y(n_674) );
INVxp67_ASAP7_75t_L g769 ( .A(n_675), .Y(n_769) );
INVx1_ASAP7_75t_L g682 ( .A(n_676), .Y(n_682) );
OR2x2_ASAP7_75t_L g696 ( .A(n_676), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g766 ( .A(n_676), .B(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI21xp33_ASAP7_75t_SL g806 ( .A1(n_678), .A2(n_807), .B(n_809), .Y(n_806) );
INVx2_ASAP7_75t_L g685 ( .A(n_679), .Y(n_685) );
AND2x2_ASAP7_75t_L g789 ( .A(n_679), .B(n_737), .Y(n_789) );
OAI21xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B(n_686), .Y(n_681) );
INVx1_ASAP7_75t_L g811 ( .A(n_684), .Y(n_811) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI21xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_696), .B(n_698), .Y(n_690) );
INVx2_ASAP7_75t_L g829 ( .A(n_691), .Y(n_829) );
NAND2x1p5_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
AND2x2_ASAP7_75t_L g820 ( .A(n_692), .B(n_748), .Y(n_820) );
BUFx3_ASAP7_75t_L g713 ( .A(n_693), .Y(n_713) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NOR2x1p5_ASAP7_75t_L g798 ( .A(n_697), .B(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI211xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B(n_715), .C(n_726), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_711), .Y(n_703) );
OAI21xp33_ASAP7_75t_L g831 ( .A1(n_704), .A2(n_832), .B(n_834), .Y(n_831) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVxp67_ASAP7_75t_L g791 ( .A(n_707), .Y(n_791) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g783 ( .A(n_709), .B(n_714), .Y(n_783) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g800 ( .A(n_710), .B(n_748), .Y(n_800) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx2_ASAP7_75t_L g717 ( .A(n_713), .Y(n_717) );
NOR2xp67_ASAP7_75t_L g722 ( .A(n_713), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g812 ( .A(n_714), .Y(n_812) );
AOI21xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_720), .B(n_724), .Y(n_715) );
OR2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
AND2x4_ASAP7_75t_L g805 ( .A(n_717), .B(n_719), .Y(n_805) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g747 ( .A(n_719), .Y(n_747) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
OAI22xp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_731), .B1(n_734), .B2(n_738), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g768 ( .A(n_733), .Y(n_768) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AOI21xp5_ASAP7_75t_R g741 ( .A1(n_742), .A2(n_744), .B(n_745), .Y(n_741) );
OAI221xp5_ASAP7_75t_L g822 ( .A1(n_746), .A2(n_823), .B1(n_826), .B2(n_827), .C(n_830), .Y(n_822) );
OR2x6_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NOR2xp33_ASAP7_75t_SL g816 ( .A(n_750), .B(n_817), .Y(n_816) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
AND2x2_ASAP7_75t_L g824 ( .A(n_751), .B(n_825), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_752), .B(n_771), .Y(n_770) );
AND2x2_ASAP7_75t_L g777 ( .A(n_752), .B(n_778), .Y(n_777) );
NAND3xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_792), .C(n_821), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_775), .Y(n_755) );
OAI221xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_765), .B1(n_769), .B2(n_770), .C(n_772), .Y(n_756) );
NOR3xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_761), .C(n_762), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g823 ( .A1(n_760), .A2(n_778), .B(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_SL g774 ( .A(n_764), .Y(n_774) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_767), .B(n_773), .Y(n_772) );
NOR2xp67_ASAP7_75t_L g817 ( .A(n_771), .B(n_818), .Y(n_817) );
OAI21xp5_ASAP7_75t_L g834 ( .A1(n_773), .A2(n_835), .B(n_839), .Y(n_834) );
NAND2xp5_ASAP7_75t_SL g775 ( .A(n_776), .B(n_784), .Y(n_775) );
OAI21xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_781), .B(n_783), .Y(n_776) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_781), .B(n_851), .Y(n_850) );
OAI21xp33_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_789), .B(n_790), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_787), .B(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
BUFx2_ASAP7_75t_L g839 ( .A(n_791), .Y(n_839) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_810), .Y(n_792) );
OAI221xp5_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_797), .B1(n_801), .B2(n_804), .C(n_806), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NOR2xp33_ASAP7_75t_SL g841 ( .A(n_802), .B(n_842), .Y(n_841) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVxp67_ASAP7_75t_SL g807 ( .A(n_808), .Y(n_807) );
OR2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
INVx2_ASAP7_75t_L g845 ( .A(n_815), .Y(n_845) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
NOR3xp33_ASAP7_75t_SL g821 ( .A(n_822), .B(n_831), .C(n_840), .Y(n_821) );
INVx1_ASAP7_75t_L g826 ( .A(n_825), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
BUFx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
AND2x4_ASAP7_75t_L g847 ( .A(n_829), .B(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
OAI22xp33_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_846), .B1(n_850), .B2(n_853), .Y(n_840) );
NOR2x1_ASAP7_75t_L g842 ( .A(n_843), .B(n_845), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_SL g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx2_ASAP7_75t_SL g851 ( .A(n_852), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_858), .Y(n_854) );
CKINVDCx5p33_ASAP7_75t_R g899 ( .A(n_855), .Y(n_899) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
BUFx12f_ASAP7_75t_SL g898 ( .A(n_860), .Y(n_898) );
OR2x6_ASAP7_75t_L g860 ( .A(n_861), .B(n_863), .Y(n_860) );
OR2x2_ASAP7_75t_L g869 ( .A(n_861), .B(n_870), .Y(n_869) );
HB1xp67_ASAP7_75t_SL g894 ( .A(n_861), .Y(n_894) );
INVx2_ASAP7_75t_SL g861 ( .A(n_862), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g902 ( .A(n_862), .Y(n_902) );
INVx2_ASAP7_75t_L g889 ( .A(n_863), .Y(n_889) );
AND2x4_ASAP7_75t_L g863 ( .A(n_864), .B(n_865), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g866 ( .A(n_867), .B(n_868), .Y(n_866) );
BUFx12f_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
NAND2xp5_ASAP7_75t_SL g871 ( .A(n_872), .B(n_894), .Y(n_871) );
OAI21xp5_ASAP7_75t_L g872 ( .A1(n_873), .A2(n_880), .B(n_890), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
NOR2xp33_ASAP7_75t_SL g903 ( .A(n_874), .B(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_885), .Y(n_880) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_881), .B(n_901), .Y(n_900) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_883), .Y(n_882) );
INVx4_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx4_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
BUFx6f_ASAP7_75t_L g893 ( .A(n_887), .Y(n_893) );
INVx5_ASAP7_75t_L g906 ( .A(n_887), .Y(n_906) );
BUFx6f_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
NAND2xp5_ASAP7_75t_SL g895 ( .A(n_890), .B(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_892), .B(n_893), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .Y(n_897) );
CKINVDCx5p33_ASAP7_75t_R g901 ( .A(n_902), .Y(n_901) );
INVx4_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx6_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
BUFx6f_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx2_ASAP7_75t_L g918 ( .A(n_908), .Y(n_918) );
AND2x2_ASAP7_75t_SL g908 ( .A(n_909), .B(n_911), .Y(n_908) );
INVx4_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
CKINVDCx5p33_ASAP7_75t_R g916 ( .A(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
endmodule