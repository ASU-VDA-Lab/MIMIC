module real_jpeg_24874_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_0),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_0),
.B(n_49),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_0),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_0),
.B(n_47),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_1),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_1),
.B(n_47),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_1),
.B(n_67),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_1),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_1),
.B(n_33),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_1),
.B(n_52),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_1),
.B(n_49),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_2),
.B(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_2),
.B(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_2),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_2),
.B(n_33),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_2),
.B(n_52),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_7),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_7),
.B(n_27),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_7),
.B(n_74),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_7),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_7),
.B(n_33),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_7),
.B(n_52),
.Y(n_276)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_10),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_10),
.B(n_27),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_10),
.B(n_33),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_10),
.B(n_17),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_10),
.B(n_52),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_10),
.B(n_49),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_10),
.B(n_47),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_10),
.B(n_67),
.Y(n_268)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_12),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_12),
.B(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_12),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_12),
.B(n_33),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_12),
.B(n_52),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_12),
.B(n_49),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_12),
.B(n_47),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_12),
.B(n_67),
.Y(n_291)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_13),
.B(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_14),
.B(n_47),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_14),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_14),
.B(n_52),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_14),
.B(n_67),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_14),
.B(n_232),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_15),
.B(n_49),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_15),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_15),
.B(n_33),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_15),
.B(n_47),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_15),
.B(n_67),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_15),
.B(n_27),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_16),
.B(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_16),
.B(n_52),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_16),
.B(n_33),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_16),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_16),
.B(n_49),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_16),
.B(n_47),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_16),
.B(n_67),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_16),
.B(n_27),
.Y(n_257)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_17),
.Y(n_162)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_17),
.Y(n_193)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_17),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_148),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_119),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_80),
.C(n_92),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_21),
.B(n_80),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_54),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_22),
.B(n_55),
.C(n_71),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_45),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_23),
.B(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_24),
.B(n_30),
.C(n_37),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_26),
.B(n_61),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_30),
.A2(n_38),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_SL g133 ( 
.A(n_30),
.B(n_82),
.C(n_85),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_31),
.B(n_62),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_32),
.B(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_35),
.A2(n_37),
.B1(n_40),
.B2(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_36),
.B(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_36),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_40),
.C(n_41),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_39),
.B(n_45),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_40),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_41),
.A2(n_42),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_44),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_45),
.Y(n_329)
);

FAx1_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.CI(n_51),
.CON(n_45),
.SN(n_45)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_48),
.C(n_51),
.Y(n_87)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_52),
.Y(n_179)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_71),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_66),
.C(n_70),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_56),
.A2(n_57),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_60),
.C(n_63),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_63),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_73),
.B1(n_77),
.B2(n_78),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_66),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_66),
.A2(n_70),
.B1(n_78),
.B2(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_66),
.B(n_77),
.C(n_79),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_70),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_79),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_73),
.Y(n_77)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_87),
.C(n_88),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_84),
.A2(n_85),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_88),
.Y(n_332)
);

FAx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_90),
.CI(n_91),
.CON(n_88),
.SN(n_88)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_90),
.C(n_91),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_92),
.B(n_328),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_106),
.C(n_110),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_93),
.B(n_324),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.C(n_102),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_94),
.B(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_96),
.B(n_102),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.C(n_100),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_99),
.B(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_106),
.B(n_110),
.Y(n_324)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_117),
.C(n_118),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_111),
.B(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.C(n_115),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_112),
.B(n_115),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_114),
.B(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_117),
.B(n_118),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_134),
.B2(n_135),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_130),
.B2(n_131),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_128),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_146),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_326),
.C(n_327),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_316),
.C(n_317),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_302),
.C(n_303),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_279),
.C(n_280),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_247),
.C(n_248),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_226),
.C(n_227),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_206),
.C(n_207),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_184),
.C(n_185),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_170),
.C(n_175),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_166),
.B2(n_167),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_168),
.C(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_160),
.Y(n_165)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_162),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.C(n_180),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_178),
.B(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_197),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_190),
.C(n_197),
.Y(n_206)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_190)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_191),
.Y(n_196)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_194),
.B(n_196),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_205),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_198),
.Y(n_205)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_201),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_204),
.C(n_205),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_215),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_210),
.C(n_215),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_213),
.C(n_214),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_218),
.C(n_219),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_225),
.Y(n_219)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_220),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_225),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_241),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_242),
.C(n_246),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_237),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_236),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_236),
.C(n_237),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_231),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_235),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_237),
.Y(n_333)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.CI(n_240),
.CON(n_237),
.SN(n_237)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_239),
.C(n_240),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_242),
.Y(n_264)
);

FAx1_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_244),
.CI(n_245),
.CON(n_242),
.SN(n_242)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_263),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_252),
.C(n_263),
.Y(n_279)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_259),
.C(n_262),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_254),
.Y(n_331)
);

FAx1_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_256),
.CI(n_257),
.CON(n_254),
.SN(n_254)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_256),
.C(n_257),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_270),
.C(n_277),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_270),
.B1(n_277),
.B2(n_278),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_266),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B(n_269),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_268),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_298),
.C(n_299),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_270),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_274),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_275),
.C(n_276),
.Y(n_293)
);

INVx11_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_294),
.B2(n_301),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_295),
.C(n_296),
.Y(n_302)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_285),
.C(n_287),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_293),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_292),
.C(n_293),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_291),
.Y(n_292)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_314),
.B2(n_315),
.Y(n_303)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_304),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_308),
.C(n_314),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_311),
.C(n_312),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_320),
.C(n_325),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_323),
.B2(n_325),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_323),
.Y(n_325)
);


endmodule