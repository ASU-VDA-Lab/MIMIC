module fake_aes_2233_n_23 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_23);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_23;
wire n_20;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
BUFx6f_ASAP7_75t_SL g10 ( .A(n_5), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
BUFx3_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
AND2x2_ASAP7_75t_SL g15 ( .A(n_3), .B(n_8), .Y(n_15) );
OAI21xp5_ASAP7_75t_L g16 ( .A1(n_12), .A2(n_4), .B(n_6), .Y(n_16) );
AO21x2_ASAP7_75t_L g17 ( .A1(n_11), .A2(n_1), .B(n_2), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_17), .B(n_14), .Y(n_18) );
INVxp67_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
AOI21xp5_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_16), .B(n_17), .Y(n_20) );
NOR3xp33_ASAP7_75t_L g21 ( .A(n_20), .B(n_15), .C(n_10), .Y(n_21) );
AOI31xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_10), .A3(n_2), .B(n_1), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_13), .Y(n_23) );
endmodule