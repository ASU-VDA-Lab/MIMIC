module fake_jpeg_14329_n_166 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_166);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_11),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_74),
.Y(n_81)
);

BUFx24_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_79),
.C(n_49),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_76),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_78),
.Y(n_88)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_56),
.B1(n_68),
.B2(n_61),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_67),
.C(n_56),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_83),
.C(n_89),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_59),
.B1(n_68),
.B2(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_69),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_63),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_64),
.B1(n_66),
.B2(n_55),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_92),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_76),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_3),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_65),
.B1(n_53),
.B2(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_54),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_99),
.Y(n_121)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_89),
.A2(n_60),
.B(n_58),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_12),
.B(n_13),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_106),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_9),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_57),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_105),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_51),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_22),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_0),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_2),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_10),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_117),
.A2(n_120),
.B(n_19),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_28),
.C(n_45),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_109),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_98),
.A2(n_4),
.B(n_5),
.Y(n_120)
);

AO21x1_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_125),
.B(n_133),
.Y(n_147)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_128),
.B(n_129),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_11),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_131),
.B(n_12),
.Y(n_139)
);

AO22x1_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_31),
.B1(n_42),
.B2(n_14),
.Y(n_134)
);

AO22x1_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_113),
.B1(n_100),
.B2(n_13),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_132),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_139),
.B(n_142),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_144),
.B(n_133),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_124),
.A2(n_106),
.B1(n_16),
.B2(n_18),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_SL g149 ( 
.A1(n_141),
.A2(n_148),
.B(n_125),
.C(n_134),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_15),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_146),
.B(n_119),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_23),
.B1(n_25),
.B2(n_29),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_118),
.B(n_30),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_145),
.B(n_146),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_126),
.B(n_32),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_150),
.C(n_151),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_137),
.Y(n_150)
);

AOI221xp5_ASAP7_75t_L g156 ( 
.A1(n_153),
.A2(n_155),
.B1(n_135),
.B2(n_116),
.C(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_159),
.Y(n_160)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_148),
.B1(n_147),
.B2(n_140),
.Y(n_161)
);

AOI31xp67_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_157),
.A3(n_139),
.B(n_152),
.Y(n_162)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_162),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_160),
.B1(n_161),
.B2(n_152),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_145),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_136),
.Y(n_166)
);


endmodule