module fake_ibex_1715_n_2347 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_421, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_426, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_434, n_296, n_120, n_168, n_155, n_315, n_441, n_13, n_122, n_116, n_370, n_431, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_437, n_355, n_407, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_444, n_199, n_410, n_308, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_408, n_119, n_361, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_443, n_344, n_393, n_436, n_428, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_425, n_2347);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_434;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_437;
input n_355;
input n_407;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_444;
input n_199;
input n_410;
input n_308;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2347;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_452;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2151;
wire n_1391;
wire n_884;
wire n_667;
wire n_850;
wire n_1971;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_557;
wire n_641;
wire n_1937;
wire n_2311;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_2249;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_2275;
wire n_1853;
wire n_2189;
wire n_745;
wire n_2112;
wire n_447;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_2203;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_455;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_1121;
wire n_693;
wire n_2256;
wire n_606;
wire n_737;
wire n_1571;
wire n_1980;
wire n_462;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_816;
wire n_1058;
wire n_1835;
wire n_2224;
wire n_1862;
wire n_1543;
wire n_823;
wire n_2233;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_2312;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_1210;
wire n_2319;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2006;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1566;
wire n_1464;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_1982;
wire n_2252;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_1120;
wire n_2300;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_2160;
wire n_2234;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_650;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_817;
wire n_2193;
wire n_2095;
wire n_555;
wire n_951;
wire n_2053;
wire n_468;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_502;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_532;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_2170;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2243;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_2106;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_2298;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_2110;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_2344;
wire n_2317;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2210;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_636;
wire n_1259;
wire n_490;
wire n_2108;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_1725;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1415;
wire n_1238;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_1270;
wire n_834;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_484;
wire n_1642;
wire n_1455;
wire n_1871;
wire n_480;
wire n_2182;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_1403;
wire n_2181;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_2272;
wire n_535;
wire n_1956;
wire n_681;
wire n_1718;
wire n_2225;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_786;
wire n_505;
wire n_2043;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2121;
wire n_1893;
wire n_1570;
wire n_2231;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1961;
wire n_1050;
wire n_2218;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1542;
wire n_1097;
wire n_1909;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_478;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_753;
wire n_2126;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_2131;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_755;
wire n_2091;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_2337;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2323;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2227;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_924;
wire n_2331;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2092;
wire n_566;
wire n_581;
wire n_1365;
wire n_1472;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_548;
wire n_1158;
wire n_1974;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_2327;
wire n_913;
wire n_509;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_1902;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

INVx1_ASAP7_75t_L g446 ( 
.A(n_189),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_66),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_276),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_218),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_29),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_435),
.B(n_277),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_339),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_179),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_377),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_27),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_403),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_165),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_140),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_30),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_333),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_342),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_54),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_93),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_386),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_260),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_373),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_381),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_396),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_369),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_311),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_401),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_427),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_388),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_385),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_15),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_176),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_393),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_10),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_376),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_267),
.Y(n_480)
);

INVxp33_ASAP7_75t_SL g481 ( 
.A(n_352),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_445),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_102),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_356),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_329),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_202),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_394),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_425),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_336),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_249),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_238),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_40),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_438),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_325),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_440),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_256),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_290),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_221),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_379),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_371),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_93),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_289),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_288),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_27),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_8),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_81),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_78),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_123),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_357),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_358),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_367),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_177),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_423),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_412),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_268),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_127),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_405),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_210),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_133),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_112),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_317),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_399),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_41),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_289),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_64),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_337),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_408),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_400),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_268),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_407),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_91),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_249),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_70),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_319),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_17),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_312),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_265),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_285),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_272),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_124),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_123),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_209),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_162),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_372),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_416),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_343),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_263),
.Y(n_547)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_206),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_384),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_227),
.Y(n_550)
);

CKINVDCx16_ASAP7_75t_R g551 ( 
.A(n_344),
.Y(n_551)
);

CKINVDCx16_ASAP7_75t_R g552 ( 
.A(n_153),
.Y(n_552)
);

CKINVDCx14_ASAP7_75t_R g553 ( 
.A(n_100),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_398),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_253),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_153),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_225),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_239),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_375),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_107),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_301),
.Y(n_561)
);

BUFx10_ASAP7_75t_L g562 ( 
.A(n_193),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_246),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_441),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_199),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_177),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_139),
.B(n_183),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_29),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_16),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_62),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_195),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_222),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_239),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_414),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_305),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_210),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_295),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_135),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_219),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_23),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_429),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_204),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_71),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_50),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_37),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_203),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_143),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_160),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_162),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_36),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_3),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_387),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_415),
.Y(n_593)
);

BUFx10_ASAP7_75t_L g594 ( 
.A(n_122),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_223),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_366),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_21),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_247),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_252),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_262),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_166),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_271),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_182),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_301),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_338),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_45),
.Y(n_606)
);

INVxp67_ASAP7_75t_SL g607 ( 
.A(n_186),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_345),
.Y(n_608)
);

NOR2xp67_ASAP7_75t_L g609 ( 
.A(n_264),
.B(n_219),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_395),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_418),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_156),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_159),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_279),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_178),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_96),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_103),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_276),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_359),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_103),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_166),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_20),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_277),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_288),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_402),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_413),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_179),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_432),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_67),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_114),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_193),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_11),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_267),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_72),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_228),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_328),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_64),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_433),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_20),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_74),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_242),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_332),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_40),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_349),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_444),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_151),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_195),
.Y(n_647)
);

BUFx10_ASAP7_75t_L g648 ( 
.A(n_419),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_181),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_439),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_68),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_346),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_49),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_36),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_424),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_169),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_360),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_266),
.Y(n_658)
);

CKINVDCx16_ASAP7_75t_R g659 ( 
.A(n_306),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_246),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_240),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_202),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_226),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_70),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_211),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_75),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_295),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_183),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_109),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_370),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_286),
.B(n_9),
.Y(n_671)
);

CKINVDCx16_ASAP7_75t_R g672 ( 
.A(n_78),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_363),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_101),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_128),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_256),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_274),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_213),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_111),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_65),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_227),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_147),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_13),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_3),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_361),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_230),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_284),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_312),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_59),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_57),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_62),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_111),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_18),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_58),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_261),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_274),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_431),
.Y(n_697)
);

CKINVDCx14_ASAP7_75t_R g698 ( 
.A(n_120),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_326),
.Y(n_699)
);

BUFx2_ASAP7_75t_L g700 ( 
.A(n_172),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_79),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_108),
.B(n_390),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_391),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_45),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_442),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_58),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_374),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_443),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_74),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_417),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_135),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_16),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_362),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_365),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_188),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_158),
.Y(n_716)
);

BUFx2_ASAP7_75t_SL g717 ( 
.A(n_426),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_220),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_28),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_0),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_105),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_217),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_406),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_97),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_42),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_77),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_180),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_350),
.Y(n_728)
);

BUFx5_ASAP7_75t_L g729 ( 
.A(n_230),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_110),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_137),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_104),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_12),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_287),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_50),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_39),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_283),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_257),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_186),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_174),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_198),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_152),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_113),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_23),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_553),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_463),
.B(n_1),
.Y(n_746)
);

BUFx8_ASAP7_75t_L g747 ( 
.A(n_619),
.Y(n_747)
);

BUFx12f_ASAP7_75t_L g748 ( 
.A(n_648),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_560),
.Y(n_749)
);

XNOR2x2_ASAP7_75t_L g750 ( 
.A(n_451),
.B(n_671),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_560),
.B(n_2),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_698),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_752)
);

CKINVDCx16_ASAP7_75t_R g753 ( 
.A(n_480),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_520),
.B(n_4),
.Y(n_754)
);

INVx4_ASAP7_75t_L g755 ( 
.A(n_648),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_729),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_560),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_613),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_504),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_759)
);

INVx6_ASAP7_75t_L g760 ( 
.A(n_648),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_613),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_613),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_729),
.Y(n_763)
);

AND2x2_ASAP7_75t_SL g764 ( 
.A(n_482),
.B(n_316),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_622),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_468),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_536),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_729),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_468),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_468),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_622),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_700),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_729),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_622),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_729),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_489),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_548),
.B(n_7),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_656),
.B(n_8),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_656),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_656),
.Y(n_780)
);

INVx5_ASAP7_75t_L g781 ( 
.A(n_489),
.Y(n_781)
);

AND2x2_ASAP7_75t_SL g782 ( 
.A(n_528),
.B(n_318),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_SL g783 ( 
.A1(n_450),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_484),
.B(n_12),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_484),
.B(n_14),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_489),
.Y(n_786)
);

CKINVDCx11_ASAP7_75t_R g787 ( 
.A(n_450),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_542),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_452),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_573),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_552),
.A2(n_17),
.B1(n_14),
.B2(n_15),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_618),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_452),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_489),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_526),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_701),
.Y(n_796)
);

INVx4_ASAP7_75t_L g797 ( 
.A(n_473),
.Y(n_797)
);

NAND2xp33_ASAP7_75t_L g798 ( 
.A(n_519),
.B(n_320),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_659),
.A2(n_22),
.B1(n_19),
.B2(n_21),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_467),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_467),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_487),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_487),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_478),
.Y(n_804)
);

INVx5_ASAP7_75t_L g805 ( 
.A(n_526),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_701),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_701),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_493),
.Y(n_808)
);

OA21x2_ASAP7_75t_L g809 ( 
.A1(n_544),
.A2(n_322),
.B(n_321),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_672),
.B(n_19),
.Y(n_810)
);

OAI22x1_ASAP7_75t_R g811 ( 
.A1(n_555),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_449),
.B(n_24),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_497),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_497),
.Y(n_814)
);

INVx5_ASAP7_75t_L g815 ( 
.A(n_526),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_544),
.B(n_25),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_456),
.B(n_26),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_526),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_668),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_668),
.B(n_26),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_449),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_551),
.B(n_31),
.Y(n_822)
);

CKINVDCx6p67_ASAP7_75t_R g823 ( 
.A(n_473),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_458),
.B(n_32),
.Y(n_824)
);

OAI21x1_ASAP7_75t_L g825 ( 
.A1(n_545),
.A2(n_324),
.B(n_323),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_628),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_SL g827 ( 
.A(n_454),
.B(n_327),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_545),
.B(n_32),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_720),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_720),
.B(n_33),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_490),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_472),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_453),
.B(n_465),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_453),
.B(n_33),
.Y(n_834)
);

INVx4_ASAP7_75t_L g835 ( 
.A(n_628),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_465),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_490),
.B(n_34),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_564),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_555),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_564),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_543),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_527),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_481),
.A2(n_38),
.B1(n_35),
.B2(n_37),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_543),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_547),
.Y(n_845)
);

NAND2xp33_ASAP7_75t_L g846 ( 
.A(n_767),
.B(n_592),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_766),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_834),
.A2(n_447),
.B1(n_448),
.B2(n_446),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_751),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_755),
.B(n_521),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_751),
.B(n_596),
.Y(n_851)
);

AND2x6_ASAP7_75t_L g852 ( 
.A(n_778),
.B(n_605),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_756),
.Y(n_853)
);

AND2x6_ASAP7_75t_L g854 ( 
.A(n_778),
.B(n_605),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_756),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_778),
.Y(n_856)
);

AND2x2_ASAP7_75t_SL g857 ( 
.A(n_764),
.B(n_702),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_820),
.B(n_638),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_766),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_834),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_755),
.B(n_505),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_755),
.B(n_760),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_820),
.B(n_830),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_834),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_831),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_788),
.B(n_536),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_748),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_766),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_842),
.B(n_505),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_830),
.Y(n_870)
);

OR2x2_ASAP7_75t_L g871 ( 
.A(n_790),
.B(n_792),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_772),
.A2(n_481),
.B1(n_507),
.B2(n_506),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_830),
.B(n_650),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_779),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_779),
.Y(n_875)
);

AO22x2_ASAP7_75t_L g876 ( 
.A1(n_759),
.A2(n_607),
.B1(n_643),
.B2(n_539),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_766),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_779),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_807),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_763),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_804),
.B(n_536),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_807),
.Y(n_882)
);

AND3x1_ASAP7_75t_L g883 ( 
.A(n_843),
.B(n_459),
.C(n_457),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_842),
.B(n_506),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_769),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_769),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_804),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_814),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_814),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_753),
.B(n_808),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_768),
.B(n_657),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_768),
.Y(n_892)
);

OAI22x1_ASAP7_75t_L g893 ( 
.A1(n_832),
.A2(n_512),
.B1(n_556),
.B2(n_508),
.Y(n_893)
);

BUFx8_ASAP7_75t_SL g894 ( 
.A(n_839),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_797),
.B(n_508),
.Y(n_895)
);

NAND3xp33_ASAP7_75t_L g896 ( 
.A(n_754),
.B(n_743),
.C(n_556),
.Y(n_896)
);

AND2x6_ASAP7_75t_L g897 ( 
.A(n_746),
.B(n_670),
.Y(n_897)
);

BUFx10_ASAP7_75t_L g898 ( 
.A(n_764),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_749),
.Y(n_899)
);

AND2x6_ASAP7_75t_L g900 ( 
.A(n_746),
.B(n_670),
.Y(n_900)
);

NAND2xp33_ASAP7_75t_L g901 ( 
.A(n_767),
.B(n_608),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_773),
.Y(n_902)
);

AND2x6_ASAP7_75t_L g903 ( 
.A(n_822),
.B(n_813),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_757),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_758),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_773),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_775),
.B(n_673),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_782),
.A2(n_576),
.B1(n_579),
.B2(n_557),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_748),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_775),
.B(n_673),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_769),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_833),
.B(n_547),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_769),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_761),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_776),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_762),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_777),
.B(n_562),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_832),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_765),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_833),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_771),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_L g922 ( 
.A1(n_789),
.A2(n_470),
.B1(n_475),
.B2(n_462),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_774),
.Y(n_923)
);

OR2x6_ASAP7_75t_L g924 ( 
.A(n_783),
.B(n_609),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_780),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_796),
.B(n_714),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_782),
.A2(n_576),
.B1(n_579),
.B2(n_557),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_797),
.B(n_601),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_777),
.B(n_562),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_806),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_SL g931 ( 
.A(n_747),
.B(n_472),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_776),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_813),
.Y(n_933)
);

INVx8_ASAP7_75t_L g934 ( 
.A(n_822),
.Y(n_934)
);

NAND2xp33_ASAP7_75t_L g935 ( 
.A(n_819),
.B(n_611),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_810),
.B(n_562),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_810),
.B(n_594),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_823),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_826),
.B(n_620),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_776),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_826),
.B(n_714),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_829),
.Y(n_942)
);

INVx4_ASAP7_75t_L g943 ( 
.A(n_835),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_789),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_786),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_786),
.Y(n_946)
);

NAND3xp33_ASAP7_75t_L g947 ( 
.A(n_785),
.B(n_742),
.C(n_739),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_793),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_747),
.A2(n_635),
.B1(n_639),
.B2(n_620),
.Y(n_949)
);

BUFx10_ASAP7_75t_L g950 ( 
.A(n_817),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_786),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_835),
.B(n_635),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_823),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_793),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_800),
.Y(n_955)
);

INVx4_ASAP7_75t_L g956 ( 
.A(n_835),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_786),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_800),
.A2(n_483),
.B1(n_486),
.B2(n_476),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_801),
.B(n_460),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_801),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_802),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_802),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_809),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_803),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_841),
.B(n_594),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_803),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_794),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_838),
.A2(n_496),
.B1(n_498),
.B2(n_492),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_794),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_838),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_840),
.A2(n_784),
.B1(n_845),
.B2(n_844),
.Y(n_971)
);

OR2x6_ASAP7_75t_L g972 ( 
.A(n_791),
.B(n_717),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_836),
.B(n_640),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_794),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_794),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_840),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_812),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_781),
.B(n_464),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_818),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_784),
.A2(n_502),
.B1(n_503),
.B2(n_501),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_818),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_836),
.Y(n_982)
);

OR2x6_ASAP7_75t_L g983 ( 
.A(n_799),
.B(n_558),
.Y(n_983)
);

NAND3xp33_ASAP7_75t_L g984 ( 
.A(n_824),
.B(n_651),
.C(n_640),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_837),
.B(n_469),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_747),
.B(n_651),
.Y(n_986)
);

OAI22xp33_ASAP7_75t_L g987 ( 
.A1(n_745),
.A2(n_584),
.B1(n_597),
.B2(n_571),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_781),
.Y(n_988)
);

INVxp33_ASAP7_75t_L g989 ( 
.A(n_787),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_818),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_818),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_825),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_781),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_825),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_809),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_752),
.A2(n_674),
.B1(n_679),
.B2(n_658),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_805),
.B(n_471),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_816),
.Y(n_998)
);

INVxp67_ASAP7_75t_SL g999 ( 
.A(n_811),
.Y(n_999)
);

OAI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_821),
.A2(n_584),
.B1(n_597),
.B2(n_571),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_805),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_805),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_805),
.B(n_474),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_770),
.Y(n_1004)
);

AND2x2_ASAP7_75t_SL g1005 ( 
.A(n_827),
.B(n_558),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_828),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_815),
.B(n_479),
.Y(n_1007)
);

NOR2x1p5_ASAP7_75t_L g1008 ( 
.A(n_787),
.B(n_742),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_828),
.Y(n_1009)
);

OR2x6_ASAP7_75t_L g1010 ( 
.A(n_750),
.B(n_570),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_815),
.B(n_499),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_908),
.A2(n_534),
.B1(n_559),
.B2(n_477),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_869),
.B(n_454),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_871),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_977),
.B(n_461),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_SL g1016 ( 
.A1(n_857),
.A2(n_634),
.B1(n_641),
.B2(n_627),
.Y(n_1016)
);

NOR3xp33_ASAP7_75t_L g1017 ( 
.A(n_987),
.B(n_491),
.C(n_455),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_875),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_884),
.B(n_485),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_1010),
.A2(n_523),
.B(n_529),
.C(n_516),
.Y(n_1020)
);

AND2x2_ASAP7_75t_SL g1021 ( 
.A(n_1005),
.B(n_519),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_927),
.A2(n_534),
.B1(n_559),
.B2(n_477),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_875),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_860),
.A2(n_531),
.B1(n_537),
.B2(n_533),
.Y(n_1024)
);

OR2x6_ASAP7_75t_L g1025 ( 
.A(n_934),
.B(n_570),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_861),
.B(n_485),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_933),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_938),
.B(n_488),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_977),
.B(n_488),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_862),
.B(n_494),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_862),
.B(n_494),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_938),
.B(n_495),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_985),
.B(n_495),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_849),
.A2(n_541),
.B(n_550),
.C(n_540),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_982),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_944),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_917),
.B(n_594),
.Y(n_1037)
);

INVx8_ASAP7_75t_L g1038 ( 
.A(n_934),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_850),
.B(n_511),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_985),
.B(n_511),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_L g1041 ( 
.A(n_987),
.B(n_646),
.C(n_602),
.Y(n_1041)
);

NAND3xp33_ASAP7_75t_SL g1042 ( 
.A(n_980),
.B(n_679),
.C(n_674),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_864),
.A2(n_565),
.B1(n_566),
.B2(n_563),
.Y(n_1043)
);

INVx4_ASAP7_75t_L g1044 ( 
.A(n_953),
.Y(n_1044)
);

INVxp67_ASAP7_75t_L g1045 ( 
.A(n_865),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_929),
.B(n_724),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_936),
.B(n_724),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_937),
.B(n_725),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_953),
.B(n_568),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_1010),
.A2(n_569),
.B(n_575),
.C(n_572),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_920),
.B(n_947),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_895),
.B(n_546),
.Y(n_1052)
);

CKINVDCx6p67_ASAP7_75t_R g1053 ( 
.A(n_867),
.Y(n_1053)
);

OR2x6_ASAP7_75t_L g1054 ( 
.A(n_934),
.B(n_1008),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_897),
.B(n_554),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_897),
.B(n_574),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_881),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_897),
.B(n_574),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_856),
.A2(n_578),
.B1(n_580),
.B2(n_577),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_897),
.B(n_581),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_852),
.A2(n_583),
.B1(n_585),
.B2(n_582),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_948),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_848),
.B(n_581),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_866),
.B(n_681),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_L g1065 ( 
.A(n_896),
.B(n_691),
.C(n_681),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_863),
.A2(n_798),
.B(n_509),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_857),
.A2(n_636),
.B1(n_652),
.B2(n_626),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_887),
.B(n_655),
.Y(n_1068)
);

OR2x2_ASAP7_75t_L g1069 ( 
.A(n_865),
.B(n_691),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_965),
.A2(n_636),
.B1(n_652),
.B2(n_626),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_954),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_874),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_912),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_878),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_854),
.A2(n_615),
.B1(n_616),
.B2(n_589),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_928),
.B(n_707),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_879),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_963),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_848),
.B(n_707),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_882),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_912),
.Y(n_1081)
);

OAI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_1010),
.A2(n_728),
.B1(n_634),
.B2(n_641),
.Y(n_1082)
);

INVx8_ASAP7_75t_L g1083 ( 
.A(n_903),
.Y(n_1083)
);

BUFx12f_ASAP7_75t_L g1084 ( 
.A(n_918),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_854),
.A2(n_623),
.B1(n_624),
.B2(n_621),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_888),
.B(n_728),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_900),
.B(n_708),
.Y(n_1087)
);

AND2x6_ASAP7_75t_SL g1088 ( 
.A(n_924),
.B(n_839),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_1005),
.B(n_710),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_889),
.A2(n_706),
.B1(n_712),
.B2(n_694),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_890),
.B(n_694),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_955),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_960),
.Y(n_1093)
);

O2A1O1Ixp5_ASAP7_75t_L g1094 ( 
.A1(n_863),
.A2(n_500),
.B(n_513),
.C(n_510),
.Y(n_1094)
);

OR2x6_ASAP7_75t_L g1095 ( 
.A(n_972),
.B(n_591),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_854),
.A2(n_630),
.B1(n_631),
.B2(n_629),
.Y(n_1096)
);

AND2x6_ASAP7_75t_SL g1097 ( 
.A(n_924),
.B(n_567),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_984),
.B(n_632),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_939),
.B(n_514),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_952),
.B(n_706),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_998),
.B(n_466),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_950),
.B(n_517),
.Y(n_1102)
);

AND2x2_ASAP7_75t_SL g1103 ( 
.A(n_931),
.B(n_519),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_973),
.B(n_722),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_912),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_950),
.B(n_522),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_961),
.Y(n_1107)
);

BUFx5_ASAP7_75t_L g1108 ( 
.A(n_854),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_870),
.A2(n_637),
.B1(n_647),
.B2(n_633),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_962),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_903),
.A2(n_654),
.B1(n_660),
.B2(n_653),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_899),
.Y(n_1112)
);

INVx4_ASAP7_75t_L g1113 ( 
.A(n_903),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_903),
.B(n_739),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_992),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_964),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1006),
.B(n_743),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_1009),
.B(n_530),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_966),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_872),
.B(n_949),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_904),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_983),
.A2(n_662),
.B1(n_663),
.B2(n_661),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_970),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_983),
.A2(n_851),
.B(n_873),
.C(n_858),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_976),
.Y(n_1125)
);

XOR2x2_ASAP7_75t_L g1126 ( 
.A(n_883),
.B(n_627),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_858),
.B(n_515),
.Y(n_1127)
);

NOR3xp33_ASAP7_75t_L g1128 ( 
.A(n_1000),
.B(n_704),
.C(n_524),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_905),
.B(n_549),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_914),
.B(n_518),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_916),
.B(n_593),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_926),
.A2(n_665),
.B(n_666),
.C(n_664),
.Y(n_1132)
);

NOR2x1p5_ASAP7_75t_L g1133 ( 
.A(n_999),
.B(n_525),
.Y(n_1133)
);

INVxp67_ASAP7_75t_SL g1134 ( 
.A(n_994),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_919),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_921),
.B(n_532),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_986),
.B(n_893),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_983),
.B(n_535),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_996),
.A2(n_972),
.B1(n_971),
.B2(n_922),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_923),
.B(n_538),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_898),
.A2(n_590),
.B1(n_595),
.B2(n_586),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_925),
.B(n_598),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_930),
.A2(n_669),
.B1(n_675),
.B2(n_667),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_898),
.A2(n_599),
.B1(n_603),
.B2(n_600),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_942),
.B(n_606),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_972),
.B(n_612),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_846),
.B(n_625),
.Y(n_1147)
);

NAND3xp33_ASAP7_75t_SL g1148 ( 
.A(n_922),
.B(n_617),
.C(n_649),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_959),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_943),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_959),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_926),
.A2(n_677),
.B1(n_682),
.B2(n_676),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_935),
.B(n_642),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_901),
.B(n_644),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_958),
.B(n_649),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_956),
.B(n_645),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_958),
.B(n_678),
.Y(n_1157)
);

INVxp67_ASAP7_75t_L g1158 ( 
.A(n_1011),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_968),
.B(n_685),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_941),
.B(n_697),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1002),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_894),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_968),
.B(n_699),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_891),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_894),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1002),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_891),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_941),
.B(n_703),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_995),
.B(n_705),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_853),
.B(n_713),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_924),
.B(n_683),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_907),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_855),
.B(n_723),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_876),
.B(n_680),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_876),
.A2(n_684),
.B1(n_687),
.B2(n_686),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_876),
.A2(n_690),
.B1(n_696),
.B2(n_689),
.Y(n_1176)
);

INVx5_ASAP7_75t_L g1177 ( 
.A(n_988),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_978),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_989),
.Y(n_1179)
);

AND2x4_ASAP7_75t_SL g1180 ( 
.A(n_989),
.B(n_680),
.Y(n_1180)
);

OAI221xp5_ASAP7_75t_L g1181 ( 
.A1(n_910),
.A2(n_716),
.B1(n_718),
.B2(n_715),
.C(n_709),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_880),
.B(n_591),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_892),
.B(n_604),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_902),
.B(n_604),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_910),
.A2(n_721),
.B1(n_726),
.B2(n_719),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_902),
.A2(n_731),
.B1(n_732),
.B2(n_727),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_906),
.B(n_614),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1000),
.A2(n_736),
.B1(n_738),
.B2(n_733),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1007),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_978),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_997),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1001),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_997),
.B(n_741),
.Y(n_1193)
);

AND2x6_ASAP7_75t_SL g1194 ( 
.A(n_1003),
.B(n_744),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_993),
.B(n_693),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_911),
.B(n_693),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_913),
.B(n_737),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_913),
.B(n_688),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_915),
.A2(n_734),
.B1(n_735),
.B2(n_688),
.Y(n_1199)
);

BUFx12f_ASAP7_75t_L g1200 ( 
.A(n_847),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_915),
.A2(n_735),
.B1(n_740),
.B2(n_734),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_932),
.B(n_561),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_940),
.B(n_561),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_847),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_940),
.B(n_587),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_945),
.Y(n_1206)
);

OR2x4_ASAP7_75t_L g1207 ( 
.A(n_847),
.B(n_588),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_945),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_946),
.A2(n_692),
.B1(n_695),
.B2(n_588),
.Y(n_1209)
);

NAND3xp33_ASAP7_75t_SL g1210 ( 
.A(n_951),
.B(n_740),
.C(n_957),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_SL g1211 ( 
.A1(n_859),
.A2(n_692),
.B1(n_711),
.B2(n_695),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_969),
.B(n_692),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_969),
.Y(n_1213)
);

INVx4_ASAP7_75t_L g1214 ( 
.A(n_859),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_974),
.B(n_695),
.Y(n_1215)
);

INVxp67_ASAP7_75t_L g1216 ( 
.A(n_974),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_979),
.B(n_695),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1112),
.Y(n_1218)
);

BUFx4f_ASAP7_75t_L g1219 ( 
.A(n_1038),
.Y(n_1219)
);

NAND3xp33_ASAP7_75t_L g1220 ( 
.A(n_1128),
.B(n_730),
.C(n_610),
.Y(n_1220)
);

NOR3xp33_ASAP7_75t_L g1221 ( 
.A(n_1148),
.B(n_981),
.C(n_979),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1034),
.A2(n_981),
.B(n_991),
.C(n_1004),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1121),
.B(n_730),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1014),
.B(n_730),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1014),
.B(n_35),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1135),
.B(n_1124),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1057),
.B(n_38),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1051),
.B(n_39),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1051),
.B(n_41),
.Y(n_1229)
);

CKINVDCx10_ASAP7_75t_R g1230 ( 
.A(n_1054),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1073),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1155),
.B(n_42),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1195),
.Y(n_1233)
);

AO32x1_ASAP7_75t_L g1234 ( 
.A1(n_1139),
.A2(n_795),
.A3(n_770),
.B1(n_815),
.B2(n_859),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1120),
.A2(n_815),
.B1(n_795),
.B2(n_770),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1015),
.B(n_1029),
.Y(n_1236)
);

OR2x6_ASAP7_75t_SL g1237 ( 
.A(n_1012),
.B(n_1022),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1083),
.Y(n_1238)
);

BUFx2_ASAP7_75t_SL g1239 ( 
.A(n_1044),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1038),
.Y(n_1240)
);

BUFx2_ASAP7_75t_SL g1241 ( 
.A(n_1044),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1033),
.B(n_43),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1123),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1157),
.B(n_43),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1040),
.B(n_44),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1038),
.Y(n_1246)
);

AND2x6_ASAP7_75t_L g1247 ( 
.A(n_1083),
.B(n_868),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1078),
.A2(n_877),
.B(n_868),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_1201),
.B(n_44),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1104),
.B(n_46),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1039),
.B(n_46),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1021),
.A2(n_885),
.B1(n_886),
.B2(n_877),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1039),
.B(n_47),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1099),
.A2(n_1160),
.B(n_1168),
.C(n_1094),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1069),
.B(n_47),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1025),
.B(n_48),
.Y(n_1256)
);

A2O1A1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1099),
.A2(n_886),
.B(n_967),
.C(n_885),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1064),
.A2(n_967),
.B1(n_975),
.B2(n_886),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1025),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1091),
.B(n_48),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1053),
.Y(n_1261)
);

OR2x6_ASAP7_75t_L g1262 ( 
.A(n_1025),
.B(n_49),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1046),
.B(n_51),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1049),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1083),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1037),
.A2(n_990),
.B1(n_975),
.B2(n_54),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1162),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1047),
.B(n_52),
.Y(n_1268)
);

AO22x1_ASAP7_75t_L g1269 ( 
.A1(n_1128),
.A2(n_56),
.B1(n_53),
.B2(n_55),
.Y(n_1269)
);

CKINVDCx16_ASAP7_75t_R g1270 ( 
.A(n_1165),
.Y(n_1270)
);

NAND2x1p5_ASAP7_75t_L g1271 ( 
.A(n_1103),
.B(n_990),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1115),
.A2(n_990),
.B(n_331),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1048),
.B(n_60),
.Y(n_1273)
);

NOR2xp67_ASAP7_75t_L g1274 ( 
.A(n_1188),
.B(n_60),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1150),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1013),
.B(n_61),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1019),
.B(n_63),
.Y(n_1277)
);

CKINVDCx10_ASAP7_75t_R g1278 ( 
.A(n_1054),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1177),
.Y(n_1279)
);

O2A1O1Ixp5_ASAP7_75t_L g1280 ( 
.A1(n_1089),
.A2(n_334),
.B(n_335),
.C(n_330),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1081),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1084),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1098),
.B(n_69),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1095),
.B(n_69),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1036),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1108),
.B(n_71),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1141),
.B(n_72),
.Y(n_1287)
);

NOR2xp67_ASAP7_75t_L g1288 ( 
.A(n_1148),
.B(n_73),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1066),
.A2(n_341),
.B(n_340),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1021),
.A2(n_76),
.B1(n_73),
.B2(n_75),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1144),
.B(n_76),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1052),
.B(n_77),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1111),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_1293)
);

INVx2_ASAP7_75t_SL g1294 ( 
.A(n_1049),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1132),
.A2(n_83),
.B(n_80),
.C(n_82),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1042),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_1296)
);

AO21x1_ASAP7_75t_L g1297 ( 
.A1(n_1205),
.A2(n_84),
.B(n_85),
.Y(n_1297)
);

AOI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1189),
.A2(n_348),
.B(n_347),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1158),
.A2(n_353),
.B(n_351),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1111),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1052),
.B(n_86),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1102),
.B(n_87),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1117),
.A2(n_355),
.B(n_354),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1207),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1102),
.B(n_88),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1108),
.B(n_89),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1105),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1106),
.B(n_89),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1137),
.B(n_1146),
.Y(n_1309)
);

OAI22x1_ASAP7_75t_L g1310 ( 
.A1(n_1067),
.A2(n_94),
.B1(n_90),
.B2(n_92),
.Y(n_1310)
);

AOI221xp5_ASAP7_75t_L g1311 ( 
.A1(n_1017),
.A2(n_95),
.B1(n_92),
.B2(n_94),
.C(n_96),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1076),
.B(n_95),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1160),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1062),
.Y(n_1314)
);

INVx4_ASAP7_75t_L g1315 ( 
.A(n_1177),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1071),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1068),
.B(n_98),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1072),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1086),
.B(n_99),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1164),
.A2(n_1172),
.B(n_1167),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1074),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1086),
.B(n_100),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1100),
.A2(n_368),
.B(n_364),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1138),
.B(n_102),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1207),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1090),
.B(n_104),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1024),
.B(n_105),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1042),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1092),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1024),
.B(n_1043),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1070),
.B(n_106),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1200),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_SL g1333 ( 
.A(n_1103),
.B(n_109),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1043),
.B(n_110),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1198),
.B(n_112),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1030),
.A2(n_380),
.B(n_378),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1031),
.A2(n_1156),
.B(n_1080),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1108),
.B(n_113),
.Y(n_1338)
);

AOI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1171),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1109),
.B(n_115),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1122),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1093),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1077),
.A2(n_383),
.B(n_382),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1107),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1017),
.A2(n_120),
.B(n_118),
.C(n_119),
.Y(n_1345)
);

O2A1O1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1041),
.A2(n_122),
.B(n_119),
.C(n_121),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1109),
.B(n_121),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1180),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1179),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1059),
.B(n_124),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1055),
.A2(n_392),
.B(n_389),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1056),
.A2(n_1060),
.B(n_1058),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1059),
.B(n_1026),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1035),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1028),
.B(n_125),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1032),
.B(n_126),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1087),
.A2(n_404),
.B(n_397),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1095),
.B(n_127),
.Y(n_1358)
);

AND2x6_ASAP7_75t_L g1359 ( 
.A(n_1149),
.B(n_409),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_SL g1360 ( 
.A1(n_1095),
.A2(n_411),
.B(n_410),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1122),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_1361)
);

A2O1A1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1168),
.A2(n_132),
.B(n_129),
.C(n_131),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1171),
.A2(n_133),
.B1(n_134),
.B2(n_136),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1063),
.B(n_134),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1079),
.B(n_136),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1182),
.Y(n_1366)
);

OA22x2_ASAP7_75t_L g1367 ( 
.A1(n_1175),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1054),
.B(n_138),
.Y(n_1368)
);

O2A1O1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1041),
.A2(n_141),
.B(n_142),
.C(n_143),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1129),
.B(n_141),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1129),
.B(n_144),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1110),
.Y(n_1372)
);

CKINVDCx10_ASAP7_75t_R g1373 ( 
.A(n_1088),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1145),
.B(n_144),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1163),
.B(n_145),
.Y(n_1375)
);

O2A1O1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1020),
.A2(n_145),
.B(n_146),
.C(n_148),
.Y(n_1376)
);

INVx4_ASAP7_75t_SL g1377 ( 
.A(n_1192),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1061),
.A2(n_421),
.B(n_420),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1133),
.Y(n_1379)
);

AND2x6_ASAP7_75t_L g1380 ( 
.A(n_1151),
.B(n_422),
.Y(n_1380)
);

BUFx4f_ASAP7_75t_L g1381 ( 
.A(n_1027),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1183),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1131),
.B(n_146),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1184),
.Y(n_1384)
);

NAND3xp33_ASAP7_75t_L g1385 ( 
.A(n_1065),
.B(n_148),
.C(n_149),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1131),
.B(n_149),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1050),
.A2(n_150),
.B(n_151),
.C(n_152),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1177),
.Y(n_1388)
);

OAI21xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1061),
.A2(n_154),
.B(n_155),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1075),
.A2(n_430),
.B(n_428),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1116),
.B(n_155),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1174),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1199),
.Y(n_1393)
);

OAI21xp33_ASAP7_75t_SL g1394 ( 
.A1(n_1075),
.A2(n_157),
.B(n_159),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1119),
.B(n_160),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1125),
.B(n_161),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1193),
.B(n_161),
.Y(n_1397)
);

INVx5_ASAP7_75t_L g1398 ( 
.A(n_1192),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1114),
.B(n_163),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1187),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1210),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1016),
.B(n_164),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1193),
.B(n_167),
.Y(n_1403)
);

INVxp67_ASAP7_75t_SL g1404 ( 
.A(n_1082),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1085),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_1405)
);

BUFx12f_ASAP7_75t_L g1406 ( 
.A(n_1097),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1147),
.B(n_168),
.Y(n_1407)
);

O2A1O1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1159),
.A2(n_170),
.B(n_171),
.C(n_172),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1154),
.B(n_171),
.Y(n_1409)
);

NAND3xp33_ASAP7_75t_L g1410 ( 
.A(n_1085),
.B(n_1096),
.C(n_1143),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1130),
.B(n_1136),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1127),
.A2(n_436),
.B(n_434),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1118),
.A2(n_437),
.B(n_174),
.Y(n_1413)
);

CKINVDCx16_ASAP7_75t_R g1414 ( 
.A(n_1176),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1082),
.Y(n_1415)
);

INVxp67_ASAP7_75t_L g1416 ( 
.A(n_1140),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1142),
.B(n_173),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1101),
.B(n_315),
.Y(n_1418)
);

AOI22x1_ASAP7_75t_L g1419 ( 
.A1(n_1214),
.A2(n_175),
.B1(n_176),
.B2(n_178),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1096),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1181),
.A2(n_1152),
.B1(n_1186),
.B2(n_1143),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1152),
.A2(n_184),
.B1(n_185),
.B2(n_187),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1018),
.A2(n_184),
.B(n_185),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1177),
.B(n_187),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1185),
.B(n_188),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1016),
.B(n_189),
.Y(n_1426)
);

NAND3xp33_ASAP7_75t_L g1427 ( 
.A(n_1186),
.B(n_190),
.C(n_191),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1023),
.A2(n_190),
.B(n_191),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_SL g1429 ( 
.A(n_1214),
.B(n_192),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1161),
.A2(n_194),
.B(n_196),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1178),
.B(n_194),
.Y(n_1431)
);

OR2x6_ASAP7_75t_L g1432 ( 
.A(n_1190),
.B(n_1191),
.Y(n_1432)
);

O2A1O1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1170),
.A2(n_196),
.B(n_197),
.C(n_198),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1173),
.A2(n_197),
.B(n_199),
.C(n_200),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1153),
.B(n_200),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1166),
.A2(n_201),
.B(n_203),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1194),
.B(n_205),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1211),
.B(n_206),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1211),
.B(n_207),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1196),
.B(n_207),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1197),
.A2(n_208),
.B1(n_209),
.B2(n_211),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1208),
.B(n_208),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1209),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1216),
.A2(n_215),
.B(n_216),
.Y(n_1444)
);

AOI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1202),
.A2(n_216),
.B(n_218),
.Y(n_1445)
);

OAI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1262),
.A2(n_1126),
.B1(n_1215),
.B2(n_1212),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1332),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1332),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1218),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1285),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1262),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1414),
.B(n_220),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1393),
.B(n_221),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1299),
.A2(n_1217),
.B(n_1203),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_SL g1455 ( 
.A(n_1219),
.B(n_1204),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1219),
.B(n_1206),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1240),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1262),
.Y(n_1458)
);

BUFx4f_ASAP7_75t_L g1459 ( 
.A(n_1332),
.Y(n_1459)
);

AO31x2_ASAP7_75t_L g1460 ( 
.A1(n_1297),
.A2(n_1213),
.A3(n_223),
.B(n_224),
.Y(n_1460)
);

AO21x1_ASAP7_75t_L g1461 ( 
.A1(n_1290),
.A2(n_222),
.B(n_224),
.Y(n_1461)
);

NOR2x1_ASAP7_75t_R g1462 ( 
.A(n_1261),
.B(n_1348),
.Y(n_1462)
);

O2A1O1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1353),
.A2(n_225),
.B(n_226),
.C(n_229),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1415),
.A2(n_229),
.B1(n_231),
.B2(n_232),
.Y(n_1464)
);

AO32x2_ASAP7_75t_L g1465 ( 
.A1(n_1293),
.A2(n_233),
.A3(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1230),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1318),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1320),
.A2(n_234),
.B(n_235),
.Y(n_1468)
);

A2O1A1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1302),
.A2(n_1308),
.B(n_1305),
.C(n_1374),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1315),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1278),
.Y(n_1471)
);

A2O1A1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1417),
.A2(n_237),
.B(n_238),
.C(n_240),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1404),
.B(n_237),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1248),
.A2(n_241),
.B(n_243),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1246),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1321),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1410),
.A2(n_243),
.B(n_244),
.Y(n_1477)
);

BUFx10_ASAP7_75t_L g1478 ( 
.A(n_1256),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1226),
.A2(n_245),
.B(n_247),
.Y(n_1479)
);

O2A1O1Ixp33_ASAP7_75t_SL g1480 ( 
.A1(n_1276),
.A2(n_248),
.B(n_250),
.C(n_251),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1294),
.B(n_253),
.Y(n_1481)
);

INVxp67_ASAP7_75t_SL g1482 ( 
.A(n_1256),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1284),
.Y(n_1483)
);

CKINVDCx6p67_ASAP7_75t_R g1484 ( 
.A(n_1282),
.Y(n_1484)
);

INVx2_ASAP7_75t_SL g1485 ( 
.A(n_1267),
.Y(n_1485)
);

AO31x2_ASAP7_75t_L g1486 ( 
.A1(n_1257),
.A2(n_1252),
.A3(n_1228),
.B(n_1229),
.Y(n_1486)
);

O2A1O1Ixp33_ASAP7_75t_SL g1487 ( 
.A1(n_1277),
.A2(n_254),
.B(n_255),
.C(n_257),
.Y(n_1487)
);

AO31x2_ASAP7_75t_L g1488 ( 
.A1(n_1252),
.A2(n_258),
.A3(n_259),
.B(n_260),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1330),
.B(n_259),
.Y(n_1489)
);

AO31x2_ASAP7_75t_L g1490 ( 
.A1(n_1229),
.A2(n_1223),
.A3(n_1386),
.B(n_1383),
.Y(n_1490)
);

INVx1_ASAP7_75t_SL g1491 ( 
.A(n_1264),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_1284),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1314),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1354),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1366),
.A2(n_269),
.B(n_270),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1272),
.A2(n_270),
.B(n_271),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1368),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1333),
.B(n_273),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1382),
.A2(n_273),
.B(n_275),
.Y(n_1499)
);

INVxp67_ASAP7_75t_L g1500 ( 
.A(n_1225),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1316),
.Y(n_1501)
);

A2O1A1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1317),
.A2(n_275),
.B(n_278),
.C(n_279),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1384),
.A2(n_278),
.B(n_280),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1368),
.B(n_280),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1400),
.A2(n_281),
.B(n_282),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1416),
.B(n_281),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1329),
.Y(n_1507)
);

INVx6_ASAP7_75t_SL g1508 ( 
.A(n_1432),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1421),
.B(n_284),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1309),
.B(n_285),
.Y(n_1510)
);

CKINVDCx14_ASAP7_75t_R g1511 ( 
.A(n_1349),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1342),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1344),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1407),
.A2(n_286),
.B1(n_287),
.B2(n_290),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1372),
.Y(n_1515)
);

AO21x2_ASAP7_75t_L g1516 ( 
.A1(n_1289),
.A2(n_291),
.B(n_292),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1232),
.B(n_291),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1244),
.B(n_292),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1281),
.B(n_293),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1391),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1407),
.A2(n_294),
.B1(n_296),
.B2(n_297),
.Y(n_1521)
);

AO31x2_ASAP7_75t_L g1522 ( 
.A1(n_1223),
.A2(n_296),
.A3(n_297),
.B(n_298),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1307),
.B(n_298),
.Y(n_1523)
);

AOI21xp33_ASAP7_75t_L g1524 ( 
.A1(n_1251),
.A2(n_299),
.B(n_300),
.Y(n_1524)
);

AO31x2_ASAP7_75t_L g1525 ( 
.A1(n_1383),
.A2(n_302),
.A3(n_303),
.B(n_304),
.Y(n_1525)
);

BUFx4f_ASAP7_75t_L g1526 ( 
.A(n_1406),
.Y(n_1526)
);

OAI22x1_ASAP7_75t_L g1527 ( 
.A1(n_1402),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1233),
.B(n_305),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1375),
.A2(n_306),
.B(n_307),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1391),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1263),
.B(n_307),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1260),
.B(n_308),
.Y(n_1532)
);

OR2x6_ASAP7_75t_L g1533 ( 
.A(n_1239),
.B(n_315),
.Y(n_1533)
);

OAI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1375),
.A2(n_308),
.B(n_309),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1397),
.A2(n_309),
.B(n_310),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_SL g1536 ( 
.A(n_1429),
.B(n_310),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1259),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1237),
.B(n_311),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1395),
.Y(n_1539)
);

AO31x2_ASAP7_75t_L g1540 ( 
.A1(n_1434),
.A2(n_313),
.A3(n_314),
.B(n_1351),
.Y(n_1540)
);

CKINVDCx8_ASAP7_75t_R g1541 ( 
.A(n_1373),
.Y(n_1541)
);

CKINVDCx9p33_ASAP7_75t_R g1542 ( 
.A(n_1358),
.Y(n_1542)
);

AOI221x1_ASAP7_75t_L g1543 ( 
.A1(n_1310),
.A2(n_1390),
.B1(n_1378),
.B2(n_1293),
.C(n_1300),
.Y(n_1543)
);

CKINVDCx11_ASAP7_75t_R g1544 ( 
.A(n_1270),
.Y(n_1544)
);

OAI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1249),
.A2(n_1274),
.B1(n_1288),
.B2(n_1367),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1242),
.A2(n_1245),
.B(n_1253),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1324),
.B(n_1319),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_SL g1548 ( 
.A(n_1271),
.B(n_1378),
.Y(n_1548)
);

INVx8_ASAP7_75t_L g1549 ( 
.A(n_1247),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1395),
.Y(n_1550)
);

AO31x2_ASAP7_75t_L g1551 ( 
.A1(n_1357),
.A2(n_1336),
.A3(n_1313),
.B(n_1362),
.Y(n_1551)
);

AOI221x1_ASAP7_75t_L g1552 ( 
.A1(n_1390),
.A2(n_1300),
.B1(n_1422),
.B2(n_1385),
.C(n_1341),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1241),
.Y(n_1553)
);

O2A1O1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1387),
.A2(n_1369),
.B(n_1346),
.C(n_1345),
.Y(n_1554)
);

AO21x2_ASAP7_75t_L g1555 ( 
.A1(n_1445),
.A2(n_1234),
.B(n_1235),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1396),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1331),
.B(n_1426),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1398),
.Y(n_1558)
);

AO31x2_ASAP7_75t_L g1559 ( 
.A1(n_1441),
.A2(n_1422),
.A3(n_1396),
.B(n_1323),
.Y(n_1559)
);

A2O1A1Ixp33_ASAP7_75t_L g1560 ( 
.A1(n_1268),
.A2(n_1273),
.B(n_1255),
.C(n_1409),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1389),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1326),
.B(n_1322),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1275),
.Y(n_1563)
);

OA21x2_ASAP7_75t_L g1564 ( 
.A1(n_1280),
.A2(n_1303),
.B(n_1412),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1292),
.A2(n_1312),
.B(n_1301),
.Y(n_1565)
);

CKINVDCx12_ASAP7_75t_R g1566 ( 
.A(n_1432),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1335),
.Y(n_1567)
);

A2O1A1Ixp33_ASAP7_75t_L g1568 ( 
.A1(n_1409),
.A2(n_1403),
.B(n_1397),
.C(n_1295),
.Y(n_1568)
);

A2O1A1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1403),
.A2(n_1370),
.B(n_1371),
.C(n_1222),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_1227),
.Y(n_1570)
);

BUFx10_ASAP7_75t_L g1571 ( 
.A(n_1355),
.Y(n_1571)
);

AOI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1287),
.A2(n_1291),
.B1(n_1347),
.B2(n_1334),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1243),
.B(n_1250),
.Y(n_1573)
);

AO21x1_ASAP7_75t_L g1574 ( 
.A1(n_1286),
.A2(n_1338),
.B(n_1306),
.Y(n_1574)
);

NOR2x1_ASAP7_75t_L g1575 ( 
.A(n_1427),
.B(n_1437),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_1341),
.Y(n_1576)
);

O2A1O1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1327),
.A2(n_1340),
.B(n_1350),
.C(n_1376),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1399),
.A2(n_1440),
.B(n_1364),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1224),
.B(n_1379),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1392),
.Y(n_1580)
);

AND2x2_ASAP7_75t_SL g1581 ( 
.A(n_1381),
.B(n_1296),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1283),
.B(n_1425),
.Y(n_1582)
);

INVx3_ASAP7_75t_SL g1583 ( 
.A(n_1304),
.Y(n_1583)
);

AOI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1418),
.A2(n_1356),
.B1(n_1361),
.B2(n_1435),
.Y(n_1584)
);

O2A1O1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1361),
.A2(n_1425),
.B(n_1394),
.C(n_1405),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1365),
.A2(n_1432),
.B(n_1442),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1231),
.B(n_1381),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1367),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1431),
.Y(n_1589)
);

INVx3_ASAP7_75t_SL g1590 ( 
.A(n_1325),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1419),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1339),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1405),
.A2(n_1420),
.B1(n_1266),
.B2(n_1363),
.Y(n_1593)
);

A2O1A1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1408),
.A2(n_1433),
.B(n_1444),
.C(n_1423),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1271),
.A2(n_1328),
.B1(n_1401),
.B2(n_1420),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1311),
.B(n_1428),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1258),
.A2(n_1234),
.B(n_1424),
.Y(n_1597)
);

AO21x1_ASAP7_75t_L g1598 ( 
.A1(n_1343),
.A2(n_1441),
.B(n_1430),
.Y(n_1598)
);

AOI221x1_ASAP7_75t_L g1599 ( 
.A1(n_1436),
.A2(n_1221),
.B1(n_1360),
.B2(n_1439),
.C(n_1438),
.Y(n_1599)
);

BUFx12f_ASAP7_75t_L g1600 ( 
.A(n_1238),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1269),
.A2(n_1443),
.B1(n_1279),
.B2(n_1388),
.Y(n_1601)
);

AO31x2_ASAP7_75t_L g1602 ( 
.A1(n_1234),
.A2(n_1413),
.A3(n_1380),
.B(n_1359),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_SL g1603 ( 
.A(n_1265),
.B(n_1359),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1359),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1377),
.A2(n_1359),
.B(n_1380),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1380),
.Y(n_1606)
);

BUFx10_ASAP7_75t_L g1607 ( 
.A(n_1380),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1247),
.B(n_1330),
.Y(n_1608)
);

NAND3xp33_ASAP7_75t_L g1609 ( 
.A(n_1220),
.B(n_1305),
.C(n_1302),
.Y(n_1609)
);

NAND3xp33_ASAP7_75t_L g1610 ( 
.A(n_1220),
.B(n_1305),
.C(n_1302),
.Y(n_1610)
);

AOI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1252),
.A2(n_1223),
.B(n_1298),
.Y(n_1611)
);

AO21x2_ASAP7_75t_L g1612 ( 
.A1(n_1299),
.A2(n_1257),
.B(n_1289),
.Y(n_1612)
);

AO31x2_ASAP7_75t_L g1613 ( 
.A1(n_1297),
.A2(n_1257),
.A3(n_1169),
.B(n_1254),
.Y(n_1613)
);

CKINVDCx8_ASAP7_75t_R g1614 ( 
.A(n_1230),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1230),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1294),
.B(n_1264),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1393),
.B(n_1014),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1218),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1404),
.A2(n_1045),
.B1(n_832),
.B2(n_1022),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1218),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1404),
.B(n_1014),
.Y(n_1621)
);

A2O1A1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1411),
.A2(n_1337),
.B(n_1254),
.C(n_1236),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1219),
.B(n_1045),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1330),
.B(n_1218),
.Y(n_1624)
);

INVxp67_ASAP7_75t_SL g1625 ( 
.A(n_1219),
.Y(n_1625)
);

NAND3xp33_ASAP7_75t_L g1626 ( 
.A(n_1220),
.B(n_1305),
.C(n_1302),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1330),
.B(n_1218),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_SL g1628 ( 
.A(n_1333),
.B(n_1113),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1262),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1332),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1218),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1393),
.B(n_1014),
.Y(n_1632)
);

OA21x2_ASAP7_75t_L g1633 ( 
.A1(n_1299),
.A2(n_825),
.B(n_1289),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_SL g1634 ( 
.A1(n_1414),
.A2(n_1016),
.B1(n_839),
.B2(n_1010),
.Y(n_1634)
);

AO31x2_ASAP7_75t_L g1635 ( 
.A1(n_1297),
.A2(n_1257),
.A3(n_1169),
.B(n_1254),
.Y(n_1635)
);

INVx5_ASAP7_75t_L g1636 ( 
.A(n_1332),
.Y(n_1636)
);

INVx3_ASAP7_75t_SL g1637 ( 
.A(n_1332),
.Y(n_1637)
);

O2A1O1Ixp33_ASAP7_75t_L g1638 ( 
.A1(n_1353),
.A2(n_1236),
.B(n_1387),
.C(n_1254),
.Y(n_1638)
);

AO21x2_ASAP7_75t_L g1639 ( 
.A1(n_1299),
.A2(n_1257),
.B(n_1289),
.Y(n_1639)
);

BUFx6f_ASAP7_75t_L g1640 ( 
.A(n_1332),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1332),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1294),
.B(n_1264),
.Y(n_1642)
);

BUFx2_ASAP7_75t_R g1643 ( 
.A(n_1282),
.Y(n_1643)
);

AO31x2_ASAP7_75t_L g1644 ( 
.A1(n_1297),
.A2(n_1257),
.A3(n_1169),
.B(n_1254),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1218),
.Y(n_1645)
);

AOI21xp33_ASAP7_75t_L g1646 ( 
.A1(n_1302),
.A2(n_1021),
.B(n_1305),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1330),
.B(n_1218),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1404),
.B(n_1014),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_1332),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1404),
.A2(n_1045),
.B1(n_832),
.B2(n_1022),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_SL g1651 ( 
.A1(n_1378),
.A2(n_1390),
.B(n_1299),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1330),
.B(n_1218),
.Y(n_1652)
);

AO31x2_ASAP7_75t_L g1653 ( 
.A1(n_1297),
.A2(n_1257),
.A3(n_1169),
.B(n_1254),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1337),
.A2(n_1134),
.B(n_1236),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1218),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1332),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1337),
.A2(n_1134),
.B(n_1236),
.Y(n_1657)
);

NAND3x1_ASAP7_75t_L g1658 ( 
.A(n_1402),
.B(n_1128),
.C(n_1041),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1337),
.A2(n_1134),
.B(n_1236),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1218),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1330),
.B(n_1218),
.Y(n_1661)
);

INVx5_ASAP7_75t_L g1662 ( 
.A(n_1332),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1330),
.B(n_1218),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1330),
.B(n_1218),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1218),
.Y(n_1665)
);

AO31x2_ASAP7_75t_L g1666 ( 
.A1(n_1297),
.A2(n_1257),
.A3(n_1169),
.B(n_1254),
.Y(n_1666)
);

NAND2x1p5_ASAP7_75t_L g1667 ( 
.A(n_1219),
.B(n_1332),
.Y(n_1667)
);

NOR2xp67_ASAP7_75t_L g1668 ( 
.A(n_1332),
.B(n_909),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1404),
.A2(n_1045),
.B1(n_832),
.B2(n_1022),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1337),
.A2(n_1134),
.B(n_1236),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1294),
.B(n_1264),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1337),
.A2(n_1134),
.B(n_1236),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1218),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1393),
.B(n_1014),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1330),
.B(n_1218),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1218),
.Y(n_1676)
);

AO21x1_ASAP7_75t_L g1677 ( 
.A1(n_1299),
.A2(n_1290),
.B(n_1378),
.Y(n_1677)
);

AOI21x1_ASAP7_75t_L g1678 ( 
.A1(n_1252),
.A2(n_1223),
.B(n_1298),
.Y(n_1678)
);

O2A1O1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1353),
.A2(n_1236),
.B(n_1387),
.C(n_1254),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1332),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1230),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1337),
.A2(n_1134),
.B(n_1236),
.Y(n_1682)
);

O2A1O1Ixp33_ASAP7_75t_L g1683 ( 
.A1(n_1353),
.A2(n_1236),
.B(n_1387),
.C(n_1254),
.Y(n_1683)
);

OAI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1254),
.A2(n_1352),
.B(n_1337),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_R g1685 ( 
.A(n_1230),
.B(n_1278),
.Y(n_1685)
);

CKINVDCx20_ASAP7_75t_R g1686 ( 
.A(n_1261),
.Y(n_1686)
);

OAI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1262),
.A2(n_832),
.B1(n_931),
.B2(n_1067),
.Y(n_1687)
);

O2A1O1Ixp33_ASAP7_75t_L g1688 ( 
.A1(n_1353),
.A2(n_1236),
.B(n_1387),
.C(n_1254),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1240),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1330),
.B(n_1218),
.Y(n_1690)
);

OAI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1254),
.A2(n_1352),
.B(n_1337),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1218),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1393),
.B(n_1014),
.Y(n_1693)
);

NAND2x1p5_ASAP7_75t_L g1694 ( 
.A(n_1219),
.B(n_1332),
.Y(n_1694)
);

CKINVDCx20_ASAP7_75t_R g1695 ( 
.A(n_1261),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1218),
.Y(n_1696)
);

AO21x1_ASAP7_75t_L g1697 ( 
.A1(n_1299),
.A2(n_1290),
.B(n_1378),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_1262),
.Y(n_1698)
);

AO31x2_ASAP7_75t_L g1699 ( 
.A1(n_1297),
.A2(n_1257),
.A3(n_1169),
.B(n_1254),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1218),
.Y(n_1700)
);

INVx4_ASAP7_75t_L g1701 ( 
.A(n_1219),
.Y(n_1701)
);

AO31x2_ASAP7_75t_L g1702 ( 
.A1(n_1297),
.A2(n_1257),
.A3(n_1169),
.B(n_1254),
.Y(n_1702)
);

AO31x2_ASAP7_75t_L g1703 ( 
.A1(n_1297),
.A2(n_1257),
.A3(n_1169),
.B(n_1254),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1218),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1218),
.Y(n_1705)
);

AO31x2_ASAP7_75t_L g1706 ( 
.A1(n_1297),
.A2(n_1257),
.A3(n_1169),
.B(n_1254),
.Y(n_1706)
);

AO31x2_ASAP7_75t_L g1707 ( 
.A1(n_1297),
.A2(n_1257),
.A3(n_1169),
.B(n_1254),
.Y(n_1707)
);

AO31x2_ASAP7_75t_L g1708 ( 
.A1(n_1297),
.A2(n_1257),
.A3(n_1169),
.B(n_1254),
.Y(n_1708)
);

OAI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1254),
.A2(n_1352),
.B(n_1337),
.Y(n_1709)
);

AO31x2_ASAP7_75t_L g1710 ( 
.A1(n_1297),
.A2(n_1257),
.A3(n_1169),
.B(n_1254),
.Y(n_1710)
);

NAND2x1p5_ASAP7_75t_L g1711 ( 
.A(n_1219),
.B(n_1332),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1404),
.B(n_1014),
.Y(n_1712)
);

INVx2_ASAP7_75t_SL g1713 ( 
.A(n_1332),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1218),
.Y(n_1714)
);

AO32x2_ASAP7_75t_L g1715 ( 
.A1(n_1290),
.A2(n_1300),
.A3(n_1293),
.B1(n_1361),
.B2(n_1341),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1218),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1414),
.B(n_1014),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1330),
.B(n_1218),
.Y(n_1718)
);

OR2x6_ASAP7_75t_L g1719 ( 
.A(n_1533),
.B(n_1701),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1621),
.B(n_1648),
.Y(n_1720)
);

AOI21xp33_ASAP7_75t_L g1721 ( 
.A1(n_1547),
.A2(n_1679),
.B(n_1638),
.Y(n_1721)
);

INVxp67_ASAP7_75t_SL g1722 ( 
.A(n_1482),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1618),
.Y(n_1723)
);

INVx4_ASAP7_75t_L g1724 ( 
.A(n_1636),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1557),
.B(n_1712),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1660),
.Y(n_1726)
);

NAND2xp33_ASAP7_75t_L g1727 ( 
.A(n_1604),
.B(n_1549),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1685),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1700),
.Y(n_1729)
);

OAI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1568),
.A2(n_1622),
.B(n_1560),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1592),
.B(n_1562),
.Y(n_1731)
);

NAND2x1p5_ASAP7_75t_L g1732 ( 
.A(n_1701),
.B(n_1636),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1565),
.A2(n_1546),
.B(n_1651),
.Y(n_1733)
);

A2O1A1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1683),
.A2(n_1688),
.B(n_1585),
.C(n_1577),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1619),
.B(n_1650),
.Y(n_1735)
);

OA21x2_ASAP7_75t_L g1736 ( 
.A1(n_1684),
.A2(n_1709),
.B(n_1691),
.Y(n_1736)
);

OAI21x1_ASAP7_75t_SL g1737 ( 
.A1(n_1605),
.A2(n_1697),
.B(n_1677),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1467),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1569),
.A2(n_1691),
.B(n_1684),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1634),
.A2(n_1576),
.B1(n_1461),
.B2(n_1588),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1617),
.B(n_1632),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1476),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1620),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1631),
.Y(n_1744)
);

AOI21x1_ASAP7_75t_L g1745 ( 
.A1(n_1597),
.A2(n_1591),
.B(n_1633),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1717),
.B(n_1674),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1669),
.B(n_1572),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1693),
.B(n_1491),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1593),
.A2(n_1483),
.B1(n_1492),
.B2(n_1497),
.Y(n_1749)
);

AND2x4_ASAP7_75t_SL g1750 ( 
.A(n_1478),
.B(n_1447),
.Y(n_1750)
);

AO21x2_ASAP7_75t_L g1751 ( 
.A1(n_1555),
.A2(n_1639),
.B(n_1612),
.Y(n_1751)
);

BUFx3_ASAP7_75t_L g1752 ( 
.A(n_1637),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1636),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1687),
.B(n_1500),
.Y(n_1754)
);

AOI21xp33_ASAP7_75t_SL g1755 ( 
.A1(n_1615),
.A2(n_1681),
.B(n_1471),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1645),
.Y(n_1756)
);

AO21x2_ASAP7_75t_L g1757 ( 
.A1(n_1555),
.A2(n_1639),
.B(n_1612),
.Y(n_1757)
);

AND2x6_ASAP7_75t_L g1758 ( 
.A(n_1504),
.B(n_1558),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1655),
.Y(n_1759)
);

BUFx3_ASAP7_75t_L g1760 ( 
.A(n_1662),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1616),
.B(n_1642),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1491),
.B(n_1457),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1665),
.B(n_1673),
.Y(n_1763)
);

BUFx2_ASAP7_75t_R g1764 ( 
.A(n_1614),
.Y(n_1764)
);

NAND2x1p5_ASAP7_75t_L g1765 ( 
.A(n_1662),
.B(n_1459),
.Y(n_1765)
);

OAI211xp5_ASAP7_75t_SL g1766 ( 
.A1(n_1452),
.A2(n_1538),
.B(n_1453),
.C(n_1446),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1533),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1676),
.B(n_1692),
.Y(n_1768)
);

OR2x6_ASAP7_75t_L g1769 ( 
.A(n_1533),
.B(n_1549),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1447),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1696),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1704),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1705),
.Y(n_1773)
);

BUFx2_ASAP7_75t_L g1774 ( 
.A(n_1459),
.Y(n_1774)
);

AO31x2_ASAP7_75t_L g1775 ( 
.A1(n_1543),
.A2(n_1598),
.A3(n_1552),
.B(n_1599),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1662),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1714),
.Y(n_1777)
);

INVxp67_ASAP7_75t_L g1778 ( 
.A(n_1506),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1504),
.A2(n_1451),
.B1(n_1629),
.B2(n_1458),
.Y(n_1779)
);

OAI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1654),
.A2(n_1659),
.B(n_1657),
.Y(n_1780)
);

BUFx2_ASAP7_75t_R g1781 ( 
.A(n_1541),
.Y(n_1781)
);

AND2x6_ASAP7_75t_SL g1782 ( 
.A(n_1526),
.B(n_1544),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1634),
.A2(n_1580),
.B1(n_1545),
.B2(n_1561),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1716),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1494),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1450),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1528),
.Y(n_1787)
);

OAI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1670),
.A2(n_1682),
.B(n_1672),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1528),
.Y(n_1789)
);

OR2x6_ASAP7_75t_L g1790 ( 
.A(n_1549),
.B(n_1667),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1640),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1510),
.B(n_1671),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1671),
.B(n_1567),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1519),
.Y(n_1794)
);

BUFx3_ASAP7_75t_L g1795 ( 
.A(n_1600),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1519),
.Y(n_1796)
);

OAI221xp5_ASAP7_75t_L g1797 ( 
.A1(n_1570),
.A2(n_1469),
.B1(n_1584),
.B2(n_1554),
.C(n_1596),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1603),
.B(n_1536),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1457),
.B(n_1689),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1493),
.Y(n_1800)
);

INVx3_ASAP7_75t_L g1801 ( 
.A(n_1640),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1523),
.Y(n_1802)
);

OAI21xp33_ASAP7_75t_L g1803 ( 
.A1(n_1536),
.A2(n_1477),
.B(n_1575),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1698),
.B(n_1478),
.Y(n_1804)
);

AOI21x1_ASAP7_75t_L g1805 ( 
.A1(n_1595),
.A2(n_1608),
.B(n_1564),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1506),
.B(n_1473),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1523),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1658),
.B(n_1582),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1581),
.A2(n_1582),
.B1(n_1596),
.B2(n_1550),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1649),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1623),
.B(n_1689),
.Y(n_1811)
);

BUFx8_ASAP7_75t_L g1812 ( 
.A(n_1466),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1501),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1507),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1558),
.Y(n_1815)
);

OR2x6_ASAP7_75t_L g1816 ( 
.A(n_1667),
.B(n_1694),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1512),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1578),
.A2(n_1548),
.B(n_1609),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1694),
.B(n_1711),
.Y(n_1819)
);

OAI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1594),
.A2(n_1509),
.B(n_1609),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1520),
.A2(n_1530),
.B1(n_1556),
.B2(n_1539),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1513),
.Y(n_1822)
);

BUFx2_ASAP7_75t_R g1823 ( 
.A(n_1553),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1548),
.A2(n_1626),
.B(n_1610),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1624),
.B(n_1627),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1515),
.Y(n_1826)
);

OAI222xp33_ASAP7_75t_SL g1827 ( 
.A1(n_1526),
.A2(n_1643),
.B1(n_1511),
.B2(n_1484),
.C1(n_1462),
.C2(n_1656),
.Y(n_1827)
);

A2O1A1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1479),
.A2(n_1535),
.B(n_1534),
.C(n_1529),
.Y(n_1828)
);

OA21x2_ASAP7_75t_L g1829 ( 
.A1(n_1479),
.A2(n_1474),
.B(n_1496),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1603),
.B(n_1628),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1624),
.B(n_1627),
.Y(n_1831)
);

OAI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1509),
.A2(n_1610),
.B(n_1626),
.Y(n_1832)
);

OA21x2_ASAP7_75t_L g1833 ( 
.A1(n_1489),
.A2(n_1534),
.B(n_1529),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1647),
.B(n_1652),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1586),
.A2(n_1454),
.B(n_1690),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1514),
.Y(n_1836)
);

AO21x2_ASAP7_75t_L g1837 ( 
.A1(n_1516),
.A2(n_1595),
.B(n_1601),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1514),
.Y(n_1838)
);

AO31x2_ASAP7_75t_L g1839 ( 
.A1(n_1574),
.A2(n_1661),
.A3(n_1690),
.B(n_1675),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1571),
.B(n_1537),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1647),
.A2(n_1718),
.B(n_1664),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1521),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1686),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1711),
.B(n_1448),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1521),
.A2(n_1524),
.B1(n_1527),
.B2(n_1663),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1661),
.B(n_1663),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1628),
.B(n_1607),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1713),
.B(n_1630),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1664),
.B(n_1579),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1641),
.B(n_1680),
.Y(n_1850)
);

AO21x2_ASAP7_75t_L g1851 ( 
.A1(n_1646),
.A2(n_1518),
.B(n_1517),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1563),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1607),
.B(n_1606),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1525),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1531),
.B(n_1532),
.Y(n_1855)
);

INVx4_ASAP7_75t_L g1856 ( 
.A(n_1470),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1531),
.B(n_1532),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1573),
.A2(n_1589),
.B(n_1518),
.Y(n_1858)
);

OAI21x1_ASAP7_75t_SL g1859 ( 
.A1(n_1463),
.A2(n_1495),
.B(n_1499),
.Y(n_1859)
);

BUFx8_ASAP7_75t_SL g1860 ( 
.A(n_1695),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1525),
.Y(n_1861)
);

BUFx2_ASAP7_75t_L g1862 ( 
.A(n_1508),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1625),
.B(n_1587),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1475),
.B(n_1485),
.Y(n_1864)
);

INVx3_ASAP7_75t_L g1865 ( 
.A(n_1508),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1715),
.B(n_1571),
.Y(n_1866)
);

NOR2xp67_ASAP7_75t_L g1867 ( 
.A(n_1668),
.B(n_1481),
.Y(n_1867)
);

OA21x2_ASAP7_75t_L g1868 ( 
.A1(n_1468),
.A2(n_1524),
.B(n_1472),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1566),
.Y(n_1869)
);

A2O1A1Ixp33_ASAP7_75t_L g1870 ( 
.A1(n_1503),
.A2(n_1505),
.B(n_1502),
.C(n_1464),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1715),
.B(n_1465),
.Y(n_1871)
);

BUFx2_ASAP7_75t_L g1872 ( 
.A(n_1542),
.Y(n_1872)
);

NAND3xp33_ASAP7_75t_L g1873 ( 
.A(n_1480),
.B(n_1487),
.C(n_1498),
.Y(n_1873)
);

O2A1O1Ixp33_ASAP7_75t_L g1874 ( 
.A1(n_1583),
.A2(n_1590),
.B(n_1456),
.C(n_1455),
.Y(n_1874)
);

AO31x2_ASAP7_75t_L g1875 ( 
.A1(n_1486),
.A2(n_1635),
.A3(n_1710),
.B(n_1708),
.Y(n_1875)
);

OA21x2_ASAP7_75t_L g1876 ( 
.A1(n_1602),
.A2(n_1486),
.B(n_1490),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1559),
.Y(n_1877)
);

BUFx2_ASAP7_75t_L g1878 ( 
.A(n_1715),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1559),
.A2(n_1465),
.B1(n_1602),
.B2(n_1710),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1613),
.B(n_1653),
.Y(n_1880)
);

BUFx3_ASAP7_75t_L g1881 ( 
.A(n_1540),
.Y(n_1881)
);

A2O1A1Ixp33_ASAP7_75t_L g1882 ( 
.A1(n_1460),
.A2(n_1540),
.B(n_1488),
.C(n_1653),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1635),
.B(n_1699),
.Y(n_1883)
);

OA21x2_ASAP7_75t_L g1884 ( 
.A1(n_1635),
.A2(n_1699),
.B(n_1707),
.Y(n_1884)
);

AO31x2_ASAP7_75t_L g1885 ( 
.A1(n_1644),
.A2(n_1702),
.A3(n_1707),
.B(n_1706),
.Y(n_1885)
);

AO31x2_ASAP7_75t_L g1886 ( 
.A1(n_1644),
.A2(n_1666),
.A3(n_1706),
.B(n_1703),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1653),
.B(n_1702),
.Y(n_1887)
);

AOI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1551),
.A2(n_1702),
.B1(n_1703),
.B2(n_1706),
.Y(n_1888)
);

OR2x6_ASAP7_75t_L g1889 ( 
.A(n_1522),
.B(n_1460),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1703),
.B(n_1708),
.Y(n_1890)
);

OAI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1568),
.A2(n_1410),
.B(n_1622),
.Y(n_1891)
);

OR2x6_ASAP7_75t_L g1892 ( 
.A(n_1533),
.B(n_1262),
.Y(n_1892)
);

CKINVDCx6p67_ASAP7_75t_R g1893 ( 
.A(n_1637),
.Y(n_1893)
);

BUFx3_ASAP7_75t_L g1894 ( 
.A(n_1637),
.Y(n_1894)
);

BUFx2_ASAP7_75t_L g1895 ( 
.A(n_1637),
.Y(n_1895)
);

NAND2x1p5_ASAP7_75t_L g1896 ( 
.A(n_1701),
.B(n_1219),
.Y(n_1896)
);

INVxp67_ASAP7_75t_L g1897 ( 
.A(n_1533),
.Y(n_1897)
);

OR2x6_ASAP7_75t_L g1898 ( 
.A(n_1533),
.B(n_1262),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1557),
.B(n_1014),
.Y(n_1899)
);

NOR2x1_ASAP7_75t_SL g1900 ( 
.A(n_1533),
.B(n_1262),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1449),
.Y(n_1901)
);

AOI21x1_ASAP7_75t_L g1902 ( 
.A1(n_1597),
.A2(n_1678),
.B(n_1611),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1449),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1621),
.B(n_1648),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1449),
.Y(n_1905)
);

AO21x2_ASAP7_75t_L g1906 ( 
.A1(n_1737),
.A2(n_1882),
.B(n_1733),
.Y(n_1906)
);

BUFx2_ASAP7_75t_L g1907 ( 
.A(n_1758),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1860),
.Y(n_1908)
);

HB1xp67_ASAP7_75t_L g1909 ( 
.A(n_1762),
.Y(n_1909)
);

OR2x6_ASAP7_75t_L g1910 ( 
.A(n_1892),
.B(n_1898),
.Y(n_1910)
);

BUFx3_ASAP7_75t_L g1911 ( 
.A(n_1732),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1877),
.Y(n_1912)
);

OAI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1870),
.A2(n_1721),
.B(n_1797),
.Y(n_1913)
);

AO21x2_ASAP7_75t_L g1914 ( 
.A1(n_1902),
.A2(n_1788),
.B(n_1780),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1899),
.B(n_1731),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1854),
.Y(n_1916)
);

AOI21x1_ASAP7_75t_L g1917 ( 
.A1(n_1745),
.A2(n_1824),
.B(n_1818),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1861),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1766),
.B(n_1741),
.Y(n_1919)
);

BUFx2_ASAP7_75t_L g1920 ( 
.A(n_1758),
.Y(n_1920)
);

AO21x2_ASAP7_75t_L g1921 ( 
.A1(n_1739),
.A2(n_1820),
.B(n_1832),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1725),
.B(n_1720),
.Y(n_1922)
);

INVx8_ASAP7_75t_L g1923 ( 
.A(n_1758),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1901),
.B(n_1903),
.Y(n_1924)
);

OR2x6_ASAP7_75t_L g1925 ( 
.A(n_1892),
.B(n_1898),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1799),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1901),
.B(n_1903),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1904),
.B(n_1849),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1897),
.B(n_1746),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1839),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_L g1931 ( 
.A(n_1897),
.B(n_1892),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1905),
.B(n_1826),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1905),
.B(n_1826),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1839),
.Y(n_1934)
);

OR2x6_ASAP7_75t_L g1935 ( 
.A(n_1898),
.B(n_1769),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1839),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1786),
.B(n_1800),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1839),
.Y(n_1938)
);

NOR3xp33_ASAP7_75t_L g1939 ( 
.A(n_1808),
.B(n_1779),
.C(n_1754),
.Y(n_1939)
);

BUFx3_ASAP7_75t_L g1940 ( 
.A(n_1732),
.Y(n_1940)
);

AOI222xp33_ASAP7_75t_L g1941 ( 
.A1(n_1783),
.A2(n_1747),
.B1(n_1900),
.B2(n_1735),
.C1(n_1740),
.C2(n_1754),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1786),
.B(n_1800),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1817),
.B(n_1852),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1817),
.B(n_1852),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1783),
.B(n_1821),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1878),
.B(n_1866),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_SL g1947 ( 
.A1(n_1798),
.A2(n_1828),
.B(n_1830),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1825),
.B(n_1831),
.Y(n_1948)
);

NOR2x1_ASAP7_75t_R g1949 ( 
.A(n_1728),
.B(n_1843),
.Y(n_1949)
);

BUFx2_ASAP7_75t_L g1950 ( 
.A(n_1758),
.Y(n_1950)
);

INVxp67_ASAP7_75t_SL g1951 ( 
.A(n_1722),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1767),
.B(n_1872),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1834),
.B(n_1846),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1821),
.B(n_1723),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1738),
.B(n_1742),
.Y(n_1955)
);

CKINVDCx20_ASAP7_75t_R g1956 ( 
.A(n_1860),
.Y(n_1956)
);

NAND2x1_ASAP7_75t_L g1957 ( 
.A(n_1829),
.B(n_1889),
.Y(n_1957)
);

OR2x6_ASAP7_75t_L g1958 ( 
.A(n_1769),
.B(n_1719),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1836),
.B(n_1838),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1726),
.B(n_1729),
.Y(n_1960)
);

OR2x6_ASAP7_75t_L g1961 ( 
.A(n_1769),
.B(n_1719),
.Y(n_1961)
);

OR2x6_ASAP7_75t_L g1962 ( 
.A(n_1719),
.B(n_1798),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1736),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1743),
.Y(n_1964)
);

BUFx3_ASAP7_75t_L g1965 ( 
.A(n_1761),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1815),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1815),
.Y(n_1967)
);

INVx3_ASAP7_75t_L g1968 ( 
.A(n_1724),
.Y(n_1968)
);

INVx3_ASAP7_75t_L g1969 ( 
.A(n_1724),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1744),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1756),
.Y(n_1971)
);

HB1xp67_ASAP7_75t_L g1972 ( 
.A(n_1760),
.Y(n_1972)
);

INVx3_ASAP7_75t_L g1973 ( 
.A(n_1856),
.Y(n_1973)
);

INVx4_ASAP7_75t_SL g1974 ( 
.A(n_1790),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_1782),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1759),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1842),
.B(n_1748),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1771),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1772),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1773),
.Y(n_1980)
);

AO21x2_ASAP7_75t_L g1981 ( 
.A1(n_1891),
.A2(n_1730),
.B(n_1835),
.Y(n_1981)
);

BUFx3_ASAP7_75t_L g1982 ( 
.A(n_1760),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1777),
.Y(n_1983)
);

NOR2xp33_ASAP7_75t_L g1984 ( 
.A(n_1778),
.B(n_1863),
.Y(n_1984)
);

INVx2_ASAP7_75t_SL g1985 ( 
.A(n_1765),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1784),
.B(n_1763),
.Y(n_1986)
);

BUFx12f_ASAP7_75t_L g1987 ( 
.A(n_1812),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1809),
.B(n_1787),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1785),
.Y(n_1989)
);

OR2x2_ASAP7_75t_L g1990 ( 
.A(n_1722),
.B(n_1806),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1789),
.Y(n_1991)
);

CKINVDCx20_ASAP7_75t_R g1992 ( 
.A(n_1893),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1794),
.B(n_1796),
.Y(n_1993)
);

HB1xp67_ASAP7_75t_L g1994 ( 
.A(n_1752),
.Y(n_1994)
);

AOI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1740),
.A2(n_1845),
.B1(n_1749),
.B2(n_1792),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1802),
.B(n_1807),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1871),
.B(n_1813),
.Y(n_1997)
);

HB1xp67_ASAP7_75t_L g1998 ( 
.A(n_1752),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1890),
.B(n_1875),
.Y(n_1999)
);

AO21x1_ASAP7_75t_SL g2000 ( 
.A1(n_1803),
.A2(n_1845),
.B(n_1810),
.Y(n_2000)
);

OA21x2_ASAP7_75t_L g2001 ( 
.A1(n_1880),
.A2(n_1887),
.B(n_1883),
.Y(n_2001)
);

INVx3_ASAP7_75t_L g2002 ( 
.A(n_1765),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1894),
.Y(n_2003)
);

AO21x2_ASAP7_75t_L g2004 ( 
.A1(n_1734),
.A2(n_1888),
.B(n_1805),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1894),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1814),
.B(n_1822),
.Y(n_2006)
);

INVx3_ASAP7_75t_L g2007 ( 
.A(n_1790),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_1812),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1997),
.B(n_1837),
.Y(n_2009)
);

INVx1_ASAP7_75t_SL g2010 ( 
.A(n_2008),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1916),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1997),
.B(n_1837),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1932),
.B(n_1884),
.Y(n_2013)
);

AO21x2_ASAP7_75t_L g2014 ( 
.A1(n_1917),
.A2(n_1913),
.B(n_1914),
.Y(n_2014)
);

INVxp67_ASAP7_75t_SL g2015 ( 
.A(n_1951),
.Y(n_2015)
);

AND2x2_ASAP7_75t_SL g2016 ( 
.A(n_1907),
.B(n_1727),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1916),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1918),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1918),
.Y(n_2019)
);

OAI21xp5_ASAP7_75t_SL g2020 ( 
.A1(n_1941),
.A2(n_1778),
.B(n_1896),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1932),
.B(n_1933),
.Y(n_2021)
);

HB1xp67_ASAP7_75t_L g2022 ( 
.A(n_1966),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1933),
.B(n_1884),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1948),
.B(n_1768),
.Y(n_2024)
);

AOI22xp33_ASAP7_75t_L g2025 ( 
.A1(n_1939),
.A2(n_1851),
.B1(n_1859),
.B2(n_1855),
.Y(n_2025)
);

NOR2xp33_ASAP7_75t_L g2026 ( 
.A(n_1922),
.B(n_1755),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1948),
.B(n_1857),
.Y(n_2027)
);

BUFx3_ASAP7_75t_L g2028 ( 
.A(n_1982),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1953),
.B(n_1793),
.Y(n_2029)
);

AOI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_1945),
.A2(n_1851),
.B1(n_1811),
.B2(n_1833),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1953),
.B(n_1811),
.Y(n_2031)
);

NOR2x1_ASAP7_75t_SL g2032 ( 
.A(n_1958),
.B(n_1847),
.Y(n_2032)
);

OR2x2_ASAP7_75t_L g2033 ( 
.A(n_1946),
.B(n_1885),
.Y(n_2033)
);

INVxp67_ASAP7_75t_SL g2034 ( 
.A(n_1967),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1963),
.Y(n_2035)
);

INVx2_ASAP7_75t_SL g2036 ( 
.A(n_1911),
.Y(n_2036)
);

INVx3_ASAP7_75t_L g2037 ( 
.A(n_1957),
.Y(n_2037)
);

HB1xp67_ASAP7_75t_L g2038 ( 
.A(n_1972),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1924),
.B(n_1876),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1924),
.B(n_1876),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1927),
.B(n_1885),
.Y(n_2041)
);

OR2x2_ASAP7_75t_L g2042 ( 
.A(n_1977),
.B(n_1885),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1937),
.B(n_1886),
.Y(n_2043)
);

INVxp67_ASAP7_75t_SL g2044 ( 
.A(n_1990),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1993),
.B(n_1841),
.Y(n_2045)
);

OR2x6_ASAP7_75t_L g2046 ( 
.A(n_1923),
.B(n_1830),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1937),
.B(n_1886),
.Y(n_2047)
);

HB1xp67_ASAP7_75t_L g2048 ( 
.A(n_1982),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1993),
.B(n_1858),
.Y(n_2049)
);

INVxp67_ASAP7_75t_SL g2050 ( 
.A(n_1990),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1942),
.B(n_1886),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1996),
.B(n_1869),
.Y(n_2052)
);

HB1xp67_ASAP7_75t_L g2053 ( 
.A(n_1982),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1943),
.B(n_1775),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1943),
.B(n_1775),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_1959),
.B(n_1879),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1944),
.B(n_1775),
.Y(n_2057)
);

INVx5_ASAP7_75t_L g2058 ( 
.A(n_1923),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1944),
.B(n_1988),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1996),
.B(n_1928),
.Y(n_2060)
);

BUFx3_ASAP7_75t_L g2061 ( 
.A(n_1911),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1915),
.B(n_2006),
.Y(n_2062)
);

HB1xp67_ASAP7_75t_L g2063 ( 
.A(n_1909),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1988),
.B(n_1775),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1999),
.B(n_1921),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1999),
.B(n_1921),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_2006),
.B(n_1869),
.Y(n_2067)
);

INVx3_ASAP7_75t_SL g2068 ( 
.A(n_2008),
.Y(n_2068)
);

INVx5_ASAP7_75t_SL g2069 ( 
.A(n_1958),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1921),
.B(n_1881),
.Y(n_2070)
);

AOI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_1919),
.A2(n_1833),
.B1(n_1840),
.B2(n_1868),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1960),
.B(n_1840),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1954),
.B(n_1959),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1954),
.B(n_1751),
.Y(n_2074)
);

HB1xp67_ASAP7_75t_L g2075 ( 
.A(n_1926),
.Y(n_2075)
);

INVx1_ASAP7_75t_SL g2076 ( 
.A(n_1994),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1960),
.B(n_1757),
.Y(n_2077)
);

HB1xp67_ASAP7_75t_L g2078 ( 
.A(n_1998),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2011),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_2033),
.B(n_1912),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2011),
.Y(n_2081)
);

OR2x2_ASAP7_75t_L g2082 ( 
.A(n_2033),
.B(n_1912),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2059),
.B(n_1930),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_2059),
.B(n_1934),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2021),
.B(n_1964),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2017),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_L g2087 ( 
.A(n_2010),
.B(n_1764),
.Y(n_2087)
);

INVxp67_ASAP7_75t_L g2088 ( 
.A(n_2078),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_2064),
.B(n_1934),
.Y(n_2089)
);

HB1xp67_ASAP7_75t_L g2090 ( 
.A(n_2038),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2017),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2018),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2018),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2019),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2064),
.B(n_1936),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2019),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2065),
.B(n_1936),
.Y(n_2097)
);

AND2x4_ASAP7_75t_SL g2098 ( 
.A(n_2046),
.B(n_1958),
.Y(n_2098)
);

AND2x4_ASAP7_75t_L g2099 ( 
.A(n_2013),
.B(n_2023),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2065),
.B(n_1938),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2066),
.B(n_1938),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2066),
.B(n_2054),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_2054),
.B(n_2004),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2055),
.B(n_2004),
.Y(n_2104)
);

INVx1_ASAP7_75t_SL g2105 ( 
.A(n_2068),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2055),
.B(n_2004),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2057),
.B(n_2001),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_2035),
.Y(n_2108)
);

INVxp67_ASAP7_75t_L g2109 ( 
.A(n_2076),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2021),
.B(n_1964),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2057),
.B(n_2001),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2077),
.B(n_2001),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2031),
.B(n_1970),
.Y(n_2113)
);

INVx3_ASAP7_75t_L g2114 ( 
.A(n_2037),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2077),
.B(n_2001),
.Y(n_2115)
);

INVx4_ASAP7_75t_L g2116 ( 
.A(n_2058),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2073),
.B(n_1981),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2073),
.B(n_1981),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2074),
.B(n_1981),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2062),
.B(n_1970),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2060),
.B(n_1971),
.Y(n_2121)
);

BUFx2_ASAP7_75t_L g2122 ( 
.A(n_2015),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2041),
.B(n_2043),
.Y(n_2123)
);

INVx2_ASAP7_75t_SL g2124 ( 
.A(n_2028),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2044),
.B(n_1971),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2043),
.B(n_1906),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2047),
.B(n_1906),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2050),
.B(n_1976),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2047),
.B(n_1906),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2063),
.B(n_1976),
.Y(n_2130)
);

INVx2_ASAP7_75t_SL g2131 ( 
.A(n_2028),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2079),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2099),
.B(n_2009),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2099),
.B(n_2009),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2099),
.B(n_2012),
.Y(n_2135)
);

NOR2xp67_ASAP7_75t_L g2136 ( 
.A(n_2116),
.B(n_2058),
.Y(n_2136)
);

OR2x2_ASAP7_75t_L g2137 ( 
.A(n_2102),
.B(n_2042),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2079),
.Y(n_2138)
);

AND2x4_ASAP7_75t_L g2139 ( 
.A(n_2114),
.B(n_2037),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2099),
.B(n_2012),
.Y(n_2140)
);

INVx1_ASAP7_75t_SL g2141 ( 
.A(n_2105),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_2083),
.B(n_2075),
.Y(n_2142)
);

OR2x2_ASAP7_75t_L g2143 ( 
.A(n_2102),
.B(n_2056),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2108),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2122),
.B(n_2056),
.Y(n_2145)
);

INVx2_ASAP7_75t_SL g2146 ( 
.A(n_2122),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2081),
.Y(n_2147)
);

INVx1_ASAP7_75t_SL g2148 ( 
.A(n_2090),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2083),
.B(n_2022),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2123),
.B(n_2070),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2081),
.Y(n_2151)
);

OR2x2_ASAP7_75t_L g2152 ( 
.A(n_2123),
.B(n_2051),
.Y(n_2152)
);

NAND2xp33_ASAP7_75t_R g2153 ( 
.A(n_2087),
.B(n_1975),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2117),
.B(n_2070),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2084),
.B(n_2034),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2086),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2086),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2117),
.B(n_2039),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2118),
.B(n_2039),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2084),
.B(n_2045),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2091),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2091),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2113),
.B(n_2085),
.Y(n_2163)
);

INVx1_ASAP7_75t_SL g2164 ( 
.A(n_2124),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2092),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2110),
.B(n_2071),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2120),
.B(n_2071),
.Y(n_2167)
);

NOR3xp33_ASAP7_75t_L g2168 ( 
.A(n_2109),
.B(n_2020),
.C(n_2026),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2118),
.B(n_2040),
.Y(n_2169)
);

NAND2x1_ASAP7_75t_L g2170 ( 
.A(n_2116),
.B(n_1910),
.Y(n_2170)
);

NOR2x1_ASAP7_75t_SL g2171 ( 
.A(n_2116),
.B(n_1935),
.Y(n_2171)
);

NOR2xp33_ASAP7_75t_L g2172 ( 
.A(n_2088),
.B(n_1975),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2132),
.Y(n_2173)
);

OAI22xp5_ASAP7_75t_L g2174 ( 
.A1(n_2136),
.A2(n_1910),
.B1(n_1925),
.B2(n_2116),
.Y(n_2174)
);

AOI22xp5_ASAP7_75t_L g2175 ( 
.A1(n_2168),
.A2(n_2020),
.B1(n_1925),
.B2(n_1910),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2158),
.B(n_2159),
.Y(n_2176)
);

INVx1_ASAP7_75t_SL g2177 ( 
.A(n_2141),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2144),
.Y(n_2178)
);

OR2x2_ASAP7_75t_L g2179 ( 
.A(n_2137),
.B(n_2112),
.Y(n_2179)
);

OAI221xp5_ASAP7_75t_SL g2180 ( 
.A1(n_2143),
.A2(n_1995),
.B1(n_1910),
.B2(n_1925),
.C(n_1935),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2132),
.Y(n_2181)
);

BUFx2_ASAP7_75t_L g2182 ( 
.A(n_2146),
.Y(n_2182)
);

NAND2x1_ASAP7_75t_SL g2183 ( 
.A(n_2136),
.B(n_2114),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2167),
.B(n_2097),
.Y(n_2184)
);

AOI222xp33_ASAP7_75t_L g2185 ( 
.A1(n_2166),
.A2(n_1929),
.B1(n_2130),
.B2(n_2067),
.C1(n_2052),
.C2(n_2121),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2154),
.B(n_2097),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2138),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2144),
.Y(n_2188)
);

OAI22xp33_ASAP7_75t_SL g2189 ( 
.A1(n_2170),
.A2(n_1925),
.B1(n_1910),
.B2(n_1935),
.Y(n_2189)
);

OR2x2_ASAP7_75t_L g2190 ( 
.A(n_2137),
.B(n_2112),
.Y(n_2190)
);

AND2x4_ASAP7_75t_L g2191 ( 
.A(n_2171),
.B(n_2114),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2158),
.B(n_2159),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2154),
.B(n_2100),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2160),
.B(n_2100),
.Y(n_2194)
);

AOI21xp33_ASAP7_75t_SL g2195 ( 
.A1(n_2153),
.A2(n_2068),
.B(n_1908),
.Y(n_2195)
);

OAI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_2170),
.A2(n_1925),
.B1(n_1935),
.B2(n_1958),
.Y(n_2196)
);

OR2x2_ASAP7_75t_L g2197 ( 
.A(n_2152),
.B(n_2115),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2138),
.Y(n_2198)
);

OR2x2_ASAP7_75t_L g2199 ( 
.A(n_2152),
.B(n_2115),
.Y(n_2199)
);

OAI21xp5_ASAP7_75t_L g2200 ( 
.A1(n_2146),
.A2(n_2005),
.B(n_2003),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_2144),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2169),
.B(n_2101),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2169),
.B(n_2101),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2147),
.Y(n_2204)
);

INVx1_ASAP7_75t_SL g2205 ( 
.A(n_2148),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2147),
.Y(n_2206)
);

O2A1O1Ixp33_ASAP7_75t_L g2207 ( 
.A1(n_2195),
.A2(n_2172),
.B(n_2068),
.C(n_1952),
.Y(n_2207)
);

AOI211xp5_ASAP7_75t_SL g2208 ( 
.A1(n_2189),
.A2(n_2171),
.B(n_2145),
.C(n_1947),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_2176),
.B(n_2133),
.Y(n_2209)
);

NAND2xp33_ASAP7_75t_L g2210 ( 
.A(n_2174),
.B(n_1923),
.Y(n_2210)
);

NOR3xp33_ASAP7_75t_L g2211 ( 
.A(n_2180),
.B(n_1949),
.C(n_1865),
.Y(n_2211)
);

OR2x2_ASAP7_75t_L g2212 ( 
.A(n_2179),
.B(n_2143),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2176),
.B(n_2150),
.Y(n_2213)
);

AOI321xp33_ASAP7_75t_L g2214 ( 
.A1(n_2175),
.A2(n_2149),
.A3(n_2142),
.B1(n_2155),
.B2(n_2163),
.C(n_2145),
.Y(n_2214)
);

AOI32xp33_ASAP7_75t_L g2215 ( 
.A1(n_2182),
.A2(n_2150),
.A3(n_2135),
.B1(n_2140),
.B2(n_2134),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2173),
.Y(n_2216)
);

INVx1_ASAP7_75t_SL g2217 ( 
.A(n_2177),
.Y(n_2217)
);

AOI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_2185),
.A2(n_2133),
.B1(n_2135),
.B2(n_2134),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2181),
.Y(n_2219)
);

NOR2xp67_ASAP7_75t_L g2220 ( 
.A(n_2191),
.B(n_1987),
.Y(n_2220)
);

AOI322xp5_ASAP7_75t_L g2221 ( 
.A1(n_2192),
.A2(n_2205),
.A3(n_2203),
.B1(n_2202),
.B2(n_2186),
.C1(n_2193),
.C2(n_2184),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2192),
.B(n_2182),
.Y(n_2222)
);

AOI31xp33_ASAP7_75t_L g2223 ( 
.A1(n_2196),
.A2(n_1949),
.A3(n_1908),
.B(n_1728),
.Y(n_2223)
);

OAI21xp33_ASAP7_75t_L g2224 ( 
.A1(n_2197),
.A2(n_2140),
.B(n_2164),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2187),
.Y(n_2225)
);

XNOR2x1_ASAP7_75t_L g2226 ( 
.A(n_2197),
.B(n_1935),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2198),
.Y(n_2227)
);

AOI221xp5_ASAP7_75t_SL g2228 ( 
.A1(n_2194),
.A2(n_1956),
.B1(n_1931),
.B2(n_2072),
.C(n_1992),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2204),
.Y(n_2229)
);

AOI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_2191),
.A2(n_2119),
.B1(n_2089),
.B2(n_2095),
.Y(n_2230)
);

OAI21xp5_ASAP7_75t_SL g2231 ( 
.A1(n_2191),
.A2(n_2098),
.B(n_2025),
.Y(n_2231)
);

OAI321xp33_ASAP7_75t_L g2232 ( 
.A1(n_2200),
.A2(n_1961),
.A3(n_2124),
.B1(n_2131),
.B2(n_2030),
.C(n_1962),
.Y(n_2232)
);

HB1xp67_ASAP7_75t_L g2233 ( 
.A(n_2178),
.Y(n_2233)
);

AND2x4_ASAP7_75t_L g2234 ( 
.A(n_2199),
.B(n_2139),
.Y(n_2234)
);

NOR2x1_ASAP7_75t_L g2235 ( 
.A(n_2199),
.B(n_1961),
.Y(n_2235)
);

OAI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_2179),
.A2(n_1961),
.B1(n_2098),
.B2(n_2016),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_SL g2237 ( 
.A(n_2178),
.B(n_2139),
.Y(n_2237)
);

INVx1_ASAP7_75t_SL g2238 ( 
.A(n_2190),
.Y(n_2238)
);

OAI22xp5_ASAP7_75t_L g2239 ( 
.A1(n_2220),
.A2(n_2190),
.B1(n_2098),
.B2(n_2016),
.Y(n_2239)
);

OAI21xp5_ASAP7_75t_SL g2240 ( 
.A1(n_2208),
.A2(n_1827),
.B(n_1987),
.Y(n_2240)
);

O2A1O1Ixp33_ASAP7_75t_L g2241 ( 
.A1(n_2223),
.A2(n_1961),
.B(n_2027),
.C(n_1865),
.Y(n_2241)
);

AOI22xp33_ASAP7_75t_SL g2242 ( 
.A1(n_2210),
.A2(n_2032),
.B1(n_2016),
.B2(n_2069),
.Y(n_2242)
);

O2A1O1Ixp33_ASAP7_75t_L g2243 ( 
.A1(n_2211),
.A2(n_1961),
.B(n_2024),
.C(n_1962),
.Y(n_2243)
);

O2A1O1Ixp33_ASAP7_75t_L g2244 ( 
.A1(n_2211),
.A2(n_1962),
.B(n_1984),
.C(n_1991),
.Y(n_2244)
);

O2A1O1Ixp33_ASAP7_75t_L g2245 ( 
.A1(n_2217),
.A2(n_1962),
.B(n_1991),
.C(n_1986),
.Y(n_2245)
);

OAI221xp5_ASAP7_75t_SL g2246 ( 
.A1(n_2231),
.A2(n_1962),
.B1(n_2030),
.B2(n_2082),
.C(n_2080),
.Y(n_2246)
);

AOI221xp5_ASAP7_75t_L g2247 ( 
.A1(n_2218),
.A2(n_2206),
.B1(n_2128),
.B2(n_2125),
.C(n_2156),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2212),
.Y(n_2248)
);

AOI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_2210),
.A2(n_2119),
.B1(n_2089),
.B2(n_2095),
.Y(n_2249)
);

OAI221xp5_ASAP7_75t_L g2250 ( 
.A1(n_2214),
.A2(n_2183),
.B1(n_2131),
.B2(n_2157),
.C(n_2156),
.Y(n_2250)
);

AOI32xp33_ASAP7_75t_L g2251 ( 
.A1(n_2235),
.A2(n_2061),
.A3(n_2111),
.B1(n_2107),
.B2(n_2028),
.Y(n_2251)
);

NOR2xp33_ASAP7_75t_L g2252 ( 
.A(n_2224),
.B(n_1781),
.Y(n_2252)
);

AOI211xp5_ASAP7_75t_SL g2253 ( 
.A1(n_2232),
.A2(n_1947),
.B(n_2053),
.C(n_2048),
.Y(n_2253)
);

OAI221xp5_ASAP7_75t_L g2254 ( 
.A1(n_2215),
.A2(n_2183),
.B1(n_2151),
.B2(n_2162),
.C(n_2161),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2216),
.Y(n_2255)
);

AOI221xp5_ASAP7_75t_L g2256 ( 
.A1(n_2238),
.A2(n_2161),
.B1(n_2162),
.B2(n_2157),
.C(n_2151),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2219),
.Y(n_2257)
);

OAI22xp5_ASAP7_75t_L g2258 ( 
.A1(n_2226),
.A2(n_2069),
.B1(n_2061),
.B2(n_2058),
.Y(n_2258)
);

NAND2x1p5_ASAP7_75t_L g2259 ( 
.A(n_2234),
.B(n_2058),
.Y(n_2259)
);

AOI21xp5_ASAP7_75t_L g2260 ( 
.A1(n_2240),
.A2(n_2226),
.B(n_2207),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2247),
.B(n_2221),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2248),
.B(n_2222),
.Y(n_2262)
);

NOR3xp33_ASAP7_75t_L g2263 ( 
.A(n_2246),
.B(n_2228),
.C(n_1895),
.Y(n_2263)
);

NOR2xp67_ASAP7_75t_SL g2264 ( 
.A(n_2250),
.B(n_1843),
.Y(n_2264)
);

OAI221xp5_ASAP7_75t_L g2265 ( 
.A1(n_2253),
.A2(n_2230),
.B1(n_2236),
.B2(n_2237),
.C(n_2229),
.Y(n_2265)
);

NAND3xp33_ASAP7_75t_L g2266 ( 
.A(n_2254),
.B(n_2237),
.C(n_1812),
.Y(n_2266)
);

AOI221xp5_ASAP7_75t_L g2267 ( 
.A1(n_2252),
.A2(n_2227),
.B1(n_2225),
.B2(n_2234),
.C(n_2213),
.Y(n_2267)
);

AOI222xp33_ASAP7_75t_L g2268 ( 
.A1(n_2256),
.A2(n_2233),
.B1(n_2209),
.B2(n_2127),
.C1(n_2129),
.C2(n_2126),
.Y(n_2268)
);

AOI222xp33_ASAP7_75t_L g2269 ( 
.A1(n_2255),
.A2(n_2257),
.B1(n_2258),
.B2(n_2239),
.C1(n_2233),
.C2(n_2129),
.Y(n_2269)
);

OAI221xp5_ASAP7_75t_L g2270 ( 
.A1(n_2251),
.A2(n_1862),
.B1(n_2165),
.B2(n_2114),
.C(n_2188),
.Y(n_2270)
);

INVx1_ASAP7_75t_SL g2271 ( 
.A(n_2259),
.Y(n_2271)
);

AOI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_2249),
.A2(n_2242),
.B1(n_2259),
.B2(n_2103),
.Y(n_2272)
);

OAI211xp5_ASAP7_75t_SL g2273 ( 
.A1(n_2243),
.A2(n_1827),
.B(n_1874),
.C(n_2007),
.Y(n_2273)
);

INVxp67_ASAP7_75t_SL g2274 ( 
.A(n_2245),
.Y(n_2274)
);

NOR2x1_ASAP7_75t_L g2275 ( 
.A(n_2241),
.B(n_1911),
.Y(n_2275)
);

NOR4xp25_ASAP7_75t_SL g2276 ( 
.A(n_2244),
.B(n_1907),
.C(n_1950),
.D(n_1920),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2247),
.B(n_2165),
.Y(n_2277)
);

AOI221xp5_ASAP7_75t_L g2278 ( 
.A1(n_2247),
.A2(n_2126),
.B1(n_2127),
.B2(n_2106),
.C(n_2104),
.Y(n_2278)
);

NAND3xp33_ASAP7_75t_L g2279 ( 
.A(n_2253),
.B(n_1873),
.C(n_1978),
.Y(n_2279)
);

AND4x1_ASAP7_75t_L g2280 ( 
.A(n_2253),
.B(n_1823),
.C(n_1804),
.D(n_1795),
.Y(n_2280)
);

AOI21xp33_ASAP7_75t_L g2281 ( 
.A1(n_2240),
.A2(n_1776),
.B(n_1753),
.Y(n_2281)
);

AOI221xp5_ASAP7_75t_L g2282 ( 
.A1(n_2261),
.A2(n_2094),
.B1(n_2092),
.B2(n_2093),
.C(n_2096),
.Y(n_2282)
);

NAND3xp33_ASAP7_75t_L g2283 ( 
.A(n_2280),
.B(n_2274),
.C(n_2263),
.Y(n_2283)
);

NAND4xp25_ASAP7_75t_L g2284 ( 
.A(n_2260),
.B(n_1795),
.C(n_1867),
.D(n_1804),
.Y(n_2284)
);

NAND4xp75_ASAP7_75t_L g2285 ( 
.A(n_2275),
.B(n_1847),
.C(n_2036),
.D(n_1985),
.Y(n_2285)
);

OAI211xp5_ASAP7_75t_L g2286 ( 
.A1(n_2265),
.A2(n_1774),
.B(n_2058),
.C(n_1923),
.Y(n_2286)
);

NAND3xp33_ASAP7_75t_SL g2287 ( 
.A(n_2276),
.B(n_1896),
.C(n_1920),
.Y(n_2287)
);

NAND4xp25_ASAP7_75t_L g2288 ( 
.A(n_2266),
.B(n_1940),
.C(n_2061),
.D(n_1965),
.Y(n_2288)
);

NOR2xp33_ASAP7_75t_SL g2289 ( 
.A(n_2281),
.B(n_2058),
.Y(n_2289)
);

AOI21xp5_ASAP7_75t_L g2290 ( 
.A1(n_2271),
.A2(n_2032),
.B(n_1923),
.Y(n_2290)
);

NOR3xp33_ASAP7_75t_L g2291 ( 
.A(n_2273),
.B(n_1969),
.C(n_1968),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2269),
.B(n_2139),
.Y(n_2292)
);

NAND4xp25_ASAP7_75t_L g2293 ( 
.A(n_2273),
.B(n_1940),
.C(n_1965),
.D(n_2029),
.Y(n_2293)
);

NAND4xp25_ASAP7_75t_SL g2294 ( 
.A(n_2268),
.B(n_2272),
.C(n_2267),
.D(n_2270),
.Y(n_2294)
);

NOR4xp75_ASAP7_75t_L g2295 ( 
.A(n_2277),
.B(n_2036),
.C(n_1969),
.D(n_1968),
.Y(n_2295)
);

NOR3xp33_ASAP7_75t_L g2296 ( 
.A(n_2279),
.B(n_1969),
.C(n_1968),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2278),
.B(n_2188),
.Y(n_2297)
);

NOR2x1_ASAP7_75t_L g2298 ( 
.A(n_2284),
.B(n_1940),
.Y(n_2298)
);

AND2x4_ASAP7_75t_L g2299 ( 
.A(n_2295),
.B(n_2262),
.Y(n_2299)
);

NOR2x1_ASAP7_75t_L g2300 ( 
.A(n_2283),
.B(n_1816),
.Y(n_2300)
);

NOR4xp25_ASAP7_75t_L g2301 ( 
.A(n_2294),
.B(n_1864),
.C(n_1979),
.D(n_1978),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2297),
.Y(n_2302)
);

AND5x1_ASAP7_75t_L g2303 ( 
.A(n_2289),
.B(n_2282),
.C(n_2291),
.D(n_2296),
.E(n_2290),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2286),
.B(n_2264),
.Y(n_2304)
);

NAND4xp25_ASAP7_75t_L g2305 ( 
.A(n_2288),
.B(n_2007),
.C(n_1965),
.D(n_2002),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2292),
.B(n_2201),
.Y(n_2306)
);

NOR3xp33_ASAP7_75t_L g2307 ( 
.A(n_2293),
.B(n_2287),
.C(n_2285),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2297),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2282),
.B(n_2201),
.Y(n_2309)
);

NAND4xp75_ASAP7_75t_L g2310 ( 
.A(n_2282),
.B(n_1819),
.C(n_1844),
.D(n_1985),
.Y(n_2310)
);

NOR3xp33_ASAP7_75t_L g2311 ( 
.A(n_2283),
.B(n_1850),
.C(n_1801),
.Y(n_2311)
);

NOR3xp33_ASAP7_75t_SL g2312 ( 
.A(n_2283),
.B(n_1853),
.C(n_1955),
.Y(n_2312)
);

NAND4xp25_ASAP7_75t_SL g2313 ( 
.A(n_2283),
.B(n_2104),
.C(n_2106),
.D(n_2103),
.Y(n_2313)
);

NAND4xp25_ASAP7_75t_SL g2314 ( 
.A(n_2300),
.B(n_2049),
.C(n_2082),
.D(n_2080),
.Y(n_2314)
);

NOR4xp25_ASAP7_75t_L g2315 ( 
.A(n_2302),
.B(n_1848),
.C(n_1980),
.D(n_1979),
.Y(n_2315)
);

NAND2x1p5_ASAP7_75t_L g2316 ( 
.A(n_2298),
.B(n_2303),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2310),
.Y(n_2317)
);

NAND4xp25_ASAP7_75t_L g2318 ( 
.A(n_2307),
.B(n_2007),
.C(n_2002),
.D(n_1980),
.Y(n_2318)
);

OAI31xp33_ASAP7_75t_L g2319 ( 
.A1(n_2313),
.A2(n_1750),
.A3(n_2002),
.B(n_1973),
.Y(n_2319)
);

OA22x2_ASAP7_75t_L g2320 ( 
.A1(n_2308),
.A2(n_1816),
.B1(n_2139),
.B2(n_1790),
.Y(n_2320)
);

NAND3xp33_ASAP7_75t_SL g2321 ( 
.A(n_2301),
.B(n_1791),
.C(n_1770),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_2299),
.B(n_2107),
.Y(n_2322)
);

AOI211xp5_ASAP7_75t_SL g2323 ( 
.A1(n_2304),
.A2(n_1727),
.B(n_1810),
.C(n_1791),
.Y(n_2323)
);

OR4x2_ASAP7_75t_L g2324 ( 
.A(n_2312),
.B(n_2069),
.C(n_1974),
.D(n_2000),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2321),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2322),
.Y(n_2326)
);

NOR2xp67_ASAP7_75t_L g2327 ( 
.A(n_2317),
.B(n_2299),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2316),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2320),
.Y(n_2329)
);

AND2x2_ASAP7_75t_SL g2330 ( 
.A(n_2315),
.B(n_2311),
.Y(n_2330)
);

OAI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_2318),
.A2(n_2306),
.B1(n_2309),
.B2(n_2305),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2323),
.B(n_2111),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2314),
.Y(n_2333)
);

XNOR2xp5_ASAP7_75t_L g2334 ( 
.A(n_2327),
.B(n_2324),
.Y(n_2334)
);

OAI22xp5_ASAP7_75t_L g2335 ( 
.A1(n_2328),
.A2(n_2319),
.B1(n_2069),
.B2(n_2046),
.Y(n_2335)
);

INVxp33_ASAP7_75t_L g2336 ( 
.A(n_2328),
.Y(n_2336)
);

OAI22xp5_ASAP7_75t_L g2337 ( 
.A1(n_2329),
.A2(n_2333),
.B1(n_2326),
.B2(n_2330),
.Y(n_2337)
);

AOI21xp5_ASAP7_75t_L g2338 ( 
.A1(n_2325),
.A2(n_2319),
.B(n_1816),
.Y(n_2338)
);

XNOR2x2_ASAP7_75t_L g2339 ( 
.A(n_2331),
.B(n_1983),
.Y(n_2339)
);

XOR2x1_ASAP7_75t_L g2340 ( 
.A(n_2330),
.B(n_1983),
.Y(n_2340)
);

AOI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_2336),
.A2(n_2337),
.B(n_2334),
.Y(n_2341)
);

OAI22xp5_ASAP7_75t_L g2342 ( 
.A1(n_2338),
.A2(n_2332),
.B1(n_2069),
.B2(n_2046),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2339),
.Y(n_2343)
);

OAI22xp5_ASAP7_75t_L g2344 ( 
.A1(n_2341),
.A2(n_2335),
.B1(n_2332),
.B2(n_2340),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_2344),
.B(n_2343),
.Y(n_2345)
);

OR2x6_ASAP7_75t_L g2346 ( 
.A(n_2345),
.B(n_2342),
.Y(n_2346)
);

AOI22xp33_ASAP7_75t_L g2347 ( 
.A1(n_2346),
.A2(n_1989),
.B1(n_2014),
.B2(n_1973),
.Y(n_2347)
);


endmodule