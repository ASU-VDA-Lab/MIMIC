module fake_jpeg_19900_n_325 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx4f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_39),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_11),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_44),
.Y(n_54)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_19),
.A2(n_0),
.B(n_3),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_48),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_39),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_32),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_53),
.A2(n_15),
.B1(n_35),
.B2(n_48),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_31),
.B1(n_33),
.B2(n_20),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_42),
.B1(n_38),
.B2(n_40),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_36),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_29),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_16),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_67),
.B(n_97),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_31),
.B1(n_41),
.B2(n_44),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_17),
.B(n_28),
.C(n_23),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_72),
.B(n_108),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_79),
.Y(n_116)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_74),
.Y(n_118)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_83),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

NAND2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_22),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_82),
.A2(n_87),
.B1(n_93),
.B2(n_104),
.Y(n_138)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_29),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_86),
.Y(n_131)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_18),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_89),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_22),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_92),
.Y(n_142)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_57),
.A2(n_41),
.B1(n_44),
.B2(n_35),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_38),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_45),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_53),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_95),
.B(n_96),
.Y(n_147)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_53),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_99),
.Y(n_136)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_62),
.B1(n_40),
.B2(n_42),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_47),
.B1(n_34),
.B2(n_37),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_27),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_102),
.Y(n_145)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

BUFx8_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_60),
.A2(n_35),
.B1(n_32),
.B2(n_15),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_107),
.Y(n_144)
);

BUFx4f_ASAP7_75t_SL g106 ( 
.A(n_50),
.Y(n_106)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_60),
.B(n_27),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_51),
.B(n_27),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_66),
.A2(n_48),
.B1(n_30),
.B2(n_28),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_30),
.B1(n_23),
.B2(n_11),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_53),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_110),
.A2(n_113),
.B(n_45),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_51),
.B(n_17),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_112),
.Y(n_128)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_55),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_119),
.A2(n_132),
.B1(n_87),
.B2(n_112),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_71),
.B1(n_77),
.B2(n_78),
.Y(n_163)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_105),
.B(n_101),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_68),
.B(n_34),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_140),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_95),
.A2(n_47),
.B1(n_34),
.B2(n_37),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_0),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_47),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_69),
.A2(n_37),
.B1(n_45),
.B2(n_33),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_141),
.A2(n_83),
.B1(n_92),
.B2(n_75),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_72),
.B(n_26),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_105),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_79),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_151),
.B(n_155),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_175),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_105),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_157),
.A2(n_161),
.B(n_180),
.Y(n_200)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_160),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_165),
.B1(n_173),
.B2(n_176),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_10),
.C(n_9),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_113),
.B1(n_98),
.B2(n_96),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_100),
.C(n_74),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_149),
.C(n_133),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_171),
.B1(n_122),
.B2(n_114),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_130),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_169),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_106),
.B(n_24),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_144),
.B(n_141),
.Y(n_184)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_121),
.Y(n_167)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_126),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_106),
.C(n_90),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_133),
.C(n_148),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_85),
.B1(n_33),
.B2(n_26),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_123),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_172),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_124),
.A2(n_26),
.B1(n_20),
.B2(n_24),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_81),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_129),
.A2(n_20),
.B1(n_81),
.B2(n_4),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_119),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_10),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_179),
.Y(n_196)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_144),
.B(n_10),
.CI(n_3),
.CON(n_179),
.SN(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_0),
.B(n_3),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_182),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_116),
.B(n_0),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_180),
.B(n_161),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_154),
.A2(n_143),
.B1(n_146),
.B2(n_138),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_186),
.A2(n_205),
.B1(n_167),
.B2(n_163),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_189),
.B(n_206),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_125),
.B1(n_135),
.B2(n_142),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_190),
.A2(n_201),
.B1(n_209),
.B2(n_139),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_135),
.B(n_147),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_195),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_170),
.A2(n_137),
.B(n_148),
.Y(n_195)
);

AO22x1_ASAP7_75t_L g197 ( 
.A1(n_153),
.A2(n_133),
.B1(n_123),
.B2(n_114),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_207),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_165),
.B1(n_156),
.B2(n_175),
.Y(n_201)
);

XOR2x2_ASAP7_75t_SL g236 ( 
.A(n_202),
.B(n_204),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_179),
.B(n_162),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_131),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_115),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_161),
.A2(n_115),
.B1(n_118),
.B2(n_149),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_118),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_212),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_139),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_7),
.Y(n_237)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_228),
.B(n_233),
.Y(n_249)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_218),
.A2(n_219),
.B1(n_224),
.B2(n_225),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_213),
.B1(n_192),
.B2(n_187),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_220),
.Y(n_254)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_221),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_152),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_223),
.B(n_232),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_164),
.B1(n_169),
.B2(n_174),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_158),
.B1(n_5),
.B2(n_6),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_227),
.A2(n_185),
.B1(n_201),
.B2(n_210),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_R g228 ( 
.A1(n_204),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

OAI21x1_ASAP7_75t_L g233 ( 
.A1(n_191),
.A2(n_4),
.B(n_6),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_234),
.B(n_238),
.Y(n_255)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_237),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_203),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_209),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_212),
.C(n_206),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_257),
.C(n_259),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_242),
.A2(n_218),
.B1(n_239),
.B2(n_222),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_215),
.B(n_196),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_243),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_202),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_246),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_195),
.Y(n_246)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_189),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_256),
.B(n_241),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_200),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_184),
.C(n_197),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_235),
.C(n_215),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_200),
.C(n_227),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_262),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_242),
.A2(n_222),
.B1(n_225),
.B2(n_224),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_268),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_259),
.A2(n_237),
.B(n_214),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_267),
.A2(n_278),
.B(n_257),
.Y(n_281)
);

O2A1O1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_250),
.A2(n_245),
.B(n_258),
.C(n_254),
.Y(n_269)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_244),
.B(n_196),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_270),
.B(n_276),
.Y(n_280)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_271),
.Y(n_284)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_273),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_248),
.A2(n_185),
.B1(n_220),
.B2(n_221),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_247),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_199),
.C(n_211),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_246),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_260),
.B(n_199),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_249),
.A2(n_194),
.B(n_208),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_279),
.B(n_265),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_253),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_286),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_263),
.B(n_240),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_274),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_240),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

NOR3xp33_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_247),
.C(n_208),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_289),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_293),
.B(n_294),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_268),
.C(n_266),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_285),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_275),
.C(n_277),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_291),
.Y(n_308)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_264),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_297),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_308),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_301),
.B(n_284),
.Y(n_305)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_305),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_309),
.B1(n_298),
.B2(n_296),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_307),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_282),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_280),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_300),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_304),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_287),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_318),
.C(n_314),
.Y(n_320)
);

AOI21x1_ASAP7_75t_L g317 ( 
.A1(n_315),
.A2(n_307),
.B(n_299),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_SL g319 ( 
.A1(n_317),
.A2(n_311),
.B(n_267),
.C(n_273),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_319),
.A2(n_320),
.B(n_312),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_321),
.A2(n_290),
.B(n_280),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

NAND2x1_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_270),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_324),
.Y(n_325)
);


endmodule