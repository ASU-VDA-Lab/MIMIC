module fake_jpeg_31844_n_237 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_237);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_7),
.B(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_11),
.B(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_2),
.B(n_3),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_10),
.B(n_4),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_53),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_65),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_17),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_58),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx5_ASAP7_75t_SL g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_1),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g66 ( 
.A(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_67),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_16),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_77),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_34),
.B1(n_18),
.B2(n_22),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_71),
.A2(n_72),
.B1(n_84),
.B2(n_48),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_34),
.B1(n_22),
.B2(n_28),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_41),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_59),
.B1(n_60),
.B2(n_56),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_78),
.A2(n_98),
.B1(n_50),
.B2(n_45),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_22),
.B1(n_28),
.B2(n_38),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_5),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_89),
.C(n_63),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_53),
.B(n_31),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_23),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_35),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_52),
.A2(n_37),
.B1(n_36),
.B2(n_35),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_31),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_37),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_102),
.A2(n_111),
.B1(n_83),
.B2(n_101),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_97),
.B(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_103),
.B(n_131),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_119),
.Y(n_144)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_76),
.A2(n_47),
.B1(n_42),
.B2(n_65),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_107),
.A2(n_122),
.B1(n_82),
.B2(n_91),
.Y(n_148)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_110),
.B(n_102),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_80),
.A2(n_52),
.B1(n_44),
.B2(n_45),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_96),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_113),
.B(n_123),
.Y(n_139)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_32),
.B1(n_20),
.B2(n_27),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_116),
.B1(n_21),
.B2(n_19),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_32),
.B1(n_20),
.B2(n_27),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_96),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_87),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_124),
.Y(n_152)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

NAND2xp33_ASAP7_75t_SL g147 ( 
.A(n_125),
.B(n_126),
.Y(n_147)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_127),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_142)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_129),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_36),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_78),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_23),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_70),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_145),
.C(n_116),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_169)
);

OAI32xp33_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_73),
.A3(n_89),
.B1(n_80),
.B2(n_57),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_57),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_148),
.A2(n_156),
.B1(n_120),
.B2(n_46),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_82),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_158),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_109),
.A2(n_95),
.B1(n_81),
.B2(n_21),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_95),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_107),
.A2(n_81),
.B1(n_62),
.B2(n_63),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_116),
.A2(n_54),
.B1(n_57),
.B2(n_64),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_38),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_176),
.C(n_136),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_121),
.B1(n_105),
.B2(n_127),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_168),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_111),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_118),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_177),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_133),
.B1(n_130),
.B2(n_124),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_172),
.B1(n_154),
.B2(n_152),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_108),
.B1(n_19),
.B2(n_117),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_SL g187 ( 
.A1(n_173),
.A2(n_159),
.B(n_142),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_174),
.A2(n_175),
.B1(n_152),
.B2(n_138),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_96),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_119),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_144),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_179),
.Y(n_184)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_161),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_183),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_96),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_163),
.B(n_154),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_188),
.B1(n_192),
.B2(n_173),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_162),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_190),
.A2(n_172),
.B1(n_169),
.B2(n_183),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_171),
.Y(n_191)
);

AOI211xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_136),
.B(n_147),
.C(n_138),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_169),
.A2(n_152),
.B(n_149),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_155),
.Y(n_200)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_200),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_197),
.A2(n_170),
.B1(n_168),
.B2(n_164),
.Y(n_201)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_205),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_155),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_204),
.B(n_208),
.Y(n_217)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_181),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_197),
.A2(n_165),
.B1(n_178),
.B2(n_7),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_212),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_178),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_210),
.B(n_211),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_5),
.Y(n_211)
);

INVxp33_ASAP7_75t_SL g212 ( 
.A(n_185),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_194),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_206),
.B(n_199),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_221),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_195),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_190),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_223),
.B(n_214),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_199),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_213),
.A2(n_191),
.B1(n_195),
.B2(n_192),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_219),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_224),
.A2(n_214),
.B1(n_196),
.B2(n_193),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_226),
.A2(n_229),
.B1(n_5),
.B2(n_6),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_216),
.B(n_218),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_227),
.A2(n_6),
.B(n_8),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_231),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_228),
.A2(n_9),
.B(n_10),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_232),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_233),
.A2(n_234),
.B(n_15),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_235),
.A2(n_14),
.B1(n_16),
.B2(n_233),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_14),
.Y(n_237)
);


endmodule