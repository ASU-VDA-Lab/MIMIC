module fake_aes_2998_n_846 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_115, n_97, n_80, n_107, n_60, n_114, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_113, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_846);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_115;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_113;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_846;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_840;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_420;
wire n_446;
wire n_165;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_295;
wire n_143;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g116 ( .A(n_48), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_78), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_17), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_16), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_24), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_29), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_33), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_55), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_12), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_71), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_69), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_99), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_58), .Y(n_129) );
BUFx10_ASAP7_75t_L g130 ( .A(n_96), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_108), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_32), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_70), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_63), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_30), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_80), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_52), .Y(n_137) );
INVxp33_ASAP7_75t_SL g138 ( .A(n_46), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_98), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_85), .Y(n_140) );
CKINVDCx14_ASAP7_75t_R g141 ( .A(n_21), .Y(n_141) );
XOR2xp5_ASAP7_75t_L g142 ( .A(n_67), .B(n_42), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_49), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_107), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_25), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_15), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_102), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_41), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_89), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_57), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_54), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_59), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_6), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_103), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_73), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_27), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_50), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_82), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_86), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_64), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_112), .Y(n_161) );
INVx1_ASAP7_75t_SL g162 ( .A(n_37), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_65), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_2), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_110), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_17), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_60), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_28), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_74), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_62), .Y(n_170) );
INVxp67_ASAP7_75t_SL g171 ( .A(n_111), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_81), .Y(n_172) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_130), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_118), .B(n_0), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_152), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_144), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_130), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_122), .Y(n_180) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_119), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_150), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_124), .B(n_0), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_119), .B(n_1), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_122), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_130), .B(n_1), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_142), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_129), .Y(n_188) );
INVxp33_ASAP7_75t_SL g189 ( .A(n_142), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_150), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_166), .B(n_3), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_116), .B(n_4), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_166), .B(n_5), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_144), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_129), .Y(n_195) );
BUFx8_ASAP7_75t_L g196 ( .A(n_131), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_131), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_132), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_132), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_164), .B(n_5), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_146), .B(n_6), .Y(n_201) );
NOR2xp67_ASAP7_75t_L g202 ( .A(n_127), .B(n_7), .Y(n_202) );
OR2x2_ASAP7_75t_L g203 ( .A(n_173), .B(n_146), .Y(n_203) );
INVx1_ASAP7_75t_SL g204 ( .A(n_173), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_198), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_198), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_198), .Y(n_207) );
OR2x2_ASAP7_75t_L g208 ( .A(n_181), .B(n_153), .Y(n_208) );
BUFx10_ASAP7_75t_L g209 ( .A(n_184), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_178), .Y(n_210) );
NAND2xp33_ASAP7_75t_SL g211 ( .A(n_186), .B(n_154), .Y(n_211) );
BUFx4f_ASAP7_75t_L g212 ( .A(n_184), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_181), .B(n_153), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_174), .B(n_138), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_174), .B(n_121), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_174), .B(n_121), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_176), .Y(n_217) );
INVx1_ASAP7_75t_SL g218 ( .A(n_186), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_198), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_174), .B(n_126), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_176), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_198), .Y(n_222) );
NAND3x1_ASAP7_75t_L g223 ( .A(n_186), .B(n_167), .C(n_154), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_179), .B(n_126), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_179), .B(n_135), .Y(n_225) );
NAND2xp33_ASAP7_75t_L g226 ( .A(n_179), .B(n_135), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_198), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_179), .B(n_136), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_196), .B(n_136), .Y(n_229) );
INVx3_ASAP7_75t_L g230 ( .A(n_201), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_176), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_175), .A2(n_172), .B1(n_167), .B2(n_138), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_194), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_184), .B(n_133), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_199), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_201), .Y(n_236) );
OR2x2_ASAP7_75t_L g237 ( .A(n_175), .B(n_139), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_199), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_199), .Y(n_239) );
INVx1_ASAP7_75t_SL g240 ( .A(n_175), .Y(n_240) );
INVxp67_ASAP7_75t_SL g241 ( .A(n_191), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_191), .B(n_139), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_176), .Y(n_243) );
INVx4_ASAP7_75t_L g244 ( .A(n_184), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_193), .B(n_133), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_199), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_201), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_180), .B(n_151), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_230), .A2(n_201), .B1(n_180), .B2(n_188), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_241), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_212), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_242), .Y(n_252) );
BUFx2_ASAP7_75t_L g253 ( .A(n_218), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_242), .B(n_216), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_212), .A2(n_172), .B1(n_189), .B2(n_193), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_216), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_225), .B(n_196), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_225), .B(n_196), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_230), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_212), .A2(n_185), .B(n_188), .C(n_197), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_206), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_208), .A2(n_183), .B(n_200), .C(n_185), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_248), .B(n_196), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_230), .Y(n_264) );
AO22x1_ASAP7_75t_L g265 ( .A1(n_232), .A2(n_187), .B1(n_193), .B2(n_151), .Y(n_265) );
AOI21x1_ASAP7_75t_L g266 ( .A1(n_234), .A2(n_193), .B(n_195), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_209), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_209), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_214), .B(n_191), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_220), .B(n_202), .Y(n_270) );
NAND2x1_ASAP7_75t_L g271 ( .A(n_244), .B(n_195), .Y(n_271) );
INVxp67_ASAP7_75t_L g272 ( .A(n_204), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_240), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_237), .Y(n_274) );
INVx2_ASAP7_75t_SL g275 ( .A(n_209), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_237), .B(n_234), .Y(n_276) );
NAND2x2_ASAP7_75t_L g277 ( .A(n_203), .B(n_208), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_233), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_209), .Y(n_279) );
OR2x2_ASAP7_75t_SL g280 ( .A(n_223), .B(n_187), .Y(n_280) );
OR2x6_ASAP7_75t_L g281 ( .A(n_223), .B(n_183), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_234), .B(n_202), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_244), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_230), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_236), .A2(n_197), .B(n_195), .C(n_182), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_236), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_236), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_221), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_234), .B(n_200), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_272), .B(n_211), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_289), .B(n_213), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_259), .Y(n_292) );
AND2x2_ASAP7_75t_SL g293 ( .A(n_289), .B(n_245), .Y(n_293) );
OR2x6_ASAP7_75t_L g294 ( .A(n_281), .B(n_244), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_L g295 ( .A1(n_254), .A2(n_203), .B(n_247), .C(n_236), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_289), .A2(n_245), .B1(n_244), .B2(n_247), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_253), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_264), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_284), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_286), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_276), .B(n_213), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_279), .Y(n_302) );
HAxp5_ASAP7_75t_L g303 ( .A(n_280), .B(n_210), .CON(n_303), .SN(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_274), .B(n_245), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_287), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_263), .A2(n_245), .B(n_226), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_266), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_283), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_257), .A2(n_224), .B(n_215), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_273), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_252), .B(n_210), .Y(n_311) );
INVx4_ASAP7_75t_L g312 ( .A(n_279), .Y(n_312) );
INVx6_ASAP7_75t_L g313 ( .A(n_279), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_283), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_288), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_256), .B(n_247), .Y(n_316) );
INVxp67_ASAP7_75t_L g317 ( .A(n_273), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_288), .Y(n_318) );
INVx4_ASAP7_75t_L g319 ( .A(n_279), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_267), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_267), .Y(n_321) );
AOI21xp33_ASAP7_75t_L g322 ( .A1(n_255), .A2(n_229), .B(n_228), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_251), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_288), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_293), .B(n_250), .Y(n_325) );
OAI21x1_ASAP7_75t_L g326 ( .A1(n_307), .A2(n_282), .B(n_270), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_307), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_302), .Y(n_328) );
CKINVDCx16_ASAP7_75t_R g329 ( .A(n_297), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_302), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_302), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_294), .B(n_251), .Y(n_332) );
INVx2_ASAP7_75t_SL g333 ( .A(n_302), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_293), .A2(n_249), .B1(n_281), .B2(n_260), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_293), .A2(n_281), .B1(n_277), .B2(n_247), .Y(n_335) );
OAI21x1_ASAP7_75t_L g336 ( .A1(n_306), .A2(n_258), .B(n_262), .Y(n_336) );
OAI21x1_ASAP7_75t_L g337 ( .A1(n_309), .A2(n_197), .B(n_243), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_294), .B(n_268), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_292), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_302), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_294), .A2(n_277), .B1(n_269), .B2(n_249), .Y(n_341) );
AOI21x1_ASAP7_75t_L g342 ( .A1(n_294), .A2(n_243), .B(n_231), .Y(n_342) );
OAI21x1_ASAP7_75t_L g343 ( .A1(n_315), .A2(n_231), .B(n_217), .Y(n_343) );
AOI21xp33_ASAP7_75t_L g344 ( .A1(n_295), .A2(n_260), .B(n_285), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_310), .B(n_265), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_292), .Y(n_346) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_315), .A2(n_217), .B(n_261), .Y(n_347) );
OAI21x1_ASAP7_75t_L g348 ( .A1(n_318), .A2(n_261), .B(n_271), .Y(n_348) );
OAI21x1_ASAP7_75t_L g349 ( .A1(n_318), .A2(n_324), .B(n_299), .Y(n_349) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_324), .A2(n_182), .B(n_190), .Y(n_350) );
OAI21x1_ASAP7_75t_L g351 ( .A1(n_299), .A2(n_182), .B(n_190), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_291), .A2(n_285), .B1(n_190), .B2(n_275), .Y(n_352) );
INVx2_ASAP7_75t_SL g353 ( .A(n_338), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_339), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_329), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_334), .A2(n_310), .B1(n_317), .B2(n_304), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_329), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_341), .A2(n_311), .B1(n_297), .B2(n_290), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_341), .A2(n_334), .B1(n_344), .B2(n_335), .C(n_301), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_325), .B(n_304), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_345), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_335), .A2(n_290), .B1(n_322), .B2(n_278), .Y(n_362) );
AOI222xp33_ASAP7_75t_L g363 ( .A1(n_325), .A2(n_278), .B1(n_303), .B2(n_296), .C1(n_316), .C2(n_192), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_339), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_345), .A2(n_321), .B1(n_320), .B2(n_323), .Y(n_365) );
OA21x2_ASAP7_75t_L g366 ( .A1(n_337), .A2(n_134), .B(n_305), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_345), .A2(n_323), .B1(n_308), .B2(n_305), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_325), .B(n_298), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_332), .B(n_312), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_346), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_344), .A2(n_352), .B1(n_346), .B2(n_303), .C(n_332), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_327), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_352), .A2(n_298), .B(n_300), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_332), .A2(n_308), .B1(n_300), .B2(n_303), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_332), .A2(n_314), .B1(n_321), .B2(n_320), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_338), .A2(n_314), .B1(n_319), .B2(n_312), .Y(n_376) );
NAND3xp33_ASAP7_75t_L g377 ( .A(n_327), .B(n_199), .C(n_176), .Y(n_377) );
AOI22xp33_ASAP7_75t_SL g378 ( .A1(n_338), .A2(n_320), .B1(n_313), .B2(n_319), .Y(n_378) );
OAI22xp33_ASAP7_75t_L g379 ( .A1(n_327), .A2(n_320), .B1(n_319), .B2(n_312), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_338), .A2(n_320), .B1(n_313), .B2(n_275), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_351), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_332), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_351), .Y(n_383) );
OA21x2_ASAP7_75t_L g384 ( .A1(n_337), .A2(n_134), .B(n_205), .Y(n_384) );
BUFx4f_ASAP7_75t_SL g385 ( .A(n_338), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_336), .A2(n_313), .B1(n_268), .B2(n_199), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_336), .A2(n_313), .B1(n_163), .B2(n_117), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_336), .A2(n_120), .B1(n_123), .B2(n_125), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_326), .B(n_168), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_372), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_354), .Y(n_391) );
INVx8_ASAP7_75t_L g392 ( .A(n_369), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_355), .Y(n_393) );
AND2x4_ASAP7_75t_SL g394 ( .A(n_369), .B(n_328), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_366), .Y(n_395) );
OA21x2_ASAP7_75t_L g396 ( .A1(n_381), .A2(n_337), .B(n_326), .Y(n_396) );
NOR2x1p5_ASAP7_75t_L g397 ( .A(n_382), .B(n_389), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_357), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_354), .B(n_351), .Y(n_399) );
BUFx2_ASAP7_75t_L g400 ( .A(n_381), .Y(n_400) );
BUFx3_ASAP7_75t_L g401 ( .A(n_369), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_364), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_372), .Y(n_403) );
NAND2x1_ASAP7_75t_L g404 ( .A(n_383), .B(n_328), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_364), .B(n_350), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_370), .B(n_350), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_370), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_368), .B(n_350), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_363), .B(n_326), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_360), .B(n_340), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_358), .B(n_349), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_374), .B(n_340), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_382), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_383), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_361), .B(n_340), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_359), .B(n_328), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_356), .B(n_330), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_366), .Y(n_418) );
INVx4_ASAP7_75t_SL g419 ( .A(n_385), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_366), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_362), .B(n_349), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_371), .B(n_330), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_366), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_367), .B(n_349), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_353), .B(n_330), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_353), .Y(n_426) );
INVx4_ASAP7_75t_SL g427 ( .A(n_378), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_384), .Y(n_428) );
INVx4_ASAP7_75t_L g429 ( .A(n_384), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_384), .Y(n_430) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_384), .Y(n_431) );
BUFx3_ASAP7_75t_L g432 ( .A(n_376), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_373), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_365), .B(n_331), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_388), .B(n_331), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_376), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_375), .B(n_331), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_387), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_386), .B(n_168), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_380), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_377), .Y(n_441) );
INVx2_ASAP7_75t_SL g442 ( .A(n_379), .Y(n_442) );
AND2x2_ASAP7_75t_SL g443 ( .A(n_381), .B(n_342), .Y(n_443) );
BUFx2_ASAP7_75t_L g444 ( .A(n_381), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_355), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_372), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_361), .B(n_333), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_363), .A2(n_333), .B1(n_137), .B2(n_140), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_363), .B(n_333), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_355), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_369), .Y(n_451) );
BUFx3_ASAP7_75t_L g452 ( .A(n_369), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_355), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_363), .B(n_7), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_391), .Y(n_455) );
OAI31xp33_ASAP7_75t_SL g456 ( .A1(n_397), .A2(n_399), .A3(n_420), .B(n_418), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_413), .B(n_8), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_391), .Y(n_458) );
INVx4_ASAP7_75t_L g459 ( .A(n_419), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_401), .B(n_8), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_401), .B(n_9), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_401), .B(n_9), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_418), .Y(n_463) );
OAI31xp33_ASAP7_75t_SL g464 ( .A1(n_397), .A2(n_171), .A3(n_128), .B(n_158), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_452), .B(n_10), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_402), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_452), .B(n_10), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_402), .B(n_143), .Y(n_468) );
OAI21x1_ASAP7_75t_L g469 ( .A1(n_404), .A2(n_342), .B(n_347), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_407), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_407), .Y(n_471) );
NOR2xp67_ASAP7_75t_L g472 ( .A(n_429), .B(n_11), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_390), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_454), .B(n_145), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_403), .Y(n_475) );
BUFx2_ASAP7_75t_L g476 ( .A(n_392), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_448), .A2(n_170), .B(n_148), .C(n_149), .Y(n_477) );
AOI33xp33_ASAP7_75t_L g478 ( .A1(n_436), .A2(n_147), .A3(n_155), .B1(n_156), .B2(n_157), .B3(n_159), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_393), .B(n_160), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_452), .B(n_11), .Y(n_480) );
NOR2xp33_ASAP7_75t_SL g481 ( .A(n_392), .B(n_162), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_398), .B(n_161), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_446), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_410), .B(n_12), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_446), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_410), .B(n_13), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_445), .B(n_13), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_446), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_450), .B(n_14), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_432), .B(n_342), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_453), .Y(n_491) );
BUFx3_ASAP7_75t_L g492 ( .A(n_392), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_399), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_449), .A2(n_165), .B1(n_169), .B2(n_176), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_432), .B(n_348), .Y(n_495) );
OA211x2_ASAP7_75t_L g496 ( .A1(n_409), .A2(n_14), .B(n_15), .C(n_16), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_432), .B(n_348), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_400), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_451), .B(n_18), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_392), .B(n_18), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_423), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_423), .Y(n_502) );
INVx3_ASAP7_75t_L g503 ( .A(n_395), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_392), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_451), .B(n_19), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_438), .B(n_19), .Y(n_506) );
INVx4_ASAP7_75t_L g507 ( .A(n_419), .Y(n_507) );
OAI31xp33_ASAP7_75t_L g508 ( .A1(n_438), .A2(n_221), .A3(n_205), .B(n_227), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_414), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_415), .B(n_20), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_395), .B(n_177), .Y(n_511) );
INVxp67_ASAP7_75t_SL g512 ( .A(n_395), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_451), .B(n_20), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_405), .Y(n_514) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_395), .Y(n_515) );
INVx3_ASAP7_75t_L g516 ( .A(n_395), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_405), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_414), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_451), .B(n_21), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_436), .A2(n_348), .B1(n_347), .B2(n_343), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_414), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_406), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_440), .B(n_177), .C(n_206), .Y(n_523) );
OAI22xp5_ASAP7_75t_SL g524 ( .A1(n_419), .A2(n_22), .B1(n_177), .B2(n_26), .Y(n_524) );
INVx5_ASAP7_75t_SL g525 ( .A(n_395), .Y(n_525) );
INVxp67_ASAP7_75t_L g526 ( .A(n_420), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_400), .Y(n_527) );
BUFx3_ASAP7_75t_L g528 ( .A(n_394), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_428), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_406), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_415), .B(n_22), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_447), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_427), .B(n_343), .Y(n_533) );
OAI22xp5_ASAP7_75t_SL g534 ( .A1(n_419), .A2(n_177), .B1(n_31), .B2(n_34), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_447), .Y(n_535) );
BUFx3_ASAP7_75t_L g536 ( .A(n_394), .Y(n_536) );
NAND3xp33_ASAP7_75t_L g537 ( .A(n_422), .B(n_177), .C(n_222), .Y(n_537) );
NOR2xp67_ASAP7_75t_L g538 ( .A(n_429), .B(n_23), .Y(n_538) );
AND2x2_ASAP7_75t_SL g539 ( .A(n_429), .B(n_177), .Y(n_539) );
BUFx2_ASAP7_75t_L g540 ( .A(n_419), .Y(n_540) );
BUFx3_ASAP7_75t_L g541 ( .A(n_394), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_426), .B(n_221), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_408), .B(n_35), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_428), .Y(n_544) );
NAND2xp67_ASAP7_75t_L g545 ( .A(n_422), .B(n_36), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_444), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_428), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_416), .B(n_343), .Y(n_548) );
NAND3xp33_ASAP7_75t_L g549 ( .A(n_416), .B(n_206), .C(n_207), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_444), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_412), .B(n_38), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_430), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_412), .B(n_39), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_417), .B(n_246), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_417), .B(n_246), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_425), .B(n_40), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_552), .Y(n_557) );
NAND4xp25_ASAP7_75t_L g558 ( .A(n_464), .B(n_421), .C(n_411), .D(n_424), .Y(n_558) );
INVx1_ASAP7_75t_SL g559 ( .A(n_552), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_491), .B(n_484), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_481), .A2(n_427), .B1(n_442), .B2(n_435), .Y(n_561) );
INVx2_ASAP7_75t_SL g562 ( .A(n_492), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_514), .B(n_430), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_486), .B(n_493), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_498), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_455), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_517), .B(n_430), .Y(n_567) );
AND2x2_ASAP7_75t_SL g568 ( .A(n_456), .B(n_429), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_522), .B(n_434), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_530), .B(n_425), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_458), .B(n_433), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_498), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_527), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_532), .B(n_425), .Y(n_574) );
NAND2xp33_ASAP7_75t_SL g575 ( .A(n_459), .B(n_404), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_535), .B(n_434), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_466), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_543), .B(n_425), .Y(n_578) );
OR2x6_ASAP7_75t_L g579 ( .A(n_528), .B(n_431), .Y(n_579) );
OAI33xp33_ASAP7_75t_L g580 ( .A1(n_474), .A2(n_433), .A3(n_439), .B1(n_441), .B2(n_227), .B3(n_235), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_470), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_471), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_476), .B(n_427), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_528), .B(n_427), .Y(n_584) );
AND2x4_ASAP7_75t_L g585 ( .A(n_536), .B(n_427), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_536), .B(n_435), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_527), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_463), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_463), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_541), .B(n_443), .Y(n_590) );
OAI31xp33_ASAP7_75t_L g591 ( .A1(n_477), .A2(n_442), .A3(n_437), .B(n_441), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_526), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_541), .B(n_461), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_465), .B(n_443), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_539), .Y(n_595) );
INVxp67_ASAP7_75t_L g596 ( .A(n_472), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_526), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_546), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_550), .B(n_443), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_539), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_509), .B(n_431), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_509), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_467), .B(n_437), .Y(n_603) );
AND2x4_ASAP7_75t_SL g604 ( .A(n_459), .B(n_437), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_480), .B(n_457), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_473), .B(n_475), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_518), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_487), .B(n_437), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_489), .B(n_431), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_521), .B(n_431), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_492), .B(n_396), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_521), .B(n_396), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_485), .B(n_396), .Y(n_613) );
INVxp67_ASAP7_75t_SL g614 ( .A(n_512), .Y(n_614) );
AND2x4_ASAP7_75t_L g615 ( .A(n_495), .B(n_43), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_488), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_483), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_551), .B(n_396), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_501), .B(n_44), .Y(n_619) );
OAI322xp33_ASAP7_75t_L g620 ( .A1(n_506), .A2(n_239), .A3(n_235), .B1(n_219), .B2(n_222), .C1(n_238), .C2(n_207), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_505), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_513), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_529), .B(n_239), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_501), .B(n_45), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_502), .B(n_47), .Y(n_625) );
AND2x4_ASAP7_75t_SL g626 ( .A(n_459), .B(n_288), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_553), .B(n_51), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_504), .B(n_53), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_510), .B(n_56), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_502), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_529), .B(n_219), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_554), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_555), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_499), .B(n_61), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_479), .B(n_66), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_460), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_519), .B(n_68), .Y(n_637) );
AOI211xp5_ASAP7_75t_L g638 ( .A1(n_500), .A2(n_238), .B(n_222), .C(n_207), .Y(n_638) );
OA211x2_ASAP7_75t_L g639 ( .A1(n_511), .A2(n_72), .B(n_75), .C(n_76), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_544), .B(n_77), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_544), .B(n_238), .Y(n_641) );
NAND2x1p5_ASAP7_75t_SL g642 ( .A(n_556), .B(n_79), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_511), .A2(n_238), .B(n_222), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_547), .B(n_83), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_531), .B(n_87), .Y(n_645) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_512), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_495), .B(n_88), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_515), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_495), .B(n_90), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_525), .Y(n_650) );
NOR3xp33_ASAP7_75t_L g651 ( .A(n_478), .B(n_91), .C(n_92), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_525), .B(n_93), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_515), .Y(n_653) );
NOR2xp67_ASAP7_75t_L g654 ( .A(n_507), .B(n_94), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_525), .B(n_95), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_548), .B(n_238), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_482), .B(n_97), .Y(n_657) );
AND2x2_ASAP7_75t_SL g658 ( .A(n_507), .B(n_100), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_497), .B(n_101), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_462), .B(n_104), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_503), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g662 ( .A1(n_477), .A2(n_222), .B1(n_207), .B2(n_206), .C(n_113), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_503), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_507), .B(n_206), .Y(n_664) );
OAI31xp33_ASAP7_75t_L g665 ( .A1(n_524), .A2(n_105), .A3(n_106), .B(n_109), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_566), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_577), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_581), .Y(n_668) );
OAI21xp5_ASAP7_75t_L g669 ( .A1(n_651), .A2(n_478), .B(n_549), .Y(n_669) );
INVx1_ASAP7_75t_SL g670 ( .A(n_559), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_632), .B(n_497), .Y(n_671) );
INVxp67_ASAP7_75t_L g672 ( .A(n_560), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_582), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_588), .B(n_497), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_569), .B(n_516), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_608), .B(n_490), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_603), .B(n_490), .Y(n_677) );
INVx3_ASAP7_75t_L g678 ( .A(n_585), .Y(n_678) );
NOR2x1_ASAP7_75t_R g679 ( .A(n_585), .B(n_540), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_589), .Y(n_680) );
NAND4xp25_ASAP7_75t_L g681 ( .A(n_591), .B(n_496), .C(n_468), .D(n_494), .Y(n_681) );
NAND2xp33_ASAP7_75t_SL g682 ( .A(n_562), .B(n_534), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_592), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_609), .B(n_490), .Y(n_684) );
OAI21xp5_ASAP7_75t_SL g685 ( .A1(n_595), .A2(n_533), .B(n_537), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_564), .B(n_533), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_586), .B(n_533), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_605), .B(n_516), .Y(n_688) );
OR2x6_ASAP7_75t_L g689 ( .A(n_579), .B(n_516), .Y(n_689) );
INVxp67_ASAP7_75t_L g690 ( .A(n_557), .Y(n_690) );
INVx2_ASAP7_75t_SL g691 ( .A(n_626), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_658), .A2(n_538), .B1(n_523), .B2(n_520), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_593), .B(n_542), .Y(n_693) );
INVx1_ASAP7_75t_SL g694 ( .A(n_557), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_576), .B(n_469), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_633), .B(n_545), .Y(n_696) );
BUFx2_ASAP7_75t_L g697 ( .A(n_575), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_561), .A2(n_469), .B1(n_207), .B2(n_508), .Y(n_698) );
INVx2_ASAP7_75t_SL g699 ( .A(n_604), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_597), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_598), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_594), .B(n_114), .Y(n_702) );
AND2x4_ASAP7_75t_L g703 ( .A(n_611), .B(n_115), .Y(n_703) );
AOI211x1_ASAP7_75t_SL g704 ( .A1(n_558), .A2(n_599), .B(n_654), .C(n_571), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_570), .B(n_578), .Y(n_705) );
AND2x4_ASAP7_75t_L g706 ( .A(n_579), .B(n_587), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_616), .Y(n_707) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_565), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_574), .B(n_590), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_568), .B(n_583), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_636), .B(n_621), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_573), .B(n_587), .Y(n_712) );
INVx2_ASAP7_75t_SL g713 ( .A(n_606), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_567), .B(n_565), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_571), .Y(n_715) );
INVxp67_ASAP7_75t_SL g716 ( .A(n_646), .Y(n_716) );
OAI22xp33_ASAP7_75t_L g717 ( .A1(n_595), .A2(n_600), .B1(n_662), .B2(n_596), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_646), .Y(n_718) );
INVx1_ASAP7_75t_SL g719 ( .A(n_573), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_567), .B(n_572), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_648), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_572), .B(n_602), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_584), .B(n_600), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_563), .Y(n_724) );
AND2x4_ASAP7_75t_L g725 ( .A(n_579), .B(n_614), .Y(n_725) );
INVx1_ASAP7_75t_SL g726 ( .A(n_648), .Y(n_726) );
AO21x1_ASAP7_75t_L g727 ( .A1(n_651), .A2(n_638), .B(n_614), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_622), .B(n_618), .Y(n_728) );
BUFx2_ASAP7_75t_L g729 ( .A(n_650), .Y(n_729) );
OR2x2_ASAP7_75t_L g730 ( .A(n_599), .B(n_630), .Y(n_730) );
INVx1_ASAP7_75t_SL g731 ( .A(n_653), .Y(n_731) );
NOR2x1_ASAP7_75t_L g732 ( .A(n_664), .B(n_655), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_607), .B(n_617), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_653), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_613), .B(n_612), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_613), .B(n_612), .Y(n_736) );
O2A1O1Ixp33_ASAP7_75t_L g737 ( .A1(n_596), .A2(n_662), .B(n_657), .C(n_635), .Y(n_737) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_601), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_647), .B(n_659), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_682), .A2(n_629), .B1(n_580), .B2(n_645), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_666), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_688), .B(n_661), .Y(n_742) );
INVxp67_ASAP7_75t_L g743 ( .A(n_729), .Y(n_743) );
INVxp67_ASAP7_75t_L g744 ( .A(n_712), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_696), .A2(n_629), .B1(n_580), .B2(n_615), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_713), .B(n_656), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_667), .Y(n_747) );
OAI221xp5_ASAP7_75t_L g748 ( .A1(n_704), .A2(n_665), .B1(n_660), .B2(n_652), .C(n_649), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_726), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_668), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_673), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_701), .Y(n_752) );
AOI31xp33_ASAP7_75t_L g753 ( .A1(n_679), .A2(n_627), .A3(n_615), .B(n_637), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_714), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_728), .B(n_656), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_727), .A2(n_643), .B(n_620), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_714), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_681), .A2(n_634), .B1(n_628), .B2(n_639), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_720), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_715), .B(n_663), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_720), .Y(n_761) );
AND3x2_ASAP7_75t_L g762 ( .A(n_697), .B(n_642), .C(n_601), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_707), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_680), .Y(n_764) );
AOI221x1_ASAP7_75t_SL g765 ( .A1(n_717), .A2(n_610), .B1(n_631), .B2(n_623), .C(n_641), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_672), .B(n_610), .Y(n_766) );
NAND3xp33_ASAP7_75t_L g767 ( .A(n_708), .B(n_643), .C(n_619), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_683), .Y(n_768) );
AOI222xp33_ASAP7_75t_L g769 ( .A1(n_711), .A2(n_623), .B1(n_631), .B2(n_625), .C1(n_624), .C2(n_640), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_700), .Y(n_770) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_726), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_724), .B(n_644), .Y(n_772) );
OAI32xp33_ASAP7_75t_L g773 ( .A1(n_710), .A2(n_692), .A3(n_678), .B1(n_731), .B2(n_695), .Y(n_773) );
NAND2xp33_ASAP7_75t_SL g774 ( .A(n_699), .B(n_678), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_669), .A2(n_692), .B1(n_732), .B2(n_739), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_735), .B(n_736), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_735), .B(n_736), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_681), .A2(n_686), .B1(n_671), .B2(n_693), .Y(n_778) );
NAND2x1p5_ASAP7_75t_L g779 ( .A(n_691), .B(n_703), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_722), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_690), .B(n_738), .Y(n_781) );
AOI221xp5_ASAP7_75t_L g782 ( .A1(n_737), .A2(n_674), .B1(n_716), .B2(n_722), .C(n_694), .Y(n_782) );
NAND2x1p5_ASAP7_75t_L g783 ( .A(n_703), .B(n_670), .Y(n_783) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_731), .Y(n_784) );
NOR2x1_ASAP7_75t_L g785 ( .A(n_685), .B(n_669), .Y(n_785) );
NOR2xp67_ASAP7_75t_L g786 ( .A(n_775), .B(n_685), .Y(n_786) );
AOI221xp5_ASAP7_75t_L g787 ( .A1(n_775), .A2(n_674), .B1(n_719), .B2(n_705), .C(n_694), .Y(n_787) );
OAI21xp33_ASAP7_75t_L g788 ( .A1(n_785), .A2(n_677), .B(n_676), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g789 ( .A(n_774), .B(n_725), .Y(n_789) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_753), .A2(n_778), .B1(n_779), .B2(n_740), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_780), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_745), .A2(n_723), .B1(n_706), .B2(n_684), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_754), .Y(n_793) );
INVxp67_ASAP7_75t_L g794 ( .A(n_771), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_757), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_744), .B(n_687), .Y(n_796) );
AND2x2_ASAP7_75t_SL g797 ( .A(n_782), .B(n_725), .Y(n_797) );
AOI221xp5_ASAP7_75t_L g798 ( .A1(n_773), .A2(n_719), .B1(n_670), .B2(n_709), .C(n_706), .Y(n_798) );
O2A1O1Ixp5_ASAP7_75t_L g799 ( .A1(n_756), .A2(n_718), .B(n_721), .C(n_734), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_759), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_761), .Y(n_801) );
INVx2_ASAP7_75t_SL g802 ( .A(n_742), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_749), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_779), .A2(n_689), .B1(n_698), .B2(n_675), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_776), .Y(n_805) );
INVx1_ASAP7_75t_SL g806 ( .A(n_781), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_776), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_777), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_777), .B(n_730), .Y(n_809) );
XNOR2x1_ASAP7_75t_L g810 ( .A(n_762), .B(n_702), .Y(n_810) );
AOI21xp33_ASAP7_75t_L g811 ( .A1(n_790), .A2(n_758), .B(n_748), .Y(n_811) );
INVxp67_ASAP7_75t_L g812 ( .A(n_806), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_788), .B(n_743), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_791), .Y(n_814) );
OAI21x1_ASAP7_75t_SL g815 ( .A1(n_787), .A2(n_765), .B(n_746), .Y(n_815) );
OAI21xp33_ASAP7_75t_L g816 ( .A1(n_797), .A2(n_786), .B(n_798), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_793), .Y(n_817) );
OAI22xp33_ASAP7_75t_L g818 ( .A1(n_789), .A2(n_783), .B1(n_689), .B2(n_755), .Y(n_818) );
AND2x2_ASAP7_75t_L g819 ( .A(n_805), .B(n_784), .Y(n_819) );
INVx1_ASAP7_75t_SL g820 ( .A(n_789), .Y(n_820) );
AOI21xp33_ASAP7_75t_SL g821 ( .A1(n_797), .A2(n_783), .B(n_767), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_807), .B(n_808), .Y(n_822) );
AOI222xp33_ASAP7_75t_L g823 ( .A1(n_794), .A2(n_766), .B1(n_763), .B2(n_741), .C1(n_747), .C2(n_750), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_822), .Y(n_824) );
OAI221xp5_ASAP7_75t_SL g825 ( .A1(n_816), .A2(n_792), .B1(n_794), .B2(n_809), .C(n_769), .Y(n_825) );
NAND4xp25_ASAP7_75t_L g826 ( .A(n_811), .B(n_799), .C(n_804), .D(n_772), .Y(n_826) );
NAND3xp33_ASAP7_75t_L g827 ( .A(n_821), .B(n_799), .C(n_810), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_823), .B(n_795), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_822), .B(n_801), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_819), .B(n_800), .Y(n_830) );
NOR3xp33_ASAP7_75t_L g831 ( .A(n_825), .B(n_818), .C(n_820), .Y(n_831) );
NOR4xp75_ASAP7_75t_SL g832 ( .A(n_828), .B(n_815), .C(n_813), .D(n_812), .Y(n_832) );
NOR3xp33_ASAP7_75t_L g833 ( .A(n_827), .B(n_813), .C(n_817), .Y(n_833) );
OR2x2_ASAP7_75t_L g834 ( .A(n_824), .B(n_814), .Y(n_834) );
AND5x1_ASAP7_75t_L g835 ( .A(n_831), .B(n_826), .C(n_830), .D(n_829), .E(n_819), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_834), .Y(n_836) );
NOR3xp33_ASAP7_75t_L g837 ( .A(n_833), .B(n_770), .C(n_768), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_836), .A2(n_832), .B1(n_837), .B2(n_835), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_837), .B(n_752), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_839), .Y(n_840) );
XOR2xp5_ASAP7_75t_L g841 ( .A(n_838), .B(n_796), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_840), .B(n_751), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_841), .A2(n_803), .B(n_802), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_843), .A2(n_803), .B1(n_764), .B2(n_689), .Y(n_844) );
XNOR2xp5_ASAP7_75t_L g845 ( .A(n_844), .B(n_842), .Y(n_845) );
AOI21xp5_ASAP7_75t_L g846 ( .A1(n_845), .A2(n_760), .B(n_733), .Y(n_846) );
endmodule