module fake_jpeg_28664_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_8),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_13),
.B(n_29),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_50),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_62),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_59),
.Y(n_66)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_43),
.B(n_0),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_63),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_53),
.C(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_55),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_74),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_85),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_74),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_82),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_72),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_87),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_68),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_90),
.Y(n_95)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_39),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_39),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_90),
.A2(n_45),
.B1(n_48),
.B2(n_39),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_80),
.B1(n_15),
.B2(n_20),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_99),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_40),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_103),
.B(n_109),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_6),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_104),
.Y(n_115)
);

NOR2x1_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_41),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_9),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_26),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_10),
.B(n_12),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_110),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_14),
.B1(n_22),
.B2(n_23),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_117),
.B1(n_121),
.B2(n_36),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_94),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_114),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_24),
.B(n_25),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_120),
.B(n_31),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_102),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_93),
.B1(n_92),
.B2(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_30),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_109),
.B1(n_33),
.B2(n_35),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_125),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_119),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g129 ( 
.A1(n_128),
.A2(n_116),
.B(n_115),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_129),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_127),
.B(n_124),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_123),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_132),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);


endmodule