module fake_jpeg_30947_n_34 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_34);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_34;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_13),
.B(n_1),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_20),
.B(n_21),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_18),
.B(n_13),
.Y(n_23)
);

A2O1A1O1Ixp25_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_25),
.B(n_16),
.C(n_15),
.D(n_3),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_16),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_15),
.C(n_17),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_15),
.B(n_17),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_28),
.C(n_29),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_11),
.B1(n_9),
.B2(n_4),
.Y(n_29)
);

INVxp33_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

AOI322xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_22),
.A3(n_24),
.B1(n_4),
.B2(n_5),
.C1(n_2),
.C2(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

OAI221xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_31),
.B1(n_5),
.B2(n_6),
.C(n_8),
.Y(n_34)
);


endmodule