module real_jpeg_31442_n_16 (n_5, n_4, n_8, n_0, n_12, n_463, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_463;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_0),
.Y(n_173)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_0),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_0),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g333 ( 
.A(n_0),
.Y(n_333)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_1),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_1),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_1),
.B(n_130),
.Y(n_197)
);

OAI32xp33_ASAP7_75t_L g311 ( 
.A1(n_1),
.A2(n_312),
.A3(n_315),
.B1(n_317),
.B2(n_322),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_1),
.A2(n_161),
.B1(n_357),
.B2(n_360),
.Y(n_356)
);

OAI21xp33_ASAP7_75t_L g389 ( 
.A1(n_1),
.A2(n_183),
.B(n_390),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_2),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_2),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_2),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_3),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_3),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_3),
.A2(n_58),
.B1(n_122),
.B2(n_127),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g205 ( 
.A1(n_3),
.A2(n_58),
.B1(n_206),
.B2(n_210),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_3),
.A2(n_58),
.B1(n_336),
.B2(n_339),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_4),
.Y(n_182)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_4),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_5),
.Y(n_96)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_5),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_6),
.A2(n_235),
.B1(n_237),
.B2(n_238),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_6),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_7),
.A2(n_175),
.B1(n_179),
.B2(n_180),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_7),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_7),
.A2(n_179),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_9),
.Y(n_134)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_9),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_10),
.A2(n_108),
.B1(n_115),
.B2(n_116),
.Y(n_107)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_10),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_10),
.A2(n_115),
.B1(n_275),
.B2(n_281),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_10),
.A2(n_115),
.B1(n_363),
.B2(n_366),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_10),
.A2(n_115),
.B1(n_378),
.B2(n_382),
.Y(n_377)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_12),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_12),
.Y(n_88)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_12),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_13),
.A2(n_248),
.B1(n_251),
.B2(n_254),
.Y(n_247)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_13),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_14),
.A2(n_66),
.B1(n_71),
.B2(n_72),
.Y(n_65)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_14),
.A2(n_71),
.B1(n_192),
.B2(n_195),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_15),
.A2(n_77),
.B1(n_83),
.B2(n_84),
.Y(n_76)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_15),
.A2(n_83),
.B1(n_303),
.B2(n_306),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_15),
.A2(n_83),
.B1(n_408),
.B2(n_410),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_290),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_288),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_241),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_21),
.B(n_241),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_166),
.C(n_215),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_22),
.B(n_342),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_119),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_74),
.Y(n_23)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_24),
.B(n_74),
.C(n_119),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_53),
.B1(n_61),
.B2(n_64),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_25),
.B(n_440),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_25),
.A2(n_53),
.B1(n_309),
.B2(n_450),
.Y(n_449)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_26),
.A2(n_62),
.B1(n_65),
.B2(n_259),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_SL g301 ( 
.A1(n_26),
.A2(n_302),
.B(n_308),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_26),
.A2(n_62),
.B1(n_302),
.B2(n_362),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_41),
.Y(n_26)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

OAI22x1_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_35),
.B2(n_38),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_29),
.Y(n_384)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_34),
.Y(n_425)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_36),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_38),
.Y(n_340)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_40),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_40),
.Y(n_338)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_40),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_41)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_42),
.Y(n_316)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_49),
.Y(n_307)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_49),
.Y(n_365)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_53),
.B(n_309),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_56),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_57),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g431 ( 
.A(n_57),
.Y(n_431)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_63),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_63),
.B(n_161),
.Y(n_375)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_70),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_73),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_89),
.B1(n_100),
.B2(n_107),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OA21x2_ASAP7_75t_L g269 ( 
.A1(n_76),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_81),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_82),
.Y(n_209)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_97),
.B1(n_102),
.B2(n_106),
.Y(n_101)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_90),
.B(n_161),
.Y(n_451)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_91),
.B(n_107),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_91),
.B(n_205),
.Y(n_271)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_92)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_96),
.Y(n_328)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_100),
.B(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_100),
.Y(n_270)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_114),
.Y(n_214)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_143),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_130),
.Y(n_120)
);

NAND2x1_ASAP7_75t_SL g284 ( 
.A(n_121),
.B(n_144),
.Y(n_284)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_146),
.B1(n_149),
.B2(n_151),
.Y(n_145)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_126),
.Y(n_129)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_126),
.Y(n_283)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_130),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_135),
.B1(n_137),
.B2(n_140),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_134),
.Y(n_229)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_136),
.Y(n_359)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_140),
.Y(n_226)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_142),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_142),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_155),
.Y(n_143)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_150),
.Y(n_220)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_161),
.B(n_162),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_161),
.B(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_161),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_161),
.B(n_428),
.Y(n_427)
);

OAI21xp33_ASAP7_75t_SL g440 ( 
.A1(n_161),
.A2(n_427),
.B(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI32xp33_ASAP7_75t_L g216 ( 
.A1(n_163),
.A2(n_217),
.A3(n_219),
.B1(n_221),
.B2(n_224),
.Y(n_216)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_167),
.A2(n_215),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_197),
.B1(n_198),
.B2(n_201),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_197),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_168),
.B(n_197),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_168),
.A2(n_197),
.B1(n_198),
.B2(n_201),
.Y(n_345)
);

OAI22x1_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_174),
.B1(n_183),
.B2(n_191),
.Y(n_168)
);

INVx3_ASAP7_75t_SL g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_173),
.Y(n_395)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_178),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_181),
.Y(n_412)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_183),
.A2(n_246),
.B1(n_247),
.B2(n_255),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_183),
.A2(n_390),
.B(n_407),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_184),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_184),
.B(n_335),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_184),
.A2(n_256),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

BUFx4f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_187),
.Y(n_401)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_190),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_191),
.A2(n_330),
.B(n_334),
.Y(n_329)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_200),
.B(n_202),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_211),
.Y(n_324)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_215),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_230),
.B1(n_231),
.B2(n_240),
.Y(n_215)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

BUFx4f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_230),
.B(n_240),
.Y(n_287)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_239),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_267),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_258),
.Y(n_244)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_250),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_257),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

XNOR2x1_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_287),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_272),
.B1(n_285),
.B2(n_286),
.Y(n_268)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_270),
.A2(n_271),
.B(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_284),
.Y(n_272)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI21x1_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_346),
.B(n_460),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_341),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_295),
.B(n_461),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_300),
.C(n_310),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_297),
.B(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_300),
.A2(n_301),
.B1(n_310),
.B2(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_305),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_308),
.B(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_310),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_329),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_311),
.B(n_329),
.Y(n_353)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_325),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_331),
.Y(n_330)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx8_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_334),
.A2(n_377),
.B(n_385),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_335),
.B(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_341),
.Y(n_461)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_371),
.B(n_459),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_351),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_348),
.B(n_351),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_354),
.C(n_361),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_353),
.B(n_445),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_355),
.B(n_361),
.Y(n_445)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_362),
.Y(n_450)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx3_ASAP7_75t_SL g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

OAI321xp33_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_443),
.A3(n_452),
.B1(n_457),
.B2(n_458),
.C(n_463),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_403),
.B(n_442),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_374),
.A2(n_388),
.B(n_402),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_375),
.B(n_376),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_377),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

BUFx2_ASAP7_75t_SL g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_396),
.Y(n_388)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_399),
.Y(n_396)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_413),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_404),
.B(n_413),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_438),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_414),
.B(n_438),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_426),
.B1(n_432),
.B2(n_437),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_420),
.Y(n_415)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_416),
.Y(n_437)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx6_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_435),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_434),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

AND2x2_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_446),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_446),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.C(n_451),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_455),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_448),
.A2(n_449),
.B1(n_451),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_451),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_SL g457 ( 
.A(n_453),
.B(n_454),
.Y(n_457)
);


endmodule