module real_jpeg_30685_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_12;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_0),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_0),
.B(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_0),
.A2(n_60),
.B1(n_93),
.B2(n_95),
.Y(n_92)
);

AOI22x1_ASAP7_75t_L g126 ( 
.A1(n_0),
.A2(n_60),
.B1(n_127),
.B2(n_131),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_0),
.A2(n_138),
.A3(n_143),
.B1(n_146),
.B2(n_154),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_0),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_0),
.B(n_124),
.Y(n_272)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_1),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_1),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_2),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_2),
.Y(n_192)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_4),
.Y(n_82)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_4),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_4),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_5),
.A2(n_303),
.B1(n_306),
.B2(n_307),
.Y(n_302)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_5),
.Y(n_306)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_6),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_6),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

OAI22x1_ASAP7_75t_SL g21 ( 
.A1(n_8),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_21)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_8),
.A2(n_26),
.B1(n_79),
.B2(n_83),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_8),
.A2(n_26),
.B1(n_117),
.B2(n_120),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_8),
.A2(n_26),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_9),
.Y(n_102)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_9),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_289),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

OAI21x1_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_233),
.B(n_288),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_163),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_16),
.B(n_163),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_97),
.C(n_135),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_17),
.B(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_62),
.B2(n_63),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_18),
.B(n_64),
.C(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_18),
.B(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OA22x2_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_30),
.B1(n_46),
.B2(n_56),
.Y(n_19)
);

INVxp67_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22x1_ASAP7_75t_L g230 ( 
.A1(n_21),
.A2(n_31),
.B1(n_57),
.B2(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_24),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

AND2x4_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_46),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_39),
.B2(n_42),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_41),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_41),
.Y(n_189)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_45),
.Y(n_153)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_46),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_46),
.B(n_60),
.Y(n_258)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_49),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_49),
.Y(n_159)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_60),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_60),
.B(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_60),
.A2(n_190),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_60),
.B(n_240),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_L g247 ( 
.A1(n_60),
.A2(n_104),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_73),
.B(n_96),
.Y(n_63)
);

OAI211xp5_ASAP7_75t_L g96 ( 
.A1(n_64),
.A2(n_74),
.B(n_77),
.C(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_65),
.Y(n_204)
);

NOR2x1_ASAP7_75t_L g215 ( 
.A(n_65),
.B(n_216),
.Y(n_215)
);

AO22x1_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_68),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_68),
.Y(n_219)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_73),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_73),
.B(n_266),
.Y(n_265)
);

OA21x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B(n_87),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_75),
.Y(n_196)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_78),
.A2(n_88),
.B1(n_92),
.B2(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_82),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_82),
.Y(n_305)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_107),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_86),
.Y(n_251)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_86),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_87),
.A2(n_302),
.B(n_311),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_89),
.B(n_162),
.Y(n_161)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_92),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_97),
.A2(n_98),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_97),
.B(n_193),
.C(n_258),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_97),
.A2(n_135),
.B1(n_136),
.B2(n_286),
.Y(n_285)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_98),
.Y(n_286)
);

AOI22x1_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_115),
.B1(n_124),
.B2(n_125),
.Y(n_98)
);

AOI22x1_ASAP7_75t_L g253 ( 
.A1(n_99),
.A2(n_124),
.B1(n_125),
.B2(n_254),
.Y(n_253)
);

OA21x2_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_104),
.B(n_109),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_100),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_104),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_106),
.Y(n_242)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_109),
.B(n_225),
.C(n_226),
.Y(n_224)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_111),
.Y(n_270)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_116),
.Y(n_254)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_126),
.Y(n_228)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_160),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_137),
.B(n_160),
.Y(n_279)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

BUFx4f_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_200),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_197),
.B2(n_198),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_165),
.B(n_200),
.C(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_193),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_167),
.Y(n_314)
);

AOI21x1_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_171),
.B(n_181),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_178),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_190),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_217),
.B1(n_218),
.B2(n_220),
.Y(n_216)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_193),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_193),
.B(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_194),
.B(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_194),
.B(n_272),
.Y(n_273)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_195),
.Y(n_311)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_198),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_L g260 ( 
.A(n_199),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_199),
.B(n_261),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_222),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_203),
.Y(n_298)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B(n_211),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g316 ( 
.A1(n_204),
.A2(n_205),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_212),
.Y(n_318)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_215),
.Y(n_317)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_229),
.B1(n_230),
.B2(n_232),
.Y(n_222)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_223),
.B(n_230),
.C(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_229),
.A2(n_230),
.B1(n_252),
.B2(n_263),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_229),
.B(n_252),
.C(n_279),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_230),
.Y(n_229)
);

AOI21x1_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_282),
.B(n_287),
.Y(n_233)
);

OAI21x1_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_276),
.B(n_281),
.Y(n_234)
);

AOI21x1_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_259),
.B(n_275),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_255),
.Y(n_236)
);

NOR2xp67_ASAP7_75t_SL g275 ( 
.A(n_237),
.B(n_255),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_252),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_252),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_243),
.B(n_247),
.Y(n_238)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_252),
.A2(n_263),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI21x1_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_264),
.B(n_274),
.Y(n_259)
);

AOI21x1_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_271),
.B(n_273),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_284),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_319),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_294),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_294),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_312),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_299),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx12f_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);


endmodule