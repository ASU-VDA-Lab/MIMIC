module fake_aes_6930_n_941 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_941, n_945);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_941;
output n_945;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_925;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_232;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_476;
wire n_227;
wire n_384;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_769;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_939;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_910;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_926;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_208;
wire n_200;
wire n_573;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_899;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_924;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_916;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g113 ( .A(n_44), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_80), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_68), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_28), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_95), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_71), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_42), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_5), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_28), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_19), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_65), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_34), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_26), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_67), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_107), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_6), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_25), .Y(n_129) );
INVx1_ASAP7_75t_SL g130 ( .A(n_12), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_48), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_21), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_83), .Y(n_133) );
BUFx2_ASAP7_75t_SL g134 ( .A(n_22), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_79), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_76), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_54), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_70), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_22), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_45), .Y(n_140) );
BUFx10_ASAP7_75t_L g141 ( .A(n_23), .Y(n_141) );
CKINVDCx16_ASAP7_75t_R g142 ( .A(n_13), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_77), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_85), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_94), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_110), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_62), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_16), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_74), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_24), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_52), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_61), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_104), .Y(n_153) );
BUFx2_ASAP7_75t_SL g154 ( .A(n_109), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_4), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_13), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_73), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_120), .B(n_0), .Y(n_158) );
AND2x6_ASAP7_75t_L g159 ( .A(n_121), .B(n_0), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_121), .B(n_1), .Y(n_160) );
INVx5_ASAP7_75t_L g161 ( .A(n_113), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_115), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_121), .B(n_1), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_115), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_148), .B(n_2), .Y(n_165) );
BUFx12f_ASAP7_75t_L g166 ( .A(n_113), .Y(n_166) );
INVx5_ASAP7_75t_L g167 ( .A(n_113), .Y(n_167) );
INVx5_ASAP7_75t_L g168 ( .A(n_113), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_136), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_116), .B(n_2), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_148), .B(n_3), .Y(n_171) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_120), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_142), .B(n_3), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_148), .B(n_4), .Y(n_174) );
BUFx8_ASAP7_75t_SL g175 ( .A(n_118), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_142), .B(n_5), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_136), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_115), .B(n_6), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_116), .B(n_7), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_137), .B(n_7), .Y(n_180) );
BUFx12f_ASAP7_75t_L g181 ( .A(n_113), .Y(n_181) );
AND2x2_ASAP7_75t_SL g182 ( .A(n_180), .B(n_137), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_178), .Y(n_183) );
OAI22xp33_ASAP7_75t_SL g184 ( .A1(n_172), .A2(n_130), .B1(n_156), .B2(n_132), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_162), .Y(n_185) );
INVx2_ASAP7_75t_SL g186 ( .A(n_172), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_172), .B(n_141), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_173), .A2(n_129), .B1(n_128), .B2(n_124), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_173), .A2(n_150), .B1(n_125), .B2(n_139), .Y(n_189) );
OAI22xp33_ASAP7_75t_SL g190 ( .A1(n_170), .A2(n_130), .B1(n_139), .B2(n_149), .Y(n_190) );
CKINVDCx6p67_ASAP7_75t_R g191 ( .A(n_173), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_158), .B(n_141), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_180), .B(n_149), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_169), .B(n_114), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_173), .A2(n_140), .B1(n_151), .B2(n_126), .Y(n_195) );
CKINVDCx6p67_ASAP7_75t_R g196 ( .A(n_173), .Y(n_196) );
OAI22xp33_ASAP7_75t_SL g197 ( .A1(n_170), .A2(n_122), .B1(n_155), .B2(n_141), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_162), .Y(n_198) );
OAI22xp33_ASAP7_75t_L g199 ( .A1(n_170), .A2(n_157), .B1(n_153), .B2(n_152), .Y(n_199) );
OAI22xp33_ASAP7_75t_SL g200 ( .A1(n_179), .A2(n_141), .B1(n_119), .B2(n_123), .Y(n_200) );
OAI22xp5_ASAP7_75t_SL g201 ( .A1(n_179), .A2(n_134), .B1(n_154), .B2(n_146), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_176), .A2(n_134), .B1(n_154), .B2(n_145), .Y(n_202) );
OR2x2_ASAP7_75t_L g203 ( .A(n_158), .B(n_8), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_178), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_169), .B(n_117), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_176), .A2(n_147), .B1(n_144), .B2(n_143), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_178), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_158), .B(n_113), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_176), .A2(n_138), .B1(n_135), .B2(n_133), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_176), .A2(n_131), .B1(n_127), .B2(n_10), .Y(n_210) );
OAI22xp33_ASAP7_75t_L g211 ( .A1(n_179), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_158), .B(n_9), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_158), .B(n_11), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_166), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_178), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_178), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_178), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_176), .B(n_11), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_162), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_169), .B(n_12), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_169), .B(n_14), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_160), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_180), .A2(n_15), .B1(n_17), .B2(n_18), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_162), .Y(n_224) );
OAI22xp33_ASAP7_75t_L g225 ( .A1(n_177), .A2(n_17), .B1(n_18), .B2(n_19), .Y(n_225) );
AO22x2_ASAP7_75t_L g226 ( .A1(n_178), .A2(n_20), .B1(n_21), .B2(n_23), .Y(n_226) );
AO22x2_ASAP7_75t_L g227 ( .A1(n_178), .A2(n_20), .B1(n_24), .B2(n_25), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_178), .Y(n_228) );
OAI22xp33_ASAP7_75t_SL g229 ( .A1(n_160), .A2(n_26), .B1(n_27), .B2(n_29), .Y(n_229) );
INVx4_ASAP7_75t_L g230 ( .A(n_214), .Y(n_230) );
XOR2xp5_ASAP7_75t_L g231 ( .A(n_195), .B(n_175), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_186), .B(n_177), .Y(n_232) );
AOI21x1_ASAP7_75t_L g233 ( .A1(n_193), .A2(n_177), .B(n_180), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_220), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_212), .B(n_160), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_186), .B(n_177), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_192), .B(n_160), .Y(n_237) );
XOR2xp5_ASAP7_75t_L g238 ( .A(n_188), .B(n_175), .Y(n_238) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_193), .A2(n_180), .B(n_165), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_212), .B(n_160), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_220), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_221), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_221), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_192), .B(n_180), .Y(n_244) );
INVx4_ASAP7_75t_L g245 ( .A(n_214), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_203), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_191), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_206), .B(n_180), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_203), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_187), .B(n_180), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_208), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_212), .B(n_160), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_209), .B(n_180), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_208), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_208), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_183), .A2(n_165), .B(n_174), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_213), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_213), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_185), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_204), .A2(n_165), .B(n_174), .Y(n_260) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_191), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_185), .Y(n_262) );
XOR2xp5_ASAP7_75t_L g263 ( .A(n_210), .B(n_175), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_207), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_196), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_215), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_187), .B(n_160), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_196), .B(n_160), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_189), .B(n_160), .Y(n_269) );
INVxp33_ASAP7_75t_L g270 ( .A(n_218), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_198), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_216), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_217), .Y(n_273) );
XOR2xp5_ASAP7_75t_L g274 ( .A(n_197), .B(n_163), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_228), .A2(n_165), .B(n_174), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_218), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g277 ( .A(n_201), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_198), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_202), .B(n_163), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_223), .B(n_163), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_219), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_182), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_219), .Y(n_283) );
INVx2_ASAP7_75t_SL g284 ( .A(n_182), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_224), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_194), .B(n_163), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_222), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_200), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_224), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_184), .Y(n_290) );
INVxp33_ASAP7_75t_SL g291 ( .A(n_194), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_226), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_205), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_199), .B(n_163), .Y(n_294) );
INVx4_ASAP7_75t_SL g295 ( .A(n_226), .Y(n_295) );
AND2x2_ASAP7_75t_SL g296 ( .A(n_292), .B(n_163), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_262), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_268), .B(n_226), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_268), .B(n_226), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_264), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_284), .B(n_227), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_291), .B(n_190), .Y(n_302) );
INVxp67_ASAP7_75t_L g303 ( .A(n_235), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_266), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_262), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_295), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_272), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_284), .B(n_227), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_273), .Y(n_309) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_235), .B(n_163), .Y(n_310) );
INVxp67_ASAP7_75t_L g311 ( .A(n_235), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_295), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_247), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_256), .A2(n_229), .B(n_163), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_240), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_271), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_295), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_271), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_278), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_285), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_237), .B(n_227), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_240), .B(n_163), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_295), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_240), .B(n_165), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_237), .B(n_227), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_252), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_281), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_285), .Y(n_328) );
OR2x2_ASAP7_75t_SL g329 ( .A(n_269), .B(n_225), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_252), .B(n_165), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_293), .B(n_211), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_285), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_230), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_252), .B(n_165), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_230), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_230), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_283), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_289), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_251), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_285), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_280), .B(n_165), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_259), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_280), .B(n_165), .Y(n_343) );
OAI21xp5_ASAP7_75t_L g344 ( .A1(n_275), .A2(n_174), .B(n_171), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_259), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_259), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_280), .B(n_171), .Y(n_347) );
INVx4_ASAP7_75t_L g348 ( .A(n_245), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_245), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_247), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_326), .B(n_293), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_302), .B(n_291), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_341), .B(n_282), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_302), .B(n_270), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_300), .B(n_244), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_300), .B(n_267), .Y(n_356) );
OR2x6_ASAP7_75t_L g357 ( .A(n_306), .B(n_234), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_297), .Y(n_358) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_312), .Y(n_359) );
INVx4_ASAP7_75t_L g360 ( .A(n_306), .Y(n_360) );
NOR2xp33_ASAP7_75t_SL g361 ( .A(n_306), .B(n_261), .Y(n_361) );
NAND2x1p5_ASAP7_75t_L g362 ( .A(n_306), .B(n_241), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_297), .Y(n_363) );
INVxp67_ASAP7_75t_L g364 ( .A(n_349), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_300), .B(n_257), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_304), .B(n_258), .Y(n_366) );
AND2x2_ASAP7_75t_SL g367 ( .A(n_312), .B(n_248), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_304), .B(n_276), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_349), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_297), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_315), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_341), .B(n_270), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_326), .B(n_242), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_302), .B(n_246), .Y(n_374) );
INVx3_ASAP7_75t_L g375 ( .A(n_348), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_315), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_297), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_297), .Y(n_378) );
NAND2x1p5_ASAP7_75t_L g379 ( .A(n_348), .B(n_243), .Y(n_379) );
INVx6_ASAP7_75t_L g380 ( .A(n_348), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_326), .B(n_260), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_304), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_326), .B(n_254), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_326), .B(n_255), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_359), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_380), .Y(n_386) );
INVx1_ASAP7_75t_SL g387 ( .A(n_358), .Y(n_387) );
INVxp67_ASAP7_75t_SL g388 ( .A(n_358), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_360), .Y(n_389) );
INVx1_ASAP7_75t_SL g390 ( .A(n_358), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_358), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_359), .Y(n_392) );
BUFx12f_ASAP7_75t_L g393 ( .A(n_360), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_360), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_363), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_363), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_363), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_363), .Y(n_398) );
BUFx3_ASAP7_75t_L g399 ( .A(n_380), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_370), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_360), .Y(n_401) );
INVx6_ASAP7_75t_SL g402 ( .A(n_357), .Y(n_402) );
BUFx12f_ASAP7_75t_L g403 ( .A(n_360), .Y(n_403) );
BUFx12f_ASAP7_75t_L g404 ( .A(n_360), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_382), .B(n_381), .Y(n_405) );
INVx5_ASAP7_75t_L g406 ( .A(n_380), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_380), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_370), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_375), .B(n_319), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_380), .Y(n_410) );
BUFx12f_ASAP7_75t_L g411 ( .A(n_380), .Y(n_411) );
BUFx3_ASAP7_75t_L g412 ( .A(n_380), .Y(n_412) );
BUFx12f_ASAP7_75t_L g413 ( .A(n_379), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_379), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g415 ( .A1(n_413), .A2(n_361), .B1(n_379), .B2(n_357), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_396), .Y(n_416) );
INVx2_ASAP7_75t_SL g417 ( .A(n_413), .Y(n_417) );
INVx6_ASAP7_75t_L g418 ( .A(n_413), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_389), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_388), .A2(n_377), .B(n_370), .Y(n_420) );
INVx6_ASAP7_75t_L g421 ( .A(n_413), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_396), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_413), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_393), .A2(n_352), .B1(n_374), .B2(n_287), .Y(n_424) );
INVx6_ASAP7_75t_L g425 ( .A(n_393), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_393), .A2(n_352), .B1(n_374), .B2(n_287), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_396), .Y(n_427) );
BUFx2_ASAP7_75t_L g428 ( .A(n_385), .Y(n_428) );
INVx6_ASAP7_75t_L g429 ( .A(n_393), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g430 ( .A1(n_393), .A2(n_361), .B1(n_261), .B2(n_265), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_391), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_396), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_397), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_397), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_389), .A2(n_367), .B1(n_357), .B2(n_379), .Y(n_435) );
BUFx3_ASAP7_75t_L g436 ( .A(n_403), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_397), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_391), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_397), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_403), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_403), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_410), .Y(n_442) );
CKINVDCx6p67_ASAP7_75t_R g443 ( .A(n_403), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_403), .A2(n_354), .B1(n_367), .B2(n_274), .Y(n_444) );
BUFx10_ASAP7_75t_L g445 ( .A(n_409), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_404), .A2(n_354), .B1(n_367), .B2(n_298), .Y(n_446) );
OAI21xp5_ASAP7_75t_SL g447 ( .A1(n_394), .A2(n_231), .B(n_238), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_404), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_404), .A2(n_367), .B1(n_298), .B2(n_299), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_385), .A2(n_357), .B1(n_379), .B2(n_265), .Y(n_450) );
INVx4_ASAP7_75t_L g451 ( .A(n_404), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_400), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_404), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_414), .A2(n_298), .B1(n_299), .B2(n_290), .Y(n_454) );
INVx8_ASAP7_75t_L g455 ( .A(n_411), .Y(n_455) );
BUFx8_ASAP7_75t_L g456 ( .A(n_414), .Y(n_456) );
NAND2x1p5_ASAP7_75t_L g457 ( .A(n_414), .B(n_375), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_414), .A2(n_298), .B1(n_299), .B2(n_290), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_400), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_431), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_419), .B(n_400), .Y(n_461) );
OAI22xp33_ASAP7_75t_L g462 ( .A1(n_423), .A2(n_414), .B1(n_394), .B2(n_401), .Y(n_462) );
INVx5_ASAP7_75t_L g463 ( .A(n_418), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_416), .Y(n_464) );
BUFx4f_ASAP7_75t_SL g465 ( .A(n_419), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_428), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_431), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_435), .A2(n_394), .B1(n_401), .B2(n_392), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_424), .A2(n_402), .B1(n_394), .B2(n_401), .Y(n_469) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_418), .A2(n_401), .B1(n_410), .B2(n_385), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_423), .A2(n_392), .B1(n_385), .B2(n_402), .Y(n_471) );
CKINVDCx11_ASAP7_75t_R g472 ( .A(n_442), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_438), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_430), .A2(n_392), .B1(n_402), .B2(n_357), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_438), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_422), .Y(n_476) );
INVxp67_ASAP7_75t_L g477 ( .A(n_417), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_427), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_432), .Y(n_479) );
AOI222xp33_ASAP7_75t_L g480 ( .A1(n_447), .A2(n_249), .B1(n_350), .B2(n_288), .C1(n_341), .C2(n_343), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_426), .A2(n_402), .B1(n_299), .B2(n_325), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_456), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_433), .B(n_400), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_443), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_434), .B(n_408), .Y(n_485) );
OAI22xp5_ASAP7_75t_SL g486 ( .A1(n_442), .A2(n_313), .B1(n_263), .B2(n_350), .Y(n_486) );
OAI22xp5_ASAP7_75t_SL g487 ( .A1(n_453), .A2(n_313), .B1(n_350), .B2(n_277), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_428), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_443), .Y(n_489) );
AOI22xp33_ASAP7_75t_SL g490 ( .A1(n_418), .A2(n_392), .B1(n_411), .B2(n_406), .Y(n_490) );
BUFx2_ASAP7_75t_L g491 ( .A(n_456), .Y(n_491) );
INVx4_ASAP7_75t_SL g492 ( .A(n_418), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_453), .Y(n_493) );
INVx6_ASAP7_75t_L g494 ( .A(n_456), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_421), .A2(n_402), .B1(n_325), .B2(n_321), .Y(n_495) );
AOI22xp33_ASAP7_75t_SL g496 ( .A1(n_421), .A2(n_411), .B1(n_406), .B2(n_350), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_437), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_450), .A2(n_402), .B1(n_357), .B2(n_406), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_415), .A2(n_402), .B1(n_357), .B2(n_406), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_421), .A2(n_402), .B1(n_325), .B2(n_321), .Y(n_500) );
OAI21xp33_ASAP7_75t_L g501 ( .A1(n_444), .A2(n_288), .B(n_174), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_421), .A2(n_325), .B1(n_321), .B2(n_411), .Y(n_502) );
INVx5_ASAP7_75t_SL g503 ( .A(n_455), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_455), .A2(n_321), .B1(n_411), .B2(n_381), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_425), .A2(n_357), .B1(n_406), .B2(n_388), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_439), .Y(n_506) );
AOI22xp33_ASAP7_75t_SL g507 ( .A1(n_425), .A2(n_406), .B1(n_388), .B2(n_409), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_417), .A2(n_277), .B1(n_372), .B2(n_279), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_455), .A2(n_381), .B1(n_376), .B2(n_371), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_452), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_459), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_440), .B(n_408), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_436), .Y(n_513) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_457), .Y(n_514) );
INVx4_ASAP7_75t_L g515 ( .A(n_451), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_420), .A2(n_331), .B(n_314), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_455), .A2(n_381), .B1(n_376), .B2(n_371), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_448), .B(n_408), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_436), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_454), .B(n_408), .Y(n_520) );
NOR2x1_ASAP7_75t_L g521 ( .A(n_451), .B(n_398), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_441), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_445), .B(n_387), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_441), .Y(n_524) );
BUFx3_ASAP7_75t_L g525 ( .A(n_425), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_445), .B(n_387), .Y(n_526) );
AOI22xp33_ASAP7_75t_SL g527 ( .A1(n_425), .A2(n_406), .B1(n_409), .B2(n_375), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_429), .A2(n_381), .B1(n_376), .B2(n_371), .Y(n_528) );
BUFx4f_ASAP7_75t_SL g529 ( .A(n_451), .Y(n_529) );
INVx1_ASAP7_75t_SL g530 ( .A(n_429), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_429), .A2(n_381), .B1(n_376), .B2(n_371), .Y(n_531) );
OAI21xp5_ASAP7_75t_SL g532 ( .A1(n_457), .A2(n_314), .B(n_362), .Y(n_532) );
AOI222xp33_ASAP7_75t_L g533 ( .A1(n_429), .A2(n_341), .B1(n_343), .B2(n_314), .C1(n_159), .C2(n_372), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_457), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_480), .A2(n_446), .B1(n_449), .B2(n_458), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_464), .Y(n_536) );
INVx2_ASAP7_75t_SL g537 ( .A(n_521), .Y(n_537) );
AOI22xp33_ASAP7_75t_SL g538 ( .A1(n_474), .A2(n_445), .B1(n_406), .B2(n_405), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_478), .B(n_405), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_470), .A2(n_406), .B1(n_329), .B2(n_405), .Y(n_540) );
AO22x1_ASAP7_75t_L g541 ( .A1(n_482), .A2(n_406), .B1(n_398), .B2(n_409), .Y(n_541) );
AOI222xp33_ASAP7_75t_L g542 ( .A1(n_501), .A2(n_159), .B1(n_171), .B2(n_174), .C1(n_343), .C2(n_301), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_479), .B(n_398), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_533), .A2(n_409), .B1(n_301), .B2(n_308), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_464), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_496), .A2(n_406), .B1(n_329), .B2(n_409), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_468), .A2(n_308), .B1(n_301), .B2(n_406), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_490), .A2(n_406), .B1(n_329), .B2(n_409), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_510), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_498), .A2(n_301), .B1(n_308), .B2(n_407), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_469), .A2(n_308), .B1(n_407), .B2(n_386), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_506), .B(n_387), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_510), .B(n_390), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_519), .B(n_390), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_461), .B(n_390), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_499), .A2(n_407), .B1(n_412), .B2(n_399), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_529), .A2(n_329), .B1(n_409), .B2(n_362), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_460), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_491), .A2(n_407), .B1(n_412), .B2(n_399), .Y(n_559) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_514), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_503), .A2(n_362), .B1(n_382), .B2(n_391), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_491), .A2(n_407), .B1(n_412), .B2(n_399), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_481), .A2(n_407), .B1(n_412), .B2(n_399), .Y(n_563) );
OAI211xp5_ASAP7_75t_SL g564 ( .A1(n_472), .A2(n_269), .B(n_164), .C(n_162), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_482), .A2(n_407), .B1(n_412), .B2(n_399), .Y(n_565) );
NOR3xp33_ASAP7_75t_L g566 ( .A(n_486), .B(n_331), .C(n_164), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_460), .Y(n_567) );
OAI221xp5_ASAP7_75t_L g568 ( .A1(n_508), .A2(n_253), .B1(n_347), .B2(n_365), .C(n_366), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_482), .A2(n_386), .B1(n_375), .B2(n_159), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_503), .A2(n_362), .B1(n_382), .B2(n_391), .Y(n_570) );
OAI221xp5_ASAP7_75t_L g571 ( .A1(n_532), .A2(n_347), .B1(n_365), .B2(n_366), .C(n_368), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_471), .A2(n_494), .B1(n_505), .B2(n_504), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_494), .A2(n_375), .B1(n_386), .B2(n_391), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_494), .A2(n_386), .B1(n_375), .B2(n_159), .Y(n_574) );
OAI222xp33_ASAP7_75t_L g575 ( .A1(n_515), .A2(n_362), .B1(n_395), .B2(n_369), .C1(n_364), .C2(n_386), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_503), .A2(n_395), .B1(n_364), .B2(n_369), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_503), .A2(n_395), .B1(n_368), .B2(n_370), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_494), .A2(n_351), .B1(n_372), .B2(n_356), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_515), .A2(n_395), .B1(n_343), .B2(n_317), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_476), .B(n_395), .Y(n_580) );
AOI22xp33_ASAP7_75t_SL g581 ( .A1(n_515), .A2(n_312), .B1(n_317), .B2(n_323), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_476), .B(n_377), .Y(n_582) );
OAI222xp33_ASAP7_75t_L g583 ( .A1(n_507), .A2(n_171), .B1(n_174), .B2(n_377), .C1(n_378), .C2(n_347), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_465), .A2(n_159), .B1(n_372), .B2(n_174), .Y(n_584) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_463), .A2(n_323), .B1(n_317), .B2(n_159), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_495), .A2(n_159), .B1(n_174), .B2(n_171), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_500), .A2(n_159), .B1(n_171), .B2(n_296), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_497), .B(n_511), .Y(n_588) );
OAI222xp33_ASAP7_75t_L g589 ( .A1(n_477), .A2(n_171), .B1(n_377), .B2(n_378), .C1(n_310), .C2(n_164), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_497), .B(n_159), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_527), .A2(n_378), .B1(n_323), .B2(n_356), .Y(n_591) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_463), .A2(n_159), .B1(n_171), .B2(n_378), .Y(n_592) );
OAI221xp5_ASAP7_75t_SL g593 ( .A1(n_502), .A2(n_355), .B1(n_294), .B2(n_164), .C(n_162), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_484), .A2(n_351), .B1(n_307), .B2(n_309), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_472), .B(n_27), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_462), .A2(n_159), .B1(n_171), .B2(n_296), .Y(n_596) );
OAI222xp33_ASAP7_75t_L g597 ( .A1(n_484), .A2(n_310), .B1(n_162), .B2(n_164), .C1(n_348), .C2(n_355), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_525), .A2(n_159), .B1(n_296), .B2(n_351), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_514), .B(n_463), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_511), .B(n_159), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_467), .B(n_162), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_525), .A2(n_159), .B1(n_296), .B2(n_351), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_467), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_513), .A2(n_159), .B1(n_296), .B2(n_351), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_522), .A2(n_524), .B1(n_520), .B2(n_528), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_512), .A2(n_159), .B(n_164), .Y(n_606) );
OAI222xp33_ASAP7_75t_L g607 ( .A1(n_489), .A2(n_310), .B1(n_164), .B2(n_348), .C1(n_327), .C2(n_337), .Y(n_607) );
AOI22xp33_ASAP7_75t_SL g608 ( .A1(n_463), .A2(n_159), .B1(n_351), .B2(n_348), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_531), .A2(n_307), .B1(n_309), .B2(n_373), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_518), .B(n_164), .Y(n_610) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_463), .A2(n_348), .B1(n_324), .B2(n_373), .Y(n_611) );
OAI222xp33_ASAP7_75t_L g612 ( .A1(n_489), .A2(n_310), .B1(n_337), .B2(n_338), .C1(n_319), .C2(n_327), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_509), .A2(n_337), .B1(n_338), .B2(n_327), .Y(n_613) );
BUFx12f_ASAP7_75t_L g614 ( .A(n_493), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_517), .A2(n_307), .B1(n_309), .B2(n_373), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_534), .A2(n_338), .B1(n_319), .B2(n_310), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_483), .B(n_29), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_534), .A2(n_310), .B1(n_373), .B2(n_316), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_493), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_466), .A2(n_373), .B1(n_353), .B2(n_286), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_488), .A2(n_373), .B1(n_353), .B2(n_286), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_530), .A2(n_316), .B1(n_318), .B2(n_305), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_523), .A2(n_316), .B1(n_318), .B2(n_305), .Y(n_623) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_514), .A2(n_324), .B1(n_353), .B2(n_344), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_487), .A2(n_324), .B1(n_344), .B2(n_250), .C(n_239), .Y(n_625) );
AOI22xp33_ASAP7_75t_SL g626 ( .A1(n_514), .A2(n_324), .B1(n_344), .B2(n_349), .Y(n_626) );
OAI222xp33_ASAP7_75t_L g627 ( .A1(n_523), .A2(n_318), .B1(n_324), .B2(n_334), .C1(n_322), .C2(n_330), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_526), .A2(n_384), .B1(n_383), .B2(n_324), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_485), .B(n_30), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_473), .B(n_161), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_492), .A2(n_384), .B1(n_383), .B2(n_232), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_526), .A2(n_384), .B1(n_383), .B2(n_324), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_516), .A2(n_384), .B1(n_383), .B2(n_315), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_514), .A2(n_384), .B1(n_383), .B2(n_315), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_492), .A2(n_384), .B1(n_383), .B2(n_315), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_473), .A2(n_305), .B1(n_333), .B2(n_336), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_475), .Y(n_637) );
NAND2xp33_ASAP7_75t_SL g638 ( .A(n_561), .B(n_492), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_536), .B(n_545), .Y(n_639) );
OAI21xp5_ASAP7_75t_SL g640 ( .A1(n_538), .A2(n_492), .B(n_475), .Y(n_640) );
OA21x2_ASAP7_75t_L g641 ( .A1(n_572), .A2(n_346), .B(n_345), .Y(n_641) );
OAI21xp5_ASAP7_75t_SL g642 ( .A1(n_575), .A2(n_236), .B(n_322), .Y(n_642) );
NOR2xp33_ASAP7_75t_R g643 ( .A(n_619), .B(n_30), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_536), .B(n_31), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_545), .B(n_161), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_549), .B(n_31), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g647 ( .A1(n_595), .A2(n_334), .B1(n_322), .B2(n_330), .C(n_339), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_549), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_571), .A2(n_339), .B1(n_333), .B2(n_335), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_605), .B(n_32), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_588), .B(n_32), .Y(n_651) );
NOR2xp33_ASAP7_75t_SL g652 ( .A(n_614), .B(n_305), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g653 ( .A(n_537), .B(n_161), .C(n_167), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_539), .B(n_33), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_619), .B(n_33), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_582), .B(n_34), .Y(n_656) );
OAI21xp5_ASAP7_75t_SL g657 ( .A1(n_611), .A2(n_334), .B(n_330), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_582), .B(n_35), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_601), .B(n_35), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_601), .B(n_36), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_603), .B(n_161), .Y(n_661) );
NAND4xp25_ASAP7_75t_L g662 ( .A(n_535), .B(n_36), .C(n_37), .D(n_38), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_603), .B(n_161), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_630), .B(n_37), .Y(n_664) );
NAND4xp25_ASAP7_75t_L g665 ( .A(n_557), .B(n_38), .C(n_39), .D(n_40), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_630), .B(n_39), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_637), .B(n_161), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g668 ( .A(n_537), .B(n_161), .C(n_167), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_637), .B(n_161), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_543), .B(n_40), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g671 ( .A(n_626), .B(n_570), .C(n_617), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_555), .B(n_161), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_541), .A2(n_305), .B(n_320), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_579), .A2(n_333), .B1(n_335), .B2(n_336), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_558), .B(n_161), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_567), .B(n_161), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_567), .B(n_161), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_560), .B(n_161), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g679 ( .A(n_629), .B(n_167), .C(n_168), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_546), .A2(n_339), .B1(n_333), .B2(n_335), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_610), .B(n_167), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_552), .B(n_167), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_553), .B(n_167), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_560), .B(n_167), .Y(n_684) );
NOR2xp33_ASAP7_75t_SL g685 ( .A(n_614), .B(n_320), .Y(n_685) );
OA21x2_ASAP7_75t_L g686 ( .A1(n_556), .A2(n_346), .B(n_345), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_554), .B(n_167), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_560), .B(n_167), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_560), .B(n_167), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_577), .B(n_167), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_560), .B(n_167), .Y(n_691) );
NOR2xp67_ASAP7_75t_L g692 ( .A(n_599), .B(n_167), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_580), .B(n_167), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_548), .B(n_168), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_550), .B(n_168), .Y(n_695) );
OAI221xp5_ASAP7_75t_L g696 ( .A1(n_566), .A2(n_311), .B1(n_303), .B2(n_168), .C(n_335), .Y(n_696) );
OAI221xp5_ASAP7_75t_SL g697 ( .A1(n_544), .A2(n_303), .B1(n_311), .B2(n_333), .C(n_335), .Y(n_697) );
OAI221xp5_ASAP7_75t_L g698 ( .A1(n_608), .A2(n_544), .B1(n_584), .B2(n_594), .C(n_624), .Y(n_698) );
NAND4xp25_ASAP7_75t_L g699 ( .A(n_569), .B(n_303), .C(n_311), .D(n_335), .Y(n_699) );
NAND3xp33_ASAP7_75t_SL g700 ( .A(n_573), .B(n_332), .C(n_320), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_540), .B(n_168), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_599), .B(n_168), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_590), .B(n_168), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_541), .B(n_168), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_600), .B(n_168), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_594), .A2(n_336), .B1(n_333), .B2(n_335), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_564), .A2(n_168), .B1(n_336), .B2(n_333), .C(n_259), .Y(n_707) );
OAI221xp5_ASAP7_75t_SL g708 ( .A1(n_574), .A2(n_336), .B1(n_320), .B2(n_340), .C(n_332), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_547), .B(n_168), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_578), .B(n_168), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_578), .B(n_168), .Y(n_711) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_576), .B(n_168), .C(n_345), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_633), .B(n_41), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_551), .B(n_43), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_625), .A2(n_336), .B1(n_345), .B2(n_342), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_616), .B(n_46), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g717 ( .A1(n_618), .A2(n_336), .B1(n_166), .B2(n_181), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_628), .B(n_632), .Y(n_718) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_606), .B(n_345), .C(n_342), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_623), .B(n_47), .Y(n_720) );
NAND3xp33_ASAP7_75t_L g721 ( .A(n_631), .B(n_342), .C(n_346), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_631), .B(n_49), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_620), .B(n_50), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_621), .B(n_51), .Y(n_724) );
OAI21xp5_ASAP7_75t_L g725 ( .A1(n_612), .A2(n_233), .B(n_328), .Y(n_725) );
OAI221xp5_ASAP7_75t_L g726 ( .A1(n_592), .A2(n_320), .B1(n_328), .B2(n_340), .C(n_332), .Y(n_726) );
OAI221xp5_ASAP7_75t_L g727 ( .A1(n_596), .A2(n_328), .B1(n_332), .B2(n_340), .C(n_342), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_607), .B(n_53), .Y(n_728) );
NOR3xp33_ASAP7_75t_SL g729 ( .A(n_597), .B(n_181), .C(n_166), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_559), .B(n_55), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_563), .B(n_56), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_562), .B(n_565), .Y(n_732) );
NAND3xp33_ASAP7_75t_L g733 ( .A(n_604), .B(n_342), .C(n_346), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_591), .B(n_57), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_615), .B(n_58), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_609), .B(n_59), .Y(n_736) );
OAI221xp5_ASAP7_75t_SL g737 ( .A1(n_598), .A2(n_340), .B1(n_332), .B2(n_328), .C(n_346), .Y(n_737) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_602), .B(n_340), .C(n_328), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_613), .B(n_60), .Y(n_739) );
OAI21xp33_ASAP7_75t_L g740 ( .A1(n_586), .A2(n_259), .B(n_64), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_636), .B(n_63), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_622), .B(n_181), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_635), .B(n_66), .Y(n_743) );
OR2x2_ASAP7_75t_L g744 ( .A(n_639), .B(n_634), .Y(n_744) );
INVxp67_ASAP7_75t_L g745 ( .A(n_638), .Y(n_745) );
NAND3xp33_ASAP7_75t_L g746 ( .A(n_671), .B(n_585), .C(n_542), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_639), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_678), .B(n_581), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_648), .B(n_568), .Y(n_749) );
NOR3xp33_ASAP7_75t_L g750 ( .A(n_662), .B(n_583), .C(n_593), .Y(n_750) );
OA211x2_ASAP7_75t_L g751 ( .A1(n_652), .A2(n_627), .B(n_587), .C(n_589), .Y(n_751) );
BUFx3_ASAP7_75t_L g752 ( .A(n_678), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g753 ( .A1(n_638), .A2(n_245), .B(n_72), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_684), .B(n_69), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_684), .B(n_75), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_698), .A2(n_181), .B1(n_166), .B2(n_82), .Y(n_756) );
OR2x2_ASAP7_75t_L g757 ( .A(n_677), .B(n_78), .Y(n_757) );
AND2x4_ASAP7_75t_L g758 ( .A(n_692), .B(n_81), .Y(n_758) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_650), .B(n_84), .C(n_86), .Y(n_759) );
INVx2_ASAP7_75t_SL g760 ( .A(n_643), .Y(n_760) );
OR2x2_ASAP7_75t_L g761 ( .A(n_645), .B(n_87), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_688), .B(n_88), .Y(n_762) );
OAI211xp5_ASAP7_75t_SL g763 ( .A1(n_655), .A2(n_89), .B(n_90), .C(n_91), .Y(n_763) );
OA211x2_ASAP7_75t_L g764 ( .A1(n_685), .A2(n_92), .B(n_93), .C(n_96), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_679), .B(n_97), .C(n_98), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_688), .B(n_99), .Y(n_766) );
NAND3xp33_ASAP7_75t_L g767 ( .A(n_653), .B(n_100), .C(n_101), .Y(n_767) );
NOR3xp33_ASAP7_75t_SL g768 ( .A(n_665), .B(n_181), .C(n_166), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_641), .B(n_102), .Y(n_769) );
NAND3xp33_ASAP7_75t_L g770 ( .A(n_668), .B(n_103), .C(n_105), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_732), .A2(n_718), .B1(n_647), .B2(n_640), .Y(n_771) );
NAND4xp75_ASAP7_75t_L g772 ( .A(n_641), .B(n_106), .C(n_108), .D(n_111), .Y(n_772) );
BUFx2_ASAP7_75t_L g773 ( .A(n_643), .Y(n_773) );
OR2x2_ASAP7_75t_SL g774 ( .A(n_641), .B(n_112), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_718), .A2(n_166), .B1(n_181), .B2(n_649), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_689), .B(n_691), .Y(n_776) );
NAND4xp25_ASAP7_75t_L g777 ( .A(n_697), .B(n_680), .C(n_715), .D(n_699), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_645), .B(n_644), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_689), .B(n_691), .Y(n_779) );
AOI221xp5_ASAP7_75t_L g780 ( .A1(n_654), .A2(n_670), .B1(n_651), .B2(n_657), .C(n_672), .Y(n_780) );
INVx3_ASAP7_75t_L g781 ( .A(n_686), .Y(n_781) );
OR2x2_ASAP7_75t_L g782 ( .A(n_675), .B(n_676), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_646), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_676), .B(n_661), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_663), .B(n_669), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_663), .B(n_669), .Y(n_786) );
AOI211xp5_ASAP7_75t_L g787 ( .A1(n_642), .A2(n_728), .B(n_674), .C(n_700), .Y(n_787) );
AO21x2_ASAP7_75t_L g788 ( .A1(n_687), .A2(n_683), .B(n_682), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g789 ( .A(n_659), .B(n_660), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_667), .B(n_693), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_686), .B(n_656), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_686), .B(n_702), .Y(n_792) );
AOI22xp33_ASAP7_75t_SL g793 ( .A1(n_722), .A2(n_712), .B1(n_721), .B2(n_714), .Y(n_793) );
AOI22xp33_ASAP7_75t_SL g794 ( .A1(n_714), .A2(n_713), .B1(n_731), .B2(n_696), .Y(n_794) );
AND2x2_ASAP7_75t_L g795 ( .A(n_703), .B(n_658), .Y(n_795) );
OR2x2_ASAP7_75t_L g796 ( .A(n_664), .B(n_666), .Y(n_796) );
NAND3xp33_ASAP7_75t_L g797 ( .A(n_717), .B(n_701), .C(n_694), .Y(n_797) );
NAND3xp33_ASAP7_75t_L g798 ( .A(n_694), .B(n_729), .C(n_742), .Y(n_798) );
OA211x2_ASAP7_75t_L g799 ( .A1(n_742), .A2(n_725), .B(n_740), .C(n_704), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_681), .B(n_705), .Y(n_800) );
OR2x2_ASAP7_75t_L g801 ( .A(n_690), .B(n_710), .Y(n_801) );
OA211x2_ASAP7_75t_L g802 ( .A1(n_716), .A2(n_734), .B(n_720), .C(n_730), .Y(n_802) );
AND2x4_ASAP7_75t_L g803 ( .A(n_703), .B(n_731), .Y(n_803) );
NOR3xp33_ASAP7_75t_L g804 ( .A(n_733), .B(n_738), .C(n_707), .Y(n_804) );
BUFx3_ASAP7_75t_L g805 ( .A(n_743), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_743), .B(n_741), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_711), .B(n_673), .Y(n_807) );
OR2x2_ASAP7_75t_L g808 ( .A(n_708), .B(n_737), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_723), .B(n_724), .Y(n_809) );
CKINVDCx8_ASAP7_75t_R g810 ( .A(n_726), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_735), .B(n_736), .Y(n_811) );
INVx3_ASAP7_75t_L g812 ( .A(n_741), .Y(n_812) );
OAI211xp5_ASAP7_75t_SL g813 ( .A1(n_739), .A2(n_727), .B(n_719), .C(n_706), .Y(n_813) );
OAI211xp5_ASAP7_75t_SL g814 ( .A1(n_713), .A2(n_480), .B(n_472), .C(n_595), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_695), .B(n_709), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_695), .A2(n_698), .B1(n_662), .B2(n_665), .Y(n_816) );
INVx1_ASAP7_75t_SL g817 ( .A(n_643), .Y(n_817) );
NOR3xp33_ASAP7_75t_L g818 ( .A(n_662), .B(n_595), .C(n_665), .Y(n_818) );
NAND3xp33_ASAP7_75t_L g819 ( .A(n_671), .B(n_650), .C(n_679), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_639), .B(n_648), .Y(n_820) );
OR2x2_ASAP7_75t_L g821 ( .A(n_639), .B(n_648), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_783), .B(n_747), .Y(n_822) );
XOR2x1_ASAP7_75t_L g823 ( .A(n_760), .B(n_799), .Y(n_823) );
XNOR2xp5_ASAP7_75t_L g824 ( .A(n_817), .B(n_773), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_820), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_771), .B(n_819), .Y(n_826) );
XNOR2xp5_ASAP7_75t_L g827 ( .A(n_751), .B(n_802), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_820), .B(n_821), .Y(n_828) );
XOR2x2_ASAP7_75t_L g829 ( .A(n_818), .B(n_746), .Y(n_829) );
XNOR2x2_ASAP7_75t_L g830 ( .A(n_753), .B(n_798), .Y(n_830) );
NAND4xp75_ASAP7_75t_SL g831 ( .A(n_792), .B(n_811), .C(n_809), .D(n_814), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_744), .Y(n_832) );
AND2x2_ASAP7_75t_L g833 ( .A(n_745), .B(n_812), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_749), .B(n_745), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_749), .B(n_778), .Y(n_835) );
XOR2x2_ASAP7_75t_L g836 ( .A(n_816), .B(n_750), .Y(n_836) );
BUFx2_ASAP7_75t_L g837 ( .A(n_752), .Y(n_837) );
NAND4xp25_ASAP7_75t_L g838 ( .A(n_787), .B(n_814), .C(n_780), .D(n_756), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_793), .A2(n_753), .B1(n_812), .B2(n_810), .Y(n_839) );
INVx2_ASAP7_75t_SL g840 ( .A(n_776), .Y(n_840) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_788), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_791), .B(n_781), .Y(n_842) );
OR2x2_ASAP7_75t_L g843 ( .A(n_785), .B(n_786), .Y(n_843) );
INVx2_ASAP7_75t_SL g844 ( .A(n_779), .Y(n_844) );
NAND4xp75_ASAP7_75t_L g845 ( .A(n_780), .B(n_764), .C(n_789), .D(n_768), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_795), .B(n_790), .Y(n_846) );
NAND4xp75_ASAP7_75t_L g847 ( .A(n_800), .B(n_748), .C(n_775), .D(n_807), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_788), .B(n_784), .Y(n_848) );
NAND2xp33_ASAP7_75t_R g849 ( .A(n_808), .B(n_758), .Y(n_849) );
INVxp67_ASAP7_75t_SL g850 ( .A(n_769), .Y(n_850) );
INVx3_ASAP7_75t_L g851 ( .A(n_805), .Y(n_851) );
INVx1_ASAP7_75t_SL g852 ( .A(n_754), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_785), .Y(n_853) );
INVx2_ASAP7_75t_SL g854 ( .A(n_782), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_786), .Y(n_855) );
NAND4xp25_ASAP7_75t_L g856 ( .A(n_797), .B(n_794), .C(n_793), .D(n_777), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_801), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_774), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_803), .B(n_806), .Y(n_859) );
NAND4xp75_ASAP7_75t_L g860 ( .A(n_807), .B(n_755), .C(n_766), .D(n_762), .Y(n_860) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_796), .Y(n_861) );
XNOR2xp5_ASAP7_75t_L g862 ( .A(n_794), .B(n_815), .Y(n_862) );
OR2x2_ASAP7_75t_L g863 ( .A(n_769), .B(n_815), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_804), .B(n_761), .Y(n_864) );
INVx6_ASAP7_75t_L g865 ( .A(n_758), .Y(n_865) );
XNOR2x2_ASAP7_75t_L g866 ( .A(n_772), .B(n_765), .Y(n_866) );
INVx1_ASAP7_75t_SL g867 ( .A(n_837), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_861), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_825), .Y(n_869) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_841), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_857), .Y(n_871) );
XOR2x2_ASAP7_75t_L g872 ( .A(n_836), .B(n_759), .Y(n_872) );
NOR2xp33_ASAP7_75t_L g873 ( .A(n_856), .B(n_823), .Y(n_873) );
XOR2x2_ASAP7_75t_L g874 ( .A(n_836), .B(n_767), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_848), .B(n_757), .Y(n_875) );
INVx1_ASAP7_75t_SL g876 ( .A(n_824), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_848), .B(n_770), .Y(n_877) );
XNOR2xp5_ASAP7_75t_L g878 ( .A(n_823), .B(n_813), .Y(n_878) );
BUFx2_ASAP7_75t_SL g879 ( .A(n_851), .Y(n_879) );
XNOR2x1_ASAP7_75t_L g880 ( .A(n_829), .B(n_763), .Y(n_880) );
XOR2x2_ASAP7_75t_L g881 ( .A(n_829), .B(n_763), .Y(n_881) );
XOR2x2_ASAP7_75t_L g882 ( .A(n_862), .B(n_813), .Y(n_882) );
XOR2x2_ASAP7_75t_L g883 ( .A(n_862), .B(n_827), .Y(n_883) );
INVxp67_ASAP7_75t_L g884 ( .A(n_826), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_857), .Y(n_885) );
INVxp67_ASAP7_75t_L g886 ( .A(n_826), .Y(n_886) );
OA22x2_ASAP7_75t_L g887 ( .A1(n_839), .A2(n_833), .B1(n_849), .B2(n_834), .Y(n_887) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_842), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_828), .Y(n_889) );
NOR2xp67_ASAP7_75t_L g890 ( .A(n_838), .B(n_851), .Y(n_890) );
XOR2x2_ASAP7_75t_L g891 ( .A(n_831), .B(n_830), .Y(n_891) );
AOI22xp5_ASAP7_75t_L g892 ( .A1(n_849), .A2(n_847), .B1(n_864), .B2(n_845), .Y(n_892) );
INVx2_ASAP7_75t_SL g893 ( .A(n_840), .Y(n_893) );
INVx1_ASAP7_75t_SL g894 ( .A(n_852), .Y(n_894) );
INVxp67_ASAP7_75t_L g895 ( .A(n_864), .Y(n_895) );
AOI22x1_ASAP7_75t_L g896 ( .A1(n_878), .A2(n_830), .B1(n_858), .B2(n_833), .Y(n_896) );
AOI22x1_ASAP7_75t_SL g897 ( .A1(n_876), .A2(n_858), .B1(n_832), .B2(n_851), .Y(n_897) );
BUFx2_ASAP7_75t_SL g898 ( .A(n_867), .Y(n_898) );
INVxp67_ASAP7_75t_L g899 ( .A(n_884), .Y(n_899) );
INVx2_ASAP7_75t_SL g900 ( .A(n_893), .Y(n_900) );
XOR2x2_ASAP7_75t_L g901 ( .A(n_883), .B(n_860), .Y(n_901) );
OA22x2_ASAP7_75t_L g902 ( .A1(n_892), .A2(n_835), .B1(n_842), .B2(n_854), .Y(n_902) );
BUFx4f_ASAP7_75t_SL g903 ( .A(n_894), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_868), .Y(n_904) );
XNOR2x1_ASAP7_75t_L g905 ( .A(n_891), .B(n_866), .Y(n_905) );
XOR2x2_ASAP7_75t_L g906 ( .A(n_882), .B(n_866), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_889), .Y(n_907) );
OAI22xp33_ASAP7_75t_L g908 ( .A1(n_887), .A2(n_865), .B1(n_863), .B2(n_850), .Y(n_908) );
INVxp67_ASAP7_75t_L g909 ( .A(n_884), .Y(n_909) );
INVx2_ASAP7_75t_L g910 ( .A(n_888), .Y(n_910) );
INVxp67_ASAP7_75t_L g911 ( .A(n_886), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_898), .Y(n_912) );
OAI322xp33_ASAP7_75t_L g913 ( .A1(n_902), .A2(n_886), .A3(n_873), .B1(n_895), .B2(n_887), .C1(n_880), .C2(n_877), .Y(n_913) );
INVx2_ASAP7_75t_SL g914 ( .A(n_903), .Y(n_914) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_911), .Y(n_915) );
OAI322xp33_ASAP7_75t_L g916 ( .A1(n_902), .A2(n_895), .A3(n_877), .B1(n_875), .B2(n_870), .C1(n_881), .C2(n_863), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_903), .Y(n_917) );
INVxp33_ASAP7_75t_L g918 ( .A(n_896), .Y(n_918) );
CKINVDCx16_ASAP7_75t_R g919 ( .A(n_897), .Y(n_919) );
OAI322xp33_ASAP7_75t_L g920 ( .A1(n_908), .A2(n_875), .A3(n_870), .B1(n_871), .B2(n_885), .C1(n_869), .C2(n_822), .Y(n_920) );
AOI221xp5_ASAP7_75t_L g921 ( .A1(n_913), .A2(n_908), .B1(n_899), .B2(n_909), .C(n_911), .Y(n_921) );
AOI22xp5_ASAP7_75t_L g922 ( .A1(n_919), .A2(n_890), .B1(n_906), .B2(n_905), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_912), .A2(n_909), .B1(n_899), .B2(n_900), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_915), .Y(n_924) );
INVxp67_ASAP7_75t_L g925 ( .A(n_917), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_922), .A2(n_918), .B1(n_912), .B2(n_914), .Y(n_926) );
INVxp67_ASAP7_75t_SL g927 ( .A(n_925), .Y(n_927) );
HB1xp67_ASAP7_75t_L g928 ( .A(n_924), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_927), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g930 ( .A1(n_926), .A2(n_914), .B1(n_923), .B2(n_918), .Y(n_930) );
NOR2x1_ASAP7_75t_L g931 ( .A(n_928), .B(n_916), .Y(n_931) );
INVx2_ASAP7_75t_L g932 ( .A(n_929), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_930), .Y(n_933) );
OAI211xp5_ASAP7_75t_L g934 ( .A1(n_933), .A2(n_921), .B(n_931), .C(n_901), .Y(n_934) );
CKINVDCx5p33_ASAP7_75t_R g935 ( .A(n_932), .Y(n_935) );
INVx2_ASAP7_75t_L g936 ( .A(n_935), .Y(n_936) );
INVx2_ASAP7_75t_L g937 ( .A(n_934), .Y(n_937) );
AO22x2_ASAP7_75t_L g938 ( .A1(n_937), .A2(n_932), .B1(n_904), .B2(n_910), .Y(n_938) );
INVxp67_ASAP7_75t_L g939 ( .A(n_938), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g940 ( .A1(n_939), .A2(n_936), .B1(n_872), .B2(n_874), .Y(n_940) );
UNKNOWN g941 ( );
AO22x1_ASAP7_75t_L g942 ( .A1(n_941), .A2(n_907), .B1(n_855), .B2(n_853), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_942), .Y(n_943) );
AOI221xp5_ASAP7_75t_L g944 ( .A1(n_943), .A2(n_920), .B1(n_879), .B2(n_840), .C(n_844), .Y(n_944) );
AOI211xp5_ASAP7_75t_L g945 ( .A1(n_944), .A2(n_843), .B(n_846), .C(n_859), .Y(n_945) );
endmodule