module real_aes_16721_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_792;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_0), .Y(n_548) );
AND2x4_ASAP7_75t_L g850 ( .A(n_1), .B(n_851), .Y(n_850) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_2), .A2(n_4), .B1(n_273), .B2(n_274), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_3), .A2(n_22), .B1(n_200), .B2(n_209), .Y(n_217) );
AOI22xp33_ASAP7_75t_L g157 ( .A1(n_5), .A2(n_53), .B1(n_158), .B2(n_159), .Y(n_157) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_6), .A2(n_104), .B1(n_847), .B2(n_857), .Y(n_103) );
BUFx3_ASAP7_75t_L g499 ( .A(n_7), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_8), .A2(n_14), .B1(n_130), .B2(n_132), .Y(n_129) );
INVx1_ASAP7_75t_L g851 ( .A(n_9), .Y(n_851) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_10), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_11), .B(n_183), .Y(n_505) );
OR2x2_ASAP7_75t_L g113 ( .A(n_12), .B(n_31), .Y(n_113) );
BUFx2_ASAP7_75t_L g856 ( .A(n_12), .Y(n_856) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_13), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_15), .B(n_165), .Y(n_523) );
XNOR2xp5_ASAP7_75t_L g823 ( .A(n_16), .B(n_824), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_17), .B(n_174), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_18), .A2(n_88), .B1(n_165), .B2(n_209), .Y(n_563) );
OAI21x1_ASAP7_75t_L g142 ( .A1(n_19), .A2(n_47), .B(n_143), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g836 ( .A1(n_20), .A2(n_837), .B(n_844), .Y(n_836) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_21), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_23), .B(n_200), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_24), .B(n_135), .Y(n_229) );
INVx4_ASAP7_75t_R g182 ( .A(n_25), .Y(n_182) );
AO32x2_ASAP7_75t_L g560 ( .A1(n_26), .A2(n_211), .A3(n_212), .B1(n_561), .B2(n_564), .Y(n_560) );
AO32x1_ASAP7_75t_L g582 ( .A1(n_26), .A2(n_211), .A3(n_212), .B1(n_561), .B2(n_564), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_27), .B(n_200), .Y(n_235) );
INVx1_ASAP7_75t_L g278 ( .A(n_28), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_SL g206 ( .A1(n_29), .A2(n_130), .B(n_134), .C(n_207), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_30), .A2(n_44), .B1(n_130), .B2(n_137), .Y(n_218) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_31), .Y(n_854) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_32), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_33), .A2(n_52), .B1(n_184), .B2(n_200), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_34), .A2(n_93), .B1(n_137), .B2(n_209), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_35), .B(n_507), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_36), .B(n_529), .Y(n_573) );
INVx1_ASAP7_75t_L g232 ( .A(n_37), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_38), .B(n_130), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_39), .A2(n_70), .B1(n_137), .B2(n_554), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_40), .Y(n_251) );
INVx2_ASAP7_75t_L g108 ( .A(n_41), .Y(n_108) );
BUFx3_ASAP7_75t_L g111 ( .A(n_42), .Y(n_111) );
INVx1_ASAP7_75t_L g835 ( .A(n_42), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_43), .B(n_575), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_45), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g136 ( .A1(n_46), .A2(n_87), .B1(n_130), .B2(n_137), .Y(n_136) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_48), .A2(n_50), .B1(n_827), .B2(n_828), .Y(n_826) );
INVx1_ASAP7_75t_L g828 ( .A(n_48), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_49), .Y(n_544) );
INVx1_ASAP7_75t_L g827 ( .A(n_50), .Y(n_827) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_51), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_54), .A2(n_81), .B1(n_167), .B2(n_529), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_55), .Y(n_148) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_56), .A2(n_115), .B1(n_116), .B2(n_821), .Y(n_114) );
INVx1_ASAP7_75t_L g821 ( .A(n_56), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_57), .A2(n_85), .B1(n_165), .B2(n_209), .Y(n_495) );
INVx1_ASAP7_75t_L g143 ( .A(n_58), .Y(n_143) );
AND2x4_ASAP7_75t_L g145 ( .A(n_59), .B(n_146), .Y(n_145) );
XNOR2xp5_ASAP7_75t_L g820 ( .A(n_60), .B(n_61), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_62), .A2(n_92), .B1(n_137), .B2(n_271), .Y(n_270) );
AO22x1_ASAP7_75t_L g163 ( .A1(n_63), .A2(n_76), .B1(n_164), .B2(n_166), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_64), .B(n_209), .Y(n_504) );
INVx1_ASAP7_75t_L g146 ( .A(n_65), .Y(n_146) );
AND2x2_ASAP7_75t_L g210 ( .A(n_66), .B(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_67), .B(n_211), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_68), .A2(n_155), .B(n_158), .C(n_547), .Y(n_546) );
NAND3xp33_ASAP7_75t_L g510 ( .A(n_69), .B(n_209), .C(n_509), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_71), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_72), .B(n_158), .Y(n_257) );
AND2x2_ASAP7_75t_L g549 ( .A(n_73), .B(n_188), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_74), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_75), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_77), .B(n_200), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_78), .A2(n_98), .B1(n_165), .B2(n_167), .Y(n_531) );
INVx2_ASAP7_75t_L g135 ( .A(n_79), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_80), .B(n_253), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_82), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_83), .B(n_211), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_84), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_86), .B(n_141), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_89), .B(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_90), .A2(n_102), .B1(n_137), .B2(n_184), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_91), .B(n_529), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_94), .B(n_211), .Y(n_248) );
INVx1_ASAP7_75t_L g484 ( .A(n_95), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_95), .B(n_834), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_96), .B(n_174), .Y(n_576) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_97), .A2(n_139), .B(n_158), .C(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g187 ( .A(n_99), .B(n_188), .Y(n_187) );
NAND2xp33_ASAP7_75t_L g256 ( .A(n_100), .B(n_183), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_101), .Y(n_518) );
AO21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_114), .B(n_822), .Y(n_104) );
BUFx6f_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x6_ASAP7_75t_SL g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g830 ( .A(n_108), .B(n_831), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_108), .B(n_841), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NOR2x1_ASAP7_75t_L g843 ( .A(n_111), .B(n_113), .Y(n_843) );
NOR3x1_ASAP7_75t_L g848 ( .A(n_111), .B(n_849), .C(n_852), .Y(n_848) );
AND2x6_ASAP7_75t_SL g832 ( .A(n_112), .B(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
XOR2x1_ASAP7_75t_L g116 ( .A(n_117), .B(n_820), .Y(n_116) );
AOI22x1_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_481), .B1(n_485), .B2(n_819), .Y(n_117) );
INVx2_ASAP7_75t_L g825 ( .A(n_118), .Y(n_825) );
NOR2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_395), .Y(n_118) );
NAND4xp75_ASAP7_75t_L g119 ( .A(n_120), .B(n_300), .C(n_342), .D(n_366), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI211xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_189), .B(n_237), .C(n_279), .Y(n_121) );
INVxp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g386 ( .A(n_124), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g480 ( .A(n_124), .B(n_417), .Y(n_480) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_150), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g295 ( .A(n_126), .B(n_247), .Y(n_295) );
AND2x2_ASAP7_75t_L g336 ( .A(n_126), .B(n_297), .Y(n_336) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g243 ( .A(n_127), .B(n_172), .Y(n_243) );
OR2x2_ASAP7_75t_L g261 ( .A(n_127), .B(n_172), .Y(n_261) );
INVx2_ASAP7_75t_L g287 ( .A(n_127), .Y(n_287) );
AND2x2_ASAP7_75t_L g317 ( .A(n_127), .B(n_247), .Y(n_317) );
AND2x2_ASAP7_75t_L g346 ( .A(n_127), .B(n_171), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_127), .B(n_298), .Y(n_382) );
AO31x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_140), .A3(n_144), .B(n_147), .Y(n_127) );
OAI22x1_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_133), .B1(n_136), .B2(n_138), .Y(n_128) );
INVx4_ASAP7_75t_L g132 ( .A(n_130), .Y(n_132) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_131), .Y(n_137) );
INVx1_ASAP7_75t_L g158 ( .A(n_131), .Y(n_158) );
INVx1_ASAP7_75t_L g160 ( .A(n_131), .Y(n_160) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_131), .Y(n_165) );
INVx1_ASAP7_75t_L g167 ( .A(n_131), .Y(n_167) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_131), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_131), .Y(n_184) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_131), .Y(n_200) );
INVx1_ASAP7_75t_L g202 ( .A(n_131), .Y(n_202) );
INVx2_ASAP7_75t_L g209 ( .A(n_131), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_132), .A2(n_251), .B(n_252), .C(n_253), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_133), .A2(n_154), .B1(n_217), .B2(n_218), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_133), .A2(n_138), .B1(n_270), .B2(n_272), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_133), .A2(n_134), .B1(n_495), .B2(n_496), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_133), .A2(n_528), .B1(n_530), .B2(n_531), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_133), .A2(n_154), .B1(n_553), .B2(n_555), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_133), .A2(n_573), .B(n_574), .Y(n_572) );
INVx6_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_134), .B(n_163), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_134), .A2(n_256), .B(n_257), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g299 ( .A1(n_134), .A2(n_153), .B(n_163), .C(n_169), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_134), .A2(n_504), .B(n_505), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_134), .A2(n_204), .B1(n_562), .B2(n_563), .Y(n_561) );
BUFx8_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g139 ( .A(n_135), .Y(n_139) );
INVx2_ASAP7_75t_L g156 ( .A(n_135), .Y(n_156) );
INVx1_ASAP7_75t_L g205 ( .A(n_135), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_137), .B(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g273 ( .A(n_137), .Y(n_273) );
INVx2_ASAP7_75t_L g507 ( .A(n_137), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_138), .B(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_SL g530 ( .A(n_139), .Y(n_530) );
INVx1_ASAP7_75t_L g545 ( .A(n_139), .Y(n_545) );
INVx2_ASAP7_75t_L g501 ( .A(n_140), .Y(n_501) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g149 ( .A(n_141), .Y(n_149) );
OAI21xp33_ASAP7_75t_L g169 ( .A1(n_141), .A2(n_161), .B(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g175 ( .A(n_141), .Y(n_175) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_142), .Y(n_212) );
INVx2_ASAP7_75t_L g186 ( .A(n_144), .Y(n_186) );
BUFx10_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g170 ( .A(n_145), .Y(n_170) );
BUFx10_ASAP7_75t_L g220 ( .A(n_145), .Y(n_220) );
INVx1_ASAP7_75t_L g276 ( .A(n_145), .Y(n_276) );
AO31x2_ASAP7_75t_L g551 ( .A1(n_145), .A2(n_526), .A3(n_552), .B(n_556), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
INVx2_ASAP7_75t_L g188 ( .A(n_149), .Y(n_188) );
BUFx2_ASAP7_75t_L g195 ( .A(n_149), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_149), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_149), .B(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_149), .B(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g359 ( .A(n_150), .B(n_288), .Y(n_359) );
INVx2_ASAP7_75t_L g454 ( .A(n_150), .Y(n_454) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_171), .Y(n_150) );
INVx2_ASAP7_75t_L g242 ( .A(n_151), .Y(n_242) );
AND2x4_ASAP7_75t_L g285 ( .A(n_151), .B(n_172), .Y(n_285) );
AOI21x1_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_162), .B(n_168), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OAI21x1_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_157), .B(n_161), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_154), .A2(n_234), .B(n_235), .Y(n_233) );
AOI21x1_ASAP7_75t_L g569 ( .A1(n_154), .A2(n_570), .B(n_571), .Y(n_569) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g254 ( .A(n_156), .Y(n_254) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_160), .B(n_179), .Y(n_178) );
INVxp67_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
INVx3_ASAP7_75t_L g575 ( .A(n_165), .Y(n_575) );
OAI21xp33_ASAP7_75t_SL g228 ( .A1(n_166), .A2(n_229), .B(n_230), .Y(n_228) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_167), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_170), .A2(n_197), .B(n_206), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_170), .A2(n_541), .B(n_546), .Y(n_540) );
AND2x2_ASAP7_75t_L g444 ( .A(n_171), .B(n_242), .Y(n_444) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g308 ( .A(n_172), .Y(n_308) );
AND2x2_ASAP7_75t_L g365 ( .A(n_172), .B(n_247), .Y(n_365) );
AND2x2_ASAP7_75t_L g380 ( .A(n_172), .B(n_288), .Y(n_380) );
AND2x2_ASAP7_75t_L g402 ( .A(n_172), .B(n_242), .Y(n_402) );
AO21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_176), .B(n_187), .Y(n_172) );
AOI21x1_ASAP7_75t_L g539 ( .A1(n_173), .A2(n_540), .B(n_549), .Y(n_539) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_180), .B(n_186), .Y(n_176) );
OAI22xp33_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B1(n_184), .B2(n_185), .Y(n_181) );
INVx2_ASAP7_75t_L g271 ( .A(n_183), .Y(n_271) );
INVx1_ASAP7_75t_L g522 ( .A(n_184), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_184), .A2(n_200), .B1(n_543), .B2(n_544), .Y(n_542) );
OAI211xp5_ASAP7_75t_SL g449 ( .A1(n_189), .A2(n_450), .B(n_452), .C(n_459), .Y(n_449) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_223), .Y(n_190) );
INVxp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
OR2x2_ASAP7_75t_L g436 ( .A(n_192), .B(n_372), .Y(n_436) );
OR2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_213), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_193), .B(n_225), .Y(n_335) );
INVxp67_ASAP7_75t_L g349 ( .A(n_193), .Y(n_349) );
AND2x2_ASAP7_75t_L g369 ( .A(n_193), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_193), .B(n_282), .Y(n_376) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g265 ( .A(n_194), .Y(n_265) );
AOI21x1_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_210), .Y(n_194) );
AO31x2_ASAP7_75t_L g268 ( .A1(n_195), .A2(n_269), .A3(n_275), .B(n_277), .Y(n_268) );
OAI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_201), .B(n_204), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
INVx2_ASAP7_75t_L g554 ( .A(n_200), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
INVx2_ASAP7_75t_L g274 ( .A(n_202), .Y(n_274) );
O2A1O1Ixp5_ASAP7_75t_L g517 ( .A1(n_204), .A2(n_274), .B(n_518), .C(n_519), .Y(n_517) );
BUFx4f_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_205), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g509 ( .A(n_205), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
INVx2_ASAP7_75t_SL g529 ( .A(n_209), .Y(n_529) );
INVx2_ASAP7_75t_L g219 ( .A(n_211), .Y(n_219) );
NOR2x1_ASAP7_75t_L g258 ( .A(n_211), .B(n_259), .Y(n_258) );
INVx4_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g236 ( .A(n_212), .B(n_220), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_212), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g515 ( .A(n_212), .Y(n_515) );
BUFx3_ASAP7_75t_L g526 ( .A(n_212), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_212), .B(n_557), .Y(n_556) );
INVx2_ASAP7_75t_SL g567 ( .A(n_212), .Y(n_567) );
OR2x2_ASAP7_75t_L g310 ( .A(n_213), .B(n_292), .Y(n_310) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g358 ( .A(n_214), .B(n_265), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_214), .B(n_268), .Y(n_364) );
INVx2_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g264 ( .A(n_215), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g333 ( .A(n_215), .B(n_268), .Y(n_333) );
BUFx2_ASAP7_75t_L g340 ( .A(n_215), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_215), .B(n_268), .Y(n_420) );
AO31x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_219), .A3(n_220), .B(n_221), .Y(n_215) );
AOI31xp67_ASAP7_75t_L g493 ( .A1(n_219), .A2(n_220), .A3(n_494), .B(n_497), .Y(n_493) );
INVx1_ASAP7_75t_L g259 ( .A(n_220), .Y(n_259) );
OAI21x1_ASAP7_75t_L g502 ( .A1(n_220), .A2(n_503), .B(n_506), .Y(n_502) );
OAI21x1_ASAP7_75t_L g516 ( .A1(n_220), .A2(n_517), .B(n_520), .Y(n_516) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x4_ASAP7_75t_L g350 ( .A(n_224), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g479 ( .A(n_224), .B(n_264), .Y(n_479) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx3_ASAP7_75t_L g282 ( .A(n_225), .Y(n_282) );
AND2x2_ASAP7_75t_L g293 ( .A(n_225), .B(n_268), .Y(n_293) );
AND2x2_ASAP7_75t_L g339 ( .A(n_225), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g372 ( .A(n_225), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_225), .B(n_283), .Y(n_389) );
AND2x2_ASAP7_75t_L g428 ( .A(n_225), .B(n_429), .Y(n_428) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_233), .B(n_236), .Y(n_227) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_244), .B(n_262), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_239), .A2(n_407), .B1(n_408), .B2(n_410), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_243), .Y(n_239) );
AND2x2_ASAP7_75t_L g404 ( .A(n_240), .B(n_295), .Y(n_404) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g319 ( .A(n_241), .Y(n_319) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g468 ( .A(n_242), .B(n_288), .Y(n_468) );
AND2x2_ASAP7_75t_L g432 ( .A(n_243), .B(n_327), .Y(n_432) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_260), .Y(n_244) );
OR2x2_ASAP7_75t_L g329 ( .A(n_245), .B(n_306), .Y(n_329) );
OR2x2_ASAP7_75t_L g441 ( .A(n_245), .B(n_261), .Y(n_441) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g304 ( .A(n_246), .Y(n_304) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g288 ( .A(n_247), .Y(n_288) );
BUFx3_ASAP7_75t_L g370 ( .A(n_247), .Y(n_370) );
NAND2x1p5_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
OAI21x1_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_255), .B(n_258), .Y(n_249) );
INVx2_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_254), .A2(n_521), .B1(n_522), .B2(n_523), .Y(n_520) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g438 ( .A(n_261), .B(n_297), .Y(n_438) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
AND2x2_ASAP7_75t_L g280 ( .A(n_264), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g321 ( .A(n_264), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g458 ( .A(n_264), .Y(n_458) );
INVx1_ASAP7_75t_L g477 ( .A(n_264), .Y(n_477) );
INVx2_ASAP7_75t_L g292 ( .A(n_265), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_265), .B(n_268), .Y(n_341) );
INVx1_ASAP7_75t_L g405 ( .A(n_266), .Y(n_405) );
BUFx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g466 ( .A(n_267), .Y(n_466) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g283 ( .A(n_268), .Y(n_283) );
INVx1_ASAP7_75t_L g373 ( .A(n_268), .Y(n_373) );
AO31x2_ASAP7_75t_L g525 ( .A1(n_275), .A2(n_526), .A3(n_527), .B(n_532), .Y(n_525) );
INVx2_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_SL g564 ( .A(n_276), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_284), .B1(n_289), .B2(n_294), .Y(n_279) );
AND2x4_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx2_ASAP7_75t_L g322 ( .A(n_282), .Y(n_322) );
AND2x2_ASAP7_75t_L g324 ( .A(n_282), .B(n_309), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_282), .B(n_292), .Y(n_384) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx3_ASAP7_75t_L g315 ( .A(n_285), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_285), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g409 ( .A(n_285), .B(n_393), .Y(n_409) );
INVx1_ASAP7_75t_L g313 ( .A(n_286), .Y(n_313) );
AOI222xp33_ASAP7_75t_L g323 ( .A1(n_286), .A2(n_324), .B1(n_325), .B2(n_330), .C1(n_336), .C2(n_337), .Y(n_323) );
OAI21xp33_ASAP7_75t_SL g353 ( .A1(n_286), .A2(n_354), .B(n_355), .Y(n_353) );
AND2x2_ASAP7_75t_L g377 ( .A(n_286), .B(n_296), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_286), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
OR2x2_ASAP7_75t_L g306 ( .A(n_287), .B(n_298), .Y(n_306) );
INVx1_ASAP7_75t_L g394 ( .A(n_287), .Y(n_394) );
BUFx2_ASAP7_75t_L g328 ( .A(n_288), .Y(n_328) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_291), .B(n_332), .Y(n_361) );
OR2x2_ASAP7_75t_L g473 ( .A(n_291), .B(n_333), .Y(n_473) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g356 ( .A(n_293), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g471 ( .A(n_293), .Y(n_471) );
OAI31xp33_ASAP7_75t_L g452 ( .A1(n_294), .A2(n_453), .A3(n_455), .B(n_456), .Y(n_452) );
AND2x4_ASAP7_75t_SL g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_295), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_323), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_309), .B(n_311), .Y(n_301) );
NOR2x1_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x6_ASAP7_75t_L g422 ( .A(n_304), .B(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g354 ( .A(n_307), .Y(n_354) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g445 ( .A(n_308), .B(n_382), .Y(n_445) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_310), .A2(n_399), .B1(n_401), .B2(n_403), .Y(n_398) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_310), .A2(n_371), .B(n_433), .C(n_460), .Y(n_459) );
AOI21xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_316), .B(n_320), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND4xp25_ASAP7_75t_L g412 ( .A(n_315), .B(n_413), .C(n_414), .D(n_416), .Y(n_412) );
NAND2x1_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_317), .B(n_319), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_317), .B(n_402), .Y(n_425) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g391 ( .A(n_322), .B(n_351), .Y(n_391) );
NAND2xp33_ASAP7_75t_L g325 ( .A(n_326), .B(n_329), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_329), .A2(n_473), .B1(n_474), .B2(n_476), .Y(n_472) );
AOI221x1_ASAP7_75t_L g411 ( .A1(n_330), .A2(n_412), .B1(n_418), .B2(n_421), .C(n_424), .Y(n_411) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g351 ( .A(n_333), .Y(n_351) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g363 ( .A(n_335), .B(n_364), .Y(n_363) );
NAND2x1p5_ASAP7_75t_L g426 ( .A(n_336), .B(n_417), .Y(n_426) );
O2A1O1Ixp5_ASAP7_75t_L g439 ( .A1(n_337), .A2(n_421), .B(n_440), .C(n_442), .Y(n_439) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
INVx2_ASAP7_75t_L g388 ( .A(n_340), .Y(n_388) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_352), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_347), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_344), .A2(n_362), .B1(n_432), .B2(n_433), .C(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g368 ( .A(n_346), .B(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_346), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g467 ( .A(n_346), .B(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVxp67_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
NAND2x1_ASAP7_75t_L g446 ( .A(n_349), .B(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g470 ( .A(n_349), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g410 ( .A(n_350), .Y(n_410) );
AOI222xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_356), .B1(n_359), .B2(n_360), .C1(n_362), .C2(n_365), .Y(n_352) );
INVx1_ASAP7_75t_L g437 ( .A(n_356), .Y(n_437) );
INVx1_ASAP7_75t_L g400 ( .A(n_357), .Y(n_400) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g434 ( .A(n_358), .Y(n_434) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g375 ( .A(n_364), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g429 ( .A(n_364), .Y(n_429) );
AND2x2_ASAP7_75t_L g392 ( .A(n_365), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_385), .Y(n_366) );
AOI222xp33_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_371), .B1(n_374), .B2(n_377), .C1(n_378), .C2(n_383), .Y(n_367) );
INVx3_ASAP7_75t_L g417 ( .A(n_370), .Y(n_417) );
BUFx2_ASAP7_75t_L g475 ( .A(n_370), .Y(n_475) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g447 ( .A(n_372), .Y(n_447) );
OR2x2_ASAP7_75t_L g457 ( .A(n_372), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx2_ASAP7_75t_SL g415 ( .A(n_380), .Y(n_415) );
AND2x2_ASAP7_75t_L g460 ( .A(n_381), .B(n_417), .Y(n_460) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_382), .Y(n_413) );
INVxp67_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g419 ( .A(n_384), .B(n_420), .Y(n_419) );
NOR2x1_ASAP7_75t_L g385 ( .A(n_386), .B(n_390), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
OR2x2_ASAP7_75t_L g476 ( .A(n_389), .B(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_L g407 ( .A(n_391), .Y(n_407) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g414 ( .A(n_394), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g464 ( .A(n_394), .Y(n_464) );
NAND4xp75_ASAP7_75t_L g395 ( .A(n_396), .B(n_430), .C(n_448), .D(n_461), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_411), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_405), .B(n_406), .Y(n_397) );
INVxp33_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_400), .B(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g423 ( .A(n_402), .Y(n_423) );
AND2x2_ASAP7_75t_L g463 ( .A(n_402), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g433 ( .A(n_405), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g451 ( .A(n_416), .Y(n_451) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI22xp33_ASAP7_75t_SL g442 ( .A1(n_419), .A2(n_443), .B1(n_445), .B2(n_446), .Y(n_442) );
INVx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI21xp33_ASAP7_75t_SL g424 ( .A1(n_425), .A2(n_426), .B(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g455 ( .A(n_426), .Y(n_455) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_439), .Y(n_430) );
AOI21xp5_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_437), .B(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_478), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_465), .B1(n_467), .B2(n_469), .C(n_472), .Y(n_462) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx4_ASAP7_75t_L g819 ( .A(n_481), .Y(n_819) );
BUFx12f_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g842 ( .A(n_483), .B(n_843), .Y(n_842) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx2_ASAP7_75t_L g852 ( .A(n_484), .Y(n_852) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_720), .Y(n_485) );
AND4x1_ASAP7_75t_L g486 ( .A(n_487), .B(n_642), .C(n_675), .D(n_706), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_609), .Y(n_487) );
OAI221xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_534), .B1(n_577), .B2(n_587), .C(n_596), .Y(n_488) );
AOI21xp33_ASAP7_75t_L g714 ( .A1(n_489), .A2(n_699), .B(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_512), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_500), .Y(n_491) );
INVx2_ASAP7_75t_L g595 ( .A(n_492), .Y(n_595) );
AND2x2_ASAP7_75t_L g605 ( .A(n_492), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g641 ( .A(n_492), .B(n_525), .Y(n_641) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g630 ( .A(n_493), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g616 ( .A(n_500), .B(n_606), .Y(n_616) );
OR2x2_ASAP7_75t_L g725 ( .A(n_500), .B(n_514), .Y(n_725) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B(n_511), .Y(n_500) );
OAI21x1_ASAP7_75t_L g594 ( .A1(n_501), .A2(n_502), .B(n_511), .Y(n_594) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B(n_510), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_512), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_525), .Y(n_513) );
INVx1_ASAP7_75t_L g590 ( .A(n_514), .Y(n_590) );
INVx2_ASAP7_75t_SL g667 ( .A(n_514), .Y(n_667) );
BUFx2_ASAP7_75t_L g697 ( .A(n_514), .Y(n_697) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_524), .Y(n_514) );
OA21x2_ASAP7_75t_L g606 ( .A1(n_515), .A2(n_516), .B(n_524), .Y(n_606) );
AND2x2_ASAP7_75t_L g589 ( .A(n_525), .B(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g608 ( .A(n_525), .Y(n_608) );
OR2x2_ASAP7_75t_L g628 ( .A(n_525), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g669 ( .A(n_525), .Y(n_669) );
INVx1_ASAP7_75t_L g680 ( .A(n_525), .Y(n_680) );
AND2x2_ASAP7_75t_L g687 ( .A(n_525), .B(n_629), .Y(n_687) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2x1p5_ASAP7_75t_L g535 ( .A(n_536), .B(n_558), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_537), .B(n_550), .Y(n_536) );
INVx1_ASAP7_75t_L g601 ( .A(n_537), .Y(n_601) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_538), .Y(n_613) );
INVx1_ASAP7_75t_L g622 ( .A(n_538), .Y(n_622) );
INVx1_ASAP7_75t_L g661 ( .A(n_538), .Y(n_661) );
AND2x2_ASAP7_75t_L g691 ( .A(n_538), .B(n_551), .Y(n_691) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g585 ( .A(n_539), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_542), .B(n_545), .Y(n_541) );
INVx1_ASAP7_75t_L g597 ( .A(n_550), .Y(n_597) );
AND2x4_ASAP7_75t_L g646 ( .A(n_550), .B(n_560), .Y(n_646) );
AND2x2_ASAP7_75t_L g656 ( .A(n_550), .B(n_585), .Y(n_656) );
INVx1_ASAP7_75t_L g717 ( .A(n_550), .Y(n_717) );
INVx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g603 ( .A(n_551), .B(n_582), .Y(n_603) );
AND2x2_ASAP7_75t_L g621 ( .A(n_551), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g637 ( .A(n_551), .B(n_582), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_551), .B(n_565), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_558), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_565), .Y(n_558) );
OR2x2_ASAP7_75t_L g763 ( .A(n_559), .B(n_565), .Y(n_763) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g710 ( .A(n_560), .Y(n_710) );
AND2x2_ASAP7_75t_L g735 ( .A(n_560), .B(n_565), .Y(n_735) );
OAI21x1_ASAP7_75t_L g568 ( .A1(n_564), .A2(n_569), .B(n_572), .Y(n_568) );
INVx3_ASAP7_75t_L g586 ( .A(n_565), .Y(n_586) );
AND2x2_ASAP7_75t_L g612 ( .A(n_565), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g634 ( .A(n_565), .Y(n_634) );
INVx1_ASAP7_75t_L g648 ( .A(n_565), .Y(n_648) );
INVx1_ASAP7_75t_L g658 ( .A(n_565), .Y(n_658) );
BUFx2_ASAP7_75t_L g753 ( .A(n_565), .Y(n_753) );
OR2x2_ASAP7_75t_L g781 ( .A(n_565), .B(n_585), .Y(n_781) );
INVxp67_ASAP7_75t_L g798 ( .A(n_565), .Y(n_798) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI21x1_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B(n_576), .Y(n_566) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_583), .Y(n_578) );
AND2x4_ASAP7_75t_L g611 ( .A(n_579), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_579), .B(n_691), .Y(n_772) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g599 ( .A(n_581), .B(n_586), .Y(n_599) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_581), .Y(n_623) );
INVx1_ASAP7_75t_L g747 ( .A(n_581), .Y(n_747) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g660 ( .A(n_582), .Y(n_660) );
AND2x2_ASAP7_75t_L g674 ( .A(n_583), .B(n_637), .Y(n_674) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx1_ASAP7_75t_L g636 ( .A(n_585), .Y(n_636) );
OR2x2_ASAP7_75t_L g694 ( .A(n_585), .B(n_660), .Y(n_694) );
INVx1_ASAP7_75t_L g757 ( .A(n_585), .Y(n_757) );
AND2x2_ASAP7_75t_L g700 ( .A(n_586), .B(n_646), .Y(n_700) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x4_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
AND2x2_ASAP7_75t_L g703 ( .A(n_589), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
AND2x2_ASAP7_75t_L g607 ( .A(n_592), .B(n_608), .Y(n_607) );
NAND2x1p5_ASAP7_75t_L g652 ( .A(n_592), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g626 ( .A(n_593), .Y(n_626) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g705 ( .A(n_594), .B(n_630), .Y(n_705) );
AND2x2_ASAP7_75t_L g668 ( .A(n_595), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g739 ( .A(n_595), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_600), .C(n_604), .Y(n_596) );
INVx1_ASAP7_75t_L g731 ( .A(n_598), .Y(n_731) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x4_ASAP7_75t_L g727 ( .A(n_599), .B(n_691), .Y(n_727) );
INVx1_ASAP7_75t_L g818 ( .A(n_599), .Y(n_818) );
INVx1_ASAP7_75t_L g783 ( .A(n_600), .Y(n_783) );
AND2x4_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
AND2x2_ASAP7_75t_L g816 ( .A(n_601), .B(n_735), .Y(n_816) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g633 ( .A(n_603), .B(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g788 ( .A(n_603), .B(n_753), .Y(n_788) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVxp67_ASAP7_75t_L g678 ( .A(n_605), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_605), .B(n_640), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_605), .B(n_607), .Y(n_770) );
INVx1_ASAP7_75t_L g653 ( .A(n_606), .Y(n_653) );
INVx2_ASAP7_75t_SL g618 ( .A(n_608), .Y(n_618) );
OR2x2_ASAP7_75t_L g647 ( .A(n_608), .B(n_648), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_614), .B1(n_619), .B2(n_624), .C(n_631), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NOR2xp33_ASAP7_75t_SL g655 ( .A(n_611), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g683 ( .A(n_613), .Y(n_683) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g740 ( .A(n_616), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_616), .B(n_618), .Y(n_778) );
OR2x2_ASAP7_75t_L g760 ( .A(n_617), .B(n_750), .Y(n_760) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g729 ( .A(n_618), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g776 ( .A(n_618), .B(n_705), .Y(n_776) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
AND2x2_ASAP7_75t_L g711 ( .A(n_621), .B(n_634), .Y(n_711) );
BUFx2_ASAP7_75t_L g737 ( .A(n_621), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_625), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g640 ( .A(n_626), .Y(n_640) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g713 ( .A(n_628), .Y(n_713) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_635), .B(n_638), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g690 ( .A(n_634), .Y(n_690) );
INVxp67_ASAP7_75t_SL g693 ( .A(n_634), .Y(n_693) );
OR2x2_ASAP7_75t_L g803 ( .A(n_634), .B(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g764 ( .A(n_635), .Y(n_764) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g672 ( .A(n_636), .Y(n_672) );
AND2x2_ASAP7_75t_L g799 ( .A(n_637), .B(n_672), .Y(n_799) );
INVx2_ASAP7_75t_SL g804 ( .A(n_637), .Y(n_804) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx2_ASAP7_75t_L g686 ( .A(n_640), .Y(n_686) );
AND2x4_ASAP7_75t_L g662 ( .A(n_641), .B(n_651), .Y(n_662) );
INVx2_ASAP7_75t_L g726 ( .A(n_641), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_641), .B(n_667), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_641), .B(n_697), .Y(n_813) );
AOI221x1_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_649), .B1(n_654), .B2(n_662), .C(n_663), .Y(n_642) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx2_ASAP7_75t_L g782 ( .A(n_645), .Y(n_782) );
AOI21xp33_ASAP7_75t_L g789 ( .A1(n_645), .A2(n_790), .B(n_792), .Y(n_789) );
INVx3_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g671 ( .A(n_646), .B(n_672), .Y(n_671) );
BUFx2_ASAP7_75t_L g702 ( .A(n_646), .Y(n_702) );
AND2x4_ASAP7_75t_L g756 ( .A(n_646), .B(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g716 ( .A(n_648), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI32xp33_ASAP7_75t_L g761 ( .A1(n_650), .A2(n_759), .A3(n_762), .B1(n_764), .B2(n_765), .Y(n_761) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_651), .B(n_668), .Y(n_784) );
AND2x2_ASAP7_75t_L g800 ( .A(n_651), .B(n_680), .Y(n_800) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_655), .B(n_657), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_656), .B(n_798), .Y(n_797) );
O2A1O1Ixp33_ASAP7_75t_L g732 ( .A1(n_657), .A2(n_733), .B(n_736), .C(n_738), .Y(n_732) );
NAND2x1p5_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g681 ( .A(n_659), .Y(n_681) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
OAI21xp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_670), .B(n_673), .Y(n_663) );
OAI21xp33_ASAP7_75t_L g698 ( .A1(n_664), .A2(n_699), .B(n_701), .Y(n_698) );
INVx2_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_667), .B(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_671), .A2(n_744), .B1(n_748), .B2(n_749), .Y(n_743) );
AND2x2_ASAP7_75t_L g810 ( .A(n_671), .B(n_798), .Y(n_810) );
NOR2xp33_ASAP7_75t_SL g675 ( .A(n_676), .B(n_698), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_681), .B1(n_682), .B2(n_684), .C(n_688), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g786 ( .A1(n_677), .A2(n_787), .B(n_788), .Y(n_786) );
OR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
AND2x2_ASAP7_75t_L g769 ( .A(n_683), .B(n_735), .Y(n_769) );
INVxp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
AOI31xp33_ASAP7_75t_L g706 ( .A1(n_686), .A2(n_707), .A3(n_712), .B(n_714), .Y(n_706) );
AND2x2_ASAP7_75t_L g806 ( .A(n_686), .B(n_713), .Y(n_806) );
AND2x2_ASAP7_75t_L g695 ( .A(n_687), .B(n_696), .Y(n_695) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_687), .Y(n_759) );
INVx1_ASAP7_75t_L g793 ( .A(n_687), .Y(n_793) );
OAI21xp33_ASAP7_75t_SL g688 ( .A1(n_689), .A2(n_692), .B(n_695), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
INVx2_ASAP7_75t_L g719 ( .A(n_691), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_691), .B(n_818), .Y(n_817) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_692), .A2(n_775), .B(n_777), .Y(n_774) );
NOR2x1p5_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
O2A1O1Ixp33_ASAP7_75t_L g715 ( .A1(n_694), .A2(n_709), .B(n_716), .C(n_718), .Y(n_715) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g728 ( .A(n_697), .B(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g748 ( .A(n_697), .B(n_704), .Y(n_748) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g730 ( .A(n_705), .Y(n_730) );
INVx1_ASAP7_75t_L g766 ( .A(n_705), .Y(n_766) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_711), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_711), .A2(n_728), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g787 ( .A(n_711), .Y(n_787) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NOR2x1_ASAP7_75t_L g720 ( .A(n_721), .B(n_773), .Y(n_720) );
NAND3xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_741), .C(n_751), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_727), .B1(n_728), .B2(n_731), .C(n_732), .Y(n_722) );
INVx3_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g795 ( .A1(n_729), .A2(n_796), .B1(n_799), .B2(n_800), .Y(n_795) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OR2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
OR2x2_ASAP7_75t_L g792 ( .A(n_740), .B(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OR2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
INVx1_ASAP7_75t_L g791 ( .A(n_746), .Y(n_791) );
INVx2_ASAP7_75t_L g771 ( .A(n_748), .Y(n_771) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AOI211xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_754), .B(n_761), .C(n_767), .Y(n_751) );
BUFx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
OAI21xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_758), .B(n_760), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OR2x2_ASAP7_75t_L g762 ( .A(n_757), .B(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g805 ( .A(n_762), .Y(n_805) );
OAI22xp33_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_770), .B1(n_771), .B2(n_772), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NAND4xp75_ASAP7_75t_L g773 ( .A(n_774), .B(n_785), .C(n_794), .D(n_807), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
OAI22xp33_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B1(n_783), .B2(n_784), .Y(n_777) );
NAND2x1_ASAP7_75t_SL g779 ( .A(n_780), .B(n_782), .Y(n_779) );
INVx3_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_786), .B(n_789), .Y(n_785) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
AND2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_801), .Y(n_794) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
OAI21xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_805), .B(n_806), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_810), .B1(n_811), .B2(n_814), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVxp67_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_817), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
OAI21xp5_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_829), .B(n_836), .Y(n_822) );
XNOR2x1_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g829 ( .A(n_830), .Y(n_829) );
INVx5_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx4_ASAP7_75t_L g845 ( .A(n_832), .Y(n_845) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
BUFx10_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
AND2x2_ASAP7_75t_SL g847 ( .A(n_848), .B(n_853), .Y(n_847) );
AND2x6_ASAP7_75t_L g858 ( .A(n_848), .B(n_853), .Y(n_858) );
INVx2_ASAP7_75t_SL g849 ( .A(n_850), .Y(n_849) );
NOR2x1p5_ASAP7_75t_L g853 ( .A(n_854), .B(n_855), .Y(n_853) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx4_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
endmodule