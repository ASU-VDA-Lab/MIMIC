module fake_jpeg_10088_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_53),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_61),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_18),
.B1(n_27),
.B2(n_20),
.Y(n_83)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_30),
.B1(n_32),
.B2(n_16),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_58),
.B1(n_68),
.B2(n_18),
.Y(n_91)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_30),
.B1(n_32),
.B2(n_16),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_35),
.B(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_29),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_17),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_35),
.B(n_19),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_69),
.B(n_25),
.C(n_33),
.Y(n_95)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_70),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_30),
.B1(n_18),
.B2(n_27),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_30),
.B(n_33),
.C(n_25),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_86),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

OR2x4_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_21),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_78),
.A2(n_46),
.B(n_63),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_81)
);

AO22x1_ASAP7_75t_SL g124 ( 
.A1(n_81),
.A2(n_68),
.B1(n_26),
.B2(n_24),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_18),
.B1(n_17),
.B2(n_22),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_82),
.A2(n_90),
.B1(n_92),
.B2(n_108),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_83),
.A2(n_91),
.B1(n_99),
.B2(n_100),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_61),
.Y(n_86)
);

CKINVDCx12_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_88),
.Y(n_127)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_96),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_18),
.B1(n_22),
.B2(n_36),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_49),
.A2(n_22),
.B1(n_36),
.B2(n_20),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_47),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_62),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_48),
.A2(n_19),
.B1(n_20),
.B2(n_27),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_98),
.B1(n_103),
.B2(n_71),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_49),
.A2(n_19),
.B1(n_33),
.B2(n_25),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_69),
.A2(n_42),
.B1(n_31),
.B2(n_28),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_64),
.A2(n_31),
.B1(n_28),
.B2(n_23),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_55),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_101),
.B(n_109),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_104),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_66),
.A2(n_28),
.B1(n_23),
.B2(n_31),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_60),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_105),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_31),
.B1(n_28),
.B2(n_23),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_71),
.B1(n_56),
.B2(n_67),
.Y(n_119)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_110),
.A2(n_123),
.B(n_84),
.Y(n_153)
);

NOR2x1_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_66),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_111),
.B(n_81),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_114),
.B(n_94),
.Y(n_160)
);

AOI22x1_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_66),
.B1(n_58),
.B2(n_21),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_116),
.A2(n_81),
.B1(n_85),
.B2(n_106),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_118),
.B(n_125),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_120),
.B1(n_124),
.B2(n_128),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_46),
.B1(n_60),
.B2(n_71),
.Y(n_120)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_91),
.A2(n_80),
.B1(n_96),
.B2(n_86),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_31),
.B1(n_28),
.B2(n_23),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_130),
.A2(n_108),
.B1(n_85),
.B2(n_93),
.Y(n_142)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_73),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_76),
.B(n_0),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_76),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_84),
.B(n_9),
.C(n_15),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_11),
.C(n_14),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g136 ( 
.A(n_80),
.B(n_21),
.C(n_24),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_100),
.C(n_83),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_139),
.B(n_155),
.Y(n_204)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_140),
.B(n_144),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_148),
.B1(n_171),
.B2(n_119),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_77),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_143),
.A2(n_170),
.B(n_139),
.Y(n_203)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_150),
.Y(n_173)
);

INVxp67_ASAP7_75t_SL g194 ( 
.A(n_147),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_104),
.B1(n_77),
.B2(n_99),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_101),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_161),
.Y(n_181)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_109),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_152),
.Y(n_202)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_162),
.B(n_9),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_158),
.C(n_163),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_114),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_160),
.B(n_164),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_157),
.A2(n_165),
.B1(n_113),
.B2(n_125),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_94),
.C(n_81),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_106),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_159),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_81),
.C(n_107),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_110),
.A2(n_24),
.B(n_1),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_116),
.A2(n_88),
.B1(n_75),
.B2(n_105),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_138),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_134),
.Y(n_185)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_168),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_0),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_124),
.A2(n_75),
.B1(n_23),
.B2(n_24),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_178),
.B1(n_184),
.B2(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_180),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_190),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_163),
.A2(n_118),
.B1(n_137),
.B2(n_130),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_179),
.Y(n_222)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_137),
.B1(n_117),
.B2(n_126),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_200),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_146),
.B1(n_165),
.B2(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_193),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_134),
.B(n_24),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_188),
.A2(n_203),
.B(n_161),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_149),
.B(n_24),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_195),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_171),
.A2(n_122),
.B1(n_115),
.B2(n_133),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_191),
.A2(n_196),
.B1(n_199),
.B2(n_4),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_143),
.B(n_1),
.Y(n_192)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_153),
.B(n_24),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_24),
.B1(n_73),
.B2(n_3),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_168),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_198),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_164),
.Y(n_198)
);

AO22x1_ASAP7_75t_SL g199 ( 
.A1(n_170),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_199),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_221),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_143),
.B(n_140),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_208),
.B(n_209),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_158),
.B(n_144),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_173),
.B(n_150),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_220),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_174),
.A2(n_145),
.B(n_154),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_211),
.A2(n_188),
.B(n_189),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_152),
.Y(n_214)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_155),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_226),
.C(n_231),
.Y(n_245)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_169),
.B(n_3),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_223),
.Y(n_254)
);

OA22x2_ASAP7_75t_L g217 ( 
.A1(n_199),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_217),
.A2(n_196),
.B1(n_185),
.B2(n_180),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_204),
.B(n_13),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_172),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_2),
.Y(n_224)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_4),
.C(n_5),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_227),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_204),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_229),
.A2(n_187),
.B1(n_203),
.B2(n_192),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_236),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_208),
.B(n_195),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_244),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_193),
.B1(n_177),
.B2(n_184),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_239),
.A2(n_246),
.B1(n_248),
.B2(n_212),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_241),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_227),
.A2(n_175),
.B1(n_183),
.B2(n_176),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_252),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_253),
.C(n_226),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_186),
.B1(n_178),
.B2(n_183),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_247),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_213),
.A2(n_197),
.B1(n_201),
.B2(n_194),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_211),
.B(n_190),
.CI(n_201),
.CON(n_250),
.SN(n_250)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_251),
.Y(n_267)
);

NOR3xp33_ASAP7_75t_SL g251 ( 
.A(n_207),
.B(n_179),
.C(n_13),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_13),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_232),
.A2(n_225),
.B(n_209),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_258),
.A2(n_270),
.B(n_272),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_261),
.C(n_268),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_228),
.Y(n_260)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_260),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_215),
.C(n_232),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_262),
.A2(n_264),
.B1(n_239),
.B2(n_236),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_246),
.A2(n_206),
.B1(n_218),
.B2(n_212),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_224),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_273),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_244),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_240),
.A2(n_206),
.B(n_216),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_219),
.C(n_221),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_237),
.C(n_234),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_233),
.A2(n_216),
.B(n_222),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_248),
.B(n_254),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_275),
.A2(n_284),
.B(n_270),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_210),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_280),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_281),
.C(n_283),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_278),
.B(n_279),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_254),
.B1(n_251),
.B2(n_229),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_235),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_250),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_219),
.C(n_250),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_263),
.A2(n_205),
.B1(n_217),
.B2(n_235),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_220),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_285),
.B(n_286),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_11),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_262),
.B1(n_257),
.B2(n_269),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_289),
.A2(n_274),
.B1(n_217),
.B2(n_6),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_272),
.Y(n_291)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_291),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_278),
.B(n_273),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_301),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_295),
.A2(n_297),
.B(n_299),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_275),
.A2(n_267),
.B(n_255),
.Y(n_296)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_287),
.A2(n_255),
.B(n_258),
.Y(n_297)
);

AOI21x1_ASAP7_75t_L g299 ( 
.A1(n_281),
.A2(n_268),
.B(n_266),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_282),
.A2(n_273),
.B(n_266),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_300),
.A2(n_4),
.B(n_5),
.Y(n_310)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_284),
.A2(n_217),
.B(n_259),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_283),
.B1(n_274),
.B2(n_217),
.Y(n_302)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_306),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_10),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_309),
.B(n_310),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_298),
.B(n_297),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_307),
.A2(n_295),
.B1(n_301),
.B2(n_292),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_314),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_311),
.A2(n_292),
.B1(n_7),
.B2(n_8),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_318),
.C(n_305),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_304),
.A2(n_6),
.B(n_7),
.Y(n_317)
);

NAND2x1_ASAP7_75t_SL g321 ( 
.A(n_317),
.B(n_6),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_6),
.C(n_8),
.Y(n_318)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_322),
.C(n_303),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_303),
.B1(n_314),
.B2(n_315),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_324),
.B(n_320),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_323),
.B(n_313),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_321),
.Y(n_327)
);


endmodule