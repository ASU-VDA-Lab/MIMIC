module fake_jpeg_29237_n_387 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_387);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_387;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_292;
wire n_213;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_31),
.B(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_48),
.B(n_56),
.Y(n_122)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_53),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_60),
.Y(n_97)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_29),
.B(n_0),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_14),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_14),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_65),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_33),
.B(n_11),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_33),
.B(n_11),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_71),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_29),
.B(n_0),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_73),
.B(n_23),
.C(n_40),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_11),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

HAxp5_ASAP7_75t_SL g73 ( 
.A(n_23),
.B(n_1),
.CON(n_73),
.SN(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_83),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_44),
.B1(n_17),
.B2(n_20),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_89),
.A2(n_94),
.B1(n_125),
.B2(n_80),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_43),
.B1(n_42),
.B2(n_44),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_90),
.A2(n_95),
.B1(n_106),
.B2(n_113),
.Y(n_139)
);

OR2x4_ASAP7_75t_L g162 ( 
.A(n_91),
.B(n_125),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_43),
.B1(n_17),
.B2(n_34),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_92),
.B(n_37),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_17),
.B1(n_20),
.B2(n_24),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_25),
.B1(n_36),
.B2(n_26),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_66),
.A2(n_26),
.B1(n_28),
.B2(n_36),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_63),
.A2(n_23),
.B1(n_20),
.B2(n_40),
.Y(n_113)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_56),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_118),
.A2(n_123),
.B1(n_1),
.B2(n_2),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_70),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_126),
.Y(n_145)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_64),
.A2(n_35),
.B1(n_32),
.B2(n_24),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_69),
.A2(n_20),
.B1(n_24),
.B2(n_19),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_50),
.B(n_32),
.Y(n_126)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_68),
.A2(n_79),
.B1(n_78),
.B2(n_76),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_82),
.B1(n_59),
.B2(n_51),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_53),
.B(n_20),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_133),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_54),
.B(n_10),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_57),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_134),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_101),
.A2(n_81),
.B1(n_75),
.B2(n_74),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_135),
.B(n_144),
.Y(n_195)
);

BUFx2_ASAP7_75t_SL g136 ( 
.A(n_99),
.Y(n_136)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_136),
.Y(n_186)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx11_ASAP7_75t_L g210 ( 
.A(n_137),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_88),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_138),
.B(n_152),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx13_ASAP7_75t_L g201 ( 
.A(n_141),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_80),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_142),
.B(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_87),
.A2(n_19),
.B1(n_37),
.B2(n_10),
.Y(n_144)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

CKINVDCx12_ASAP7_75t_R g151 ( 
.A(n_86),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_151),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_122),
.B(n_9),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_80),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_176),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_154),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_156),
.A2(n_159),
.B1(n_171),
.B2(n_132),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_157),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_97),
.B(n_7),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_165),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_89),
.A2(n_47),
.B1(n_55),
.B2(n_49),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_161),
.A2(n_100),
.B1(n_119),
.B2(n_127),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_113),
.Y(n_180)
);

CKINVDCx12_ASAP7_75t_R g163 ( 
.A(n_99),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_163),
.Y(n_207)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_85),
.Y(n_164)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_109),
.B(n_110),
.C(n_9),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_166),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_167),
.A2(n_119),
.B1(n_100),
.B2(n_116),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_168),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_84),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_134),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_173),
.A2(n_144),
.B(n_171),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_6),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_174),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_105),
.B(n_4),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_175),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_4),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_157),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_181),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_112),
.B(n_103),
.Y(n_184)
);

OA21x2_ASAP7_75t_L g235 ( 
.A1(n_184),
.A2(n_146),
.B(n_137),
.Y(n_235)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_194),
.A2(n_197),
.B1(n_173),
.B2(n_135),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_151),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_163),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_139),
.A2(n_132),
.B1(n_115),
.B2(n_129),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_200),
.A2(n_140),
.B1(n_160),
.B2(n_169),
.Y(n_239)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_148),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_98),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_211),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_204),
.A2(n_205),
.B1(n_159),
.B2(n_156),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_162),
.A2(n_116),
.B1(n_102),
.B2(n_108),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_153),
.B(n_96),
.C(n_103),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_206),
.B(n_168),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_143),
.B(n_112),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_211),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_228),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_145),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_223),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_177),
.Y(n_220)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_220),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_221),
.A2(n_224),
.B(n_240),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_138),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_139),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_226),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_149),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_189),
.B(n_142),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_227),
.B(n_234),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_207),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_229),
.A2(n_230),
.B1(n_197),
.B2(n_200),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_180),
.A2(n_157),
.B1(n_148),
.B2(n_150),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_150),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_231),
.A2(n_191),
.B(n_187),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_207),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_236),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_183),
.B(n_170),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_235),
.A2(n_184),
.B(n_195),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_183),
.B(n_169),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_195),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_238),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_182),
.B(n_199),
.Y(n_238)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_195),
.A2(n_155),
.B1(n_108),
.B2(n_140),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_181),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_177),
.B(n_155),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_242),
.B(n_245),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_243),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_202),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_244),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_191),
.B(n_154),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_216),
.Y(n_251)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_262),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_187),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_266),
.C(n_237),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_260),
.A2(n_224),
.B1(n_233),
.B2(n_239),
.Y(n_272)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_216),
.Y(n_261)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_218),
.Y(n_263)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_235),
.A2(n_192),
.B(n_188),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_217),
.B(n_185),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_179),
.C(n_178),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_218),
.Y(n_267)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_220),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_242),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_272),
.A2(n_257),
.B1(n_264),
.B2(n_269),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_229),
.B1(n_233),
.B2(n_225),
.Y(n_274)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_283),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_232),
.Y(n_279)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_246),
.A2(n_214),
.B1(n_230),
.B2(n_215),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_292),
.B1(n_260),
.B2(n_262),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_248),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_281),
.B(n_255),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_231),
.C(n_221),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_291),
.C(n_294),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_221),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_288),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_270),
.B(n_228),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_287),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_245),
.Y(n_286)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_286),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_250),
.B(n_238),
.Y(n_287)
);

AOI221xp5_ASAP7_75t_L g288 ( 
.A1(n_256),
.A2(n_227),
.B1(n_226),
.B2(n_215),
.C(n_234),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_223),
.C(n_236),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_246),
.A2(n_235),
.B1(n_220),
.B2(n_204),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_219),
.C(n_178),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_264),
.B(n_258),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_295),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_307),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_299),
.B(n_289),
.C(n_290),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_301),
.A2(n_304),
.B1(n_305),
.B2(n_313),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_254),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_311),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_272),
.A2(n_257),
.B1(n_254),
.B2(n_249),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_284),
.A2(n_249),
.B1(n_247),
.B2(n_248),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_291),
.B(n_247),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_265),
.B1(n_258),
.B2(n_253),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_314),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_276),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_309),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_277),
.B(n_282),
.Y(n_311)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_312),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_273),
.A2(n_269),
.B1(n_266),
.B2(n_253),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_284),
.A2(n_266),
.B1(n_235),
.B2(n_251),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_278),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_320),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_296),
.A2(n_302),
.B1(n_310),
.B2(n_309),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_317),
.A2(n_315),
.B1(n_268),
.B2(n_271),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_SL g319 ( 
.A1(n_295),
.A2(n_280),
.B(n_293),
.C(n_290),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_319),
.A2(n_315),
.B(n_297),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_294),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_300),
.A2(n_275),
.B(n_276),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_327),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_313),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_308),
.Y(n_328)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_328),
.Y(n_335)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_329),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_311),
.B(n_275),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_332),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_333),
.A2(n_326),
.B(n_319),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_314),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_339),
.Y(n_349)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_337),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_303),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_338),
.B(n_341),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_324),
.A2(n_263),
.B1(n_261),
.B2(n_267),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_299),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_328),
.A2(n_325),
.B1(n_306),
.B2(n_318),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_343),
.B(n_344),
.Y(n_355)
);

INVx6_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_344),
.B(n_345),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_330),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_341),
.B(n_322),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_352),
.Y(n_359)
);

AO21x1_ASAP7_75t_L g363 ( 
.A1(n_351),
.A2(n_354),
.B(n_355),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_346),
.B(n_322),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_333),
.A2(n_319),
.B(n_326),
.Y(n_353)
);

OAI21x1_ASAP7_75t_L g358 ( 
.A1(n_353),
.A2(n_340),
.B(n_338),
.Y(n_358)
);

OA21x2_ASAP7_75t_SL g354 ( 
.A1(n_342),
.A2(n_306),
.B(n_316),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_332),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_357),
.B(n_334),
.Y(n_360)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_358),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_360),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_356),
.B(n_244),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_361),
.B(n_365),
.Y(n_370)
);

OAI321xp33_ASAP7_75t_L g362 ( 
.A1(n_349),
.A2(n_271),
.A3(n_346),
.B1(n_334),
.B2(n_190),
.C(n_212),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_362),
.A2(n_209),
.B1(n_213),
.B2(n_353),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_179),
.C(n_198),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_364),
.B(n_367),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_348),
.A2(n_212),
.B1(n_222),
.B2(n_198),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_351),
.A2(n_212),
.B1(n_222),
.B2(n_160),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_366),
.B(n_222),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_357),
.A2(n_192),
.B(n_193),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_360),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_369),
.B(n_375),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_371),
.Y(n_379)
);

AOI322xp5_ASAP7_75t_L g376 ( 
.A1(n_373),
.A2(n_363),
.A3(n_146),
.B1(n_193),
.B2(n_186),
.C1(n_201),
.C2(n_209),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_350),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_376),
.B(n_378),
.Y(n_381)
);

AOI322xp5_ASAP7_75t_L g378 ( 
.A1(n_374),
.A2(n_359),
.A3(n_352),
.B1(n_146),
.B2(n_186),
.C1(n_201),
.C2(n_210),
.Y(n_378)
);

AOI21x1_ASAP7_75t_L g380 ( 
.A1(n_372),
.A2(n_210),
.B(n_147),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_380),
.A2(n_370),
.B(n_368),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_382),
.B(n_379),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_377),
.A2(n_369),
.B(n_5),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_383),
.A2(n_5),
.B(n_96),
.Y(n_385)
);

NOR3xp33_ASAP7_75t_L g386 ( 
.A(n_384),
.B(n_385),
.C(n_381),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_5),
.Y(n_387)
);


endmodule