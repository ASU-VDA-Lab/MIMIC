module fake_jpeg_29422_n_347 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_21),
.B(n_9),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_49),
.B(n_56),
.Y(n_109)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_21),
.B(n_9),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_58),
.B(n_59),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_17),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_19),
.B(n_8),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_71),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_31),
.B(n_1),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_70),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_76),
.B(n_5),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_31),
.B1(n_41),
.B2(n_38),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_77),
.A2(n_83),
.B1(n_92),
.B2(n_95),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_24),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_80),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_79),
.B(n_28),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_24),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_30),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_91),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_41),
.B1(n_43),
.B2(n_42),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_19),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_88),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_25),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_36),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_35),
.B1(n_26),
.B2(n_41),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_43),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_106),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_23),
.B1(n_40),
.B2(n_39),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_57),
.A2(n_26),
.B1(n_53),
.B2(n_55),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_98),
.A2(n_107),
.B1(n_110),
.B2(n_111),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_46),
.B(n_28),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_28),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_48),
.B(n_36),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_45),
.A2(n_52),
.B1(n_65),
.B2(n_63),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_42),
.B1(n_26),
.B2(n_40),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_60),
.A2(n_44),
.B1(n_39),
.B2(n_34),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_51),
.A2(n_44),
.B1(n_34),
.B2(n_33),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_117),
.A2(n_47),
.B1(n_8),
.B2(n_12),
.Y(n_142)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_60),
.B1(n_33),
.B2(n_27),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_125),
.A2(n_96),
.B1(n_118),
.B2(n_112),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_149),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_27),
.C(n_60),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_127),
.B(n_137),
.C(n_115),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_79),
.A2(n_10),
.B(n_12),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_128),
.B(n_159),
.Y(n_173)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_76),
.A2(n_28),
.B1(n_12),
.B2(n_16),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_86),
.B(n_28),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_139),
.B(n_115),
.Y(n_186)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_114),
.B1(n_101),
.B2(n_109),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_88),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_147),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_81),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_90),
.A2(n_5),
.B(n_14),
.C(n_13),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_148),
.A2(n_109),
.B(n_13),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_86),
.B(n_1),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_75),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_152),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_102),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_153),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_95),
.B(n_2),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_157),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_100),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_132),
.Y(n_185)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_3),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_85),
.B1(n_74),
.B2(n_112),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_160),
.A2(n_164),
.B1(n_142),
.B2(n_127),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_171),
.A2(n_187),
.B1(n_189),
.B2(n_150),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_147),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_183),
.Y(n_196)
);

BUFx8_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_179),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_157),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_74),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_124),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_188),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_85),
.B1(n_74),
.B2(n_96),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_143),
.A2(n_84),
.B1(n_116),
.B2(n_108),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_101),
.B1(n_152),
.B2(n_146),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_116),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_153),
.Y(n_197)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_192),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_137),
.B(n_84),
.C(n_100),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_155),
.C(n_144),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_198),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_183),
.Y(n_198)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_126),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_202),
.B(n_208),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_203),
.A2(n_225),
.B1(n_217),
.B2(n_226),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_204),
.B(n_211),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_16),
.C(n_3),
.Y(n_245)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_139),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_210),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_139),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_213),
.B(n_214),
.Y(n_243)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_179),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_215),
.B(n_219),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_216),
.A2(n_193),
.B1(n_167),
.B2(n_184),
.Y(n_254)
);

NAND2x1p5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_134),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_218),
.A2(n_221),
.B(n_181),
.Y(n_239)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_151),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_223),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_169),
.A2(n_145),
.B(n_148),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_222),
.A2(n_177),
.B1(n_99),
.B2(n_118),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_172),
.B(n_136),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_226),
.C(n_140),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_160),
.A2(n_170),
.B1(n_176),
.B2(n_164),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_129),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_173),
.B(n_138),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_179),
.Y(n_244)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_230),
.A2(n_254),
.B1(n_202),
.B2(n_218),
.Y(n_273)
);

AOI322xp5_ASAP7_75t_L g231 ( 
.A1(n_221),
.A2(n_182),
.A3(n_194),
.B1(n_191),
.B2(n_189),
.C1(n_89),
.C2(n_177),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_244),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_252),
.C(n_211),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_238),
.A2(n_249),
.B1(n_199),
.B2(n_214),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_228),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_197),
.A2(n_181),
.B(n_166),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_240),
.A2(n_208),
.B(n_196),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_245),
.B(n_205),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_224),
.A2(n_193),
.B(n_184),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_248),
.A2(n_255),
.B(n_256),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_222),
.A2(n_167),
.B1(n_99),
.B2(n_119),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_200),
.Y(n_251)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_251),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_195),
.C(n_156),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_204),
.A2(n_195),
.B(n_122),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_218),
.A2(n_162),
.B(n_158),
.Y(n_256)
);

NAND3xp33_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_242),
.C(n_250),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_236),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_259),
.B(n_239),
.Y(n_284)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_261),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_266),
.C(n_274),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_264),
.A2(n_271),
.B1(n_277),
.B2(n_254),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_196),
.C(n_198),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_268),
.Y(n_282)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_232),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_237),
.B(n_253),
.Y(n_289)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_233),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_272),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_203),
.B1(n_199),
.B2(n_213),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_209),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_229),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_207),
.C(n_210),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_131),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_241),
.A2(n_219),
.B(n_201),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_276),
.A2(n_278),
.B(n_235),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_133),
.B1(n_212),
.B2(n_130),
.Y(n_277)
);

NAND2xp33_ASAP7_75t_SL g278 ( 
.A(n_255),
.B(n_175),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_294),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_280),
.A2(n_283),
.B1(n_288),
.B2(n_273),
.Y(n_301)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_271),
.A2(n_242),
.B1(n_250),
.B2(n_252),
.Y(n_283)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_284),
.Y(n_302)
);

NOR3xp33_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_246),
.C(n_233),
.Y(n_287)
);

NOR3xp33_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_291),
.C(n_295),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_264),
.A2(n_237),
.B1(n_248),
.B2(n_246),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_293),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_253),
.C(n_235),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_260),
.C(n_275),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_229),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_294),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_274),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_305),
.C(n_309),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_285),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_260),
.B(n_269),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_299),
.A2(n_272),
.B(n_290),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_289),
.B1(n_272),
.B2(n_281),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_308),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_266),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_262),
.C(n_276),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_277),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_280),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_296),
.B(n_270),
.Y(n_311)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_311),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_318),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_313),
.A2(n_298),
.B(n_304),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_322),
.Y(n_329)
);

OAI21xp33_ASAP7_75t_L g316 ( 
.A1(n_306),
.A2(n_282),
.B(n_285),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_258),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_317),
.A2(n_315),
.B1(n_321),
.B2(n_316),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_302),
.A2(n_282),
.B1(n_268),
.B2(n_267),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_300),
.A2(n_288),
.B1(n_283),
.B2(n_278),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_321),
.A2(n_305),
.B1(n_299),
.B2(n_309),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_303),
.B(n_258),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_324),
.A2(n_322),
.B1(n_175),
.B2(n_89),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_297),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_326),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_303),
.C(n_304),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_327),
.A2(n_330),
.B(n_97),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_328),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_320),
.B(n_179),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_4),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_323),
.A2(n_313),
.B1(n_319),
.B2(n_314),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_333),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_229),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_334),
.B(n_336),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_337),
.B(n_4),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_335),
.A2(n_330),
.B(n_332),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_340),
.B(n_342),
.Y(n_343)
);

AOI321xp33_ASAP7_75t_L g344 ( 
.A1(n_339),
.A2(n_338),
.A3(n_324),
.B1(n_334),
.B2(n_336),
.C(n_329),
.Y(n_344)
);

AOI31xp67_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_341),
.A3(n_329),
.B(n_97),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_343),
.C(n_4),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_4),
.Y(n_347)
);


endmodule