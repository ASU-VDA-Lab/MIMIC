module real_aes_5034_n_14 (n_13, n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_10, n_11, n_14);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_10;
input n_11;
output n_14;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_34;
wire n_19;
wire n_25;
wire n_32;
wire n_30;
wire n_16;
wire n_37;
wire n_35;
wire n_15;
wire n_27;
wire n_23;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g25 ( .A(n_1), .Y(n_25) );
AOI22xp33_ASAP7_75t_R g29 ( .A1(n_2), .A2(n_8), .B1(n_30), .B2(n_35), .Y(n_29) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_3), .Y(n_24) );
NOR2xp33_ASAP7_75t_R g19 ( .A(n_4), .B(n_20), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_5), .Y(n_27) );
NOR4xp25_ASAP7_75t_SL g17 ( .A(n_6), .B(n_18), .C(n_24), .D(n_25), .Y(n_17) );
NAND2xp33_ASAP7_75t_R g33 ( .A(n_6), .B(n_19), .Y(n_33) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_7), .Y(n_26) );
NAND2xp33_ASAP7_75t_R g28 ( .A(n_7), .B(n_17), .Y(n_28) );
NOR2xp33_ASAP7_75t_R g30 ( .A(n_7), .B(n_31), .Y(n_30) );
NAND2xp33_ASAP7_75t_R g37 ( .A(n_7), .B(n_32), .Y(n_37) );
NAND3xp33_ASAP7_75t_SL g20 ( .A(n_9), .B(n_21), .C(n_22), .Y(n_20) );
NOR2xp33_ASAP7_75t_R g23 ( .A(n_10), .B(n_11), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_12), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_13), .Y(n_22) );
OAI221xp5_ASAP7_75t_R g14 ( .A1(n_15), .A2(n_16), .B1(n_27), .B2(n_28), .C(n_29), .Y(n_14) );
NAND2xp33_ASAP7_75t_R g16 ( .A(n_17), .B(n_26), .Y(n_16) );
NAND2xp33_ASAP7_75t_R g18 ( .A(n_19), .B(n_23), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g34 ( .A(n_23), .Y(n_34) );
NOR4xp25_ASAP7_75t_SL g32 ( .A(n_24), .B(n_25), .C(n_33), .D(n_34), .Y(n_32) );
CKINVDCx5p33_ASAP7_75t_R g31 ( .A(n_32), .Y(n_31) );
HB1xp67_ASAP7_75t_L g35 ( .A(n_36), .Y(n_35) );
CKINVDCx5p33_ASAP7_75t_R g36 ( .A(n_37), .Y(n_36) );
endmodule