module fake_jpeg_26241_n_221 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_221);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_221;

wire n_159;
wire n_117;
wire n_144;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_12),
.B(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_31),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_0),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_30),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_20),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_23),
.A2(n_22),
.B1(n_11),
.B2(n_14),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_24),
.B1(n_28),
.B2(n_25),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_31),
.B(n_29),
.C(n_26),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_53),
.B(n_33),
.C(n_31),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_11),
.B1(n_22),
.B2(n_28),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_55),
.B1(n_25),
.B2(n_31),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_23),
.B1(n_24),
.B2(n_31),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_47),
.Y(n_73)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_33),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_11),
.B1(n_22),
.B2(n_12),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_58),
.B1(n_25),
.B2(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_54),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_31),
.B(n_15),
.C(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_23),
.B1(n_24),
.B2(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_64),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_62),
.A2(n_70),
.B1(n_77),
.B2(n_27),
.Y(n_98)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_55),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_47),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_20),
.C(n_10),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_33),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_33),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_53),
.B(n_52),
.C(n_44),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_38),
.B1(n_34),
.B2(n_30),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_80),
.B(n_98),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_72),
.B1(n_74),
.B2(n_70),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_68),
.B1(n_61),
.B2(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_46),
.B1(n_30),
.B2(n_38),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_88),
.B(n_92),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_38),
.Y(n_89)
);

OAI31xp33_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_30),
.A3(n_27),
.B(n_36),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_65),
.Y(n_101)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_71),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_95),
.Y(n_118)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_76),
.B1(n_51),
.B2(n_27),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_106),
.B(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_67),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_110),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_104),
.B(n_114),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_86),
.B(n_91),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_115),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_68),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_81),
.Y(n_132)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_119),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_87),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_36),
.B1(n_27),
.B2(n_35),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_36),
.Y(n_123)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_133),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_86),
.B1(n_85),
.B2(n_92),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_138),
.B1(n_139),
.B2(n_142),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_78),
.B(n_80),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_111),
.B(n_109),
.Y(n_148)
);

FAx1_ASAP7_75t_SL g164 ( 
.A(n_132),
.B(n_16),
.CI(n_13),
.CON(n_164),
.SN(n_164)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_90),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_104),
.B(n_30),
.CI(n_27),
.CON(n_134),
.SN(n_134)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_113),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_36),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_140),
.C(n_133),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_15),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_137),
.B(n_105),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_17),
.B1(n_19),
.B2(n_21),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_6),
.B(n_9),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_56),
.C(n_36),
.Y(n_140)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_99),
.A2(n_19),
.A3(n_17),
.B1(n_10),
.B2(n_21),
.Y(n_143)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_13),
.B1(n_16),
.B2(n_8),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_21),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_147),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_148),
.A2(n_154),
.B(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_151),
.B(n_153),
.Y(n_167)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_129),
.B(n_107),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_108),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_164),
.C(n_165),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_159),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_109),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_136),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_SL g177 ( 
.A1(n_161),
.A2(n_134),
.B(n_144),
.C(n_127),
.Y(n_177)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_130),
.B1(n_134),
.B2(n_128),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_116),
.C(n_36),
.Y(n_165)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

NOR2x1_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_143),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_172),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_157),
.B1(n_160),
.B2(n_150),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_178),
.B1(n_164),
.B2(n_36),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_132),
.C(n_140),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_128),
.C(n_135),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_179),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_16),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_160),
.B1(n_148),
.B2(n_152),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_142),
.C(n_10),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_169),
.A2(n_159),
.B1(n_164),
.B2(n_155),
.Y(n_180)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_183),
.B(n_188),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_186),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_35),
.C(n_27),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_167),
.C(n_174),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_177),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_188)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_189),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_177),
.A2(n_6),
.B(n_8),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_190),
.A2(n_7),
.B(n_8),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_195),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_196),
.A2(n_190),
.B(n_184),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_181),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_193),
.B(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_191),
.B(n_176),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_202),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_193),
.B(n_187),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_188),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_204),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_194),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_206),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_208),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_180),
.C(n_186),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_7),
.B(n_3),
.Y(n_214)
);

OA21x2_ASAP7_75t_SL g213 ( 
.A1(n_210),
.A2(n_189),
.B(n_7),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_214),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_207),
.B1(n_211),
.B2(n_208),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_216),
.A2(n_212),
.B(n_3),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_218),
.A2(n_217),
.B(n_4),
.Y(n_219)
);

OAI321xp33_ASAP7_75t_L g220 ( 
.A1(n_219),
.A2(n_1),
.A3(n_4),
.B1(n_5),
.B2(n_35),
.C(n_203),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_SL g221 ( 
.A(n_220),
.B(n_4),
.C(n_5),
.Y(n_221)
);


endmodule