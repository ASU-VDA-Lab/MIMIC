module real_aes_1872_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_755;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_0), .B(n_138), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_1), .A2(n_31), .B1(n_463), .B2(n_464), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_1), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_2), .A2(n_147), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_3), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_4), .B(n_138), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_5), .B(n_154), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_6), .B(n_154), .Y(n_546) );
INVx1_ASAP7_75t_L g145 ( .A(n_7), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_8), .B(n_154), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_9), .Y(n_109) );
NAND2xp33_ASAP7_75t_L g523 ( .A(n_10), .B(n_156), .Y(n_523) );
AND2x2_ASAP7_75t_L g175 ( .A(n_11), .B(n_163), .Y(n_175) );
AND2x2_ASAP7_75t_L g184 ( .A(n_12), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g160 ( .A(n_13), .Y(n_160) );
AOI221x1_ASAP7_75t_L g476 ( .A1(n_14), .A2(n_25), .B1(n_138), .B2(n_147), .C(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_15), .B(n_154), .Y(n_193) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_16), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_17), .B(n_138), .Y(n_519) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_18), .A2(n_163), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_19), .B(n_158), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_20), .B(n_154), .Y(n_530) );
AO21x1_ASAP7_75t_L g541 ( .A1(n_21), .A2(n_138), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_22), .B(n_138), .Y(n_218) );
INVx1_ASAP7_75t_L g106 ( .A(n_23), .Y(n_106) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_24), .A2(n_90), .B1(n_138), .B2(n_248), .Y(n_247) );
NAND2x1_ASAP7_75t_L g486 ( .A(n_26), .B(n_154), .Y(n_486) );
NAND2x1_ASAP7_75t_L g512 ( .A(n_27), .B(n_156), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_28), .Y(n_459) );
OR2x2_ASAP7_75t_L g161 ( .A(n_29), .B(n_87), .Y(n_161) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_29), .A2(n_87), .B(n_160), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_30), .B(n_156), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_31), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_32), .B(n_154), .Y(n_522) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_33), .A2(n_185), .B(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_34), .B(n_156), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_35), .A2(n_147), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_36), .B(n_154), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_37), .A2(n_147), .B(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g144 ( .A(n_38), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g148 ( .A(n_38), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g256 ( .A(n_38), .Y(n_256) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_39), .B(n_108), .C(n_110), .Y(n_107) );
OR2x6_ASAP7_75t_L g121 ( .A(n_39), .B(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_40), .B(n_138), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_41), .B(n_138), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_42), .B(n_154), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_43), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_44), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_45), .B(n_156), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_46), .B(n_138), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_47), .A2(n_147), .B(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_48), .A2(n_147), .B(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_49), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_50), .B(n_156), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_51), .B(n_138), .Y(n_190) );
INVx1_ASAP7_75t_L g141 ( .A(n_52), .Y(n_141) );
INVx1_ASAP7_75t_L g151 ( .A(n_52), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_53), .B(n_154), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_54), .A2(n_61), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_54), .Y(n_127) );
AND2x2_ASAP7_75t_L g209 ( .A(n_55), .B(n_158), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_56), .B(n_156), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_57), .B(n_154), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_58), .B(n_156), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_59), .A2(n_147), .B(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_60), .B(n_138), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_61), .Y(n_128) );
INVxp33_ASAP7_75t_L g763 ( .A(n_62), .Y(n_763) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_63), .B(n_138), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_64), .A2(n_147), .B(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g224 ( .A(n_65), .B(n_159), .Y(n_224) );
AO21x1_ASAP7_75t_L g543 ( .A1(n_66), .A2(n_147), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_67), .B(n_138), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_68), .B(n_156), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_69), .B(n_138), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_70), .B(n_156), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_71), .A2(n_95), .B1(n_147), .B2(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_72), .B(n_154), .Y(n_221) );
AND2x2_ASAP7_75t_L g497 ( .A(n_73), .B(n_159), .Y(n_497) );
INVx1_ASAP7_75t_L g143 ( .A(n_74), .Y(n_143) );
INVx1_ASAP7_75t_L g149 ( .A(n_74), .Y(n_149) );
AND2x2_ASAP7_75t_L g515 ( .A(n_75), .B(n_185), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_76), .B(n_156), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_77), .A2(n_147), .B(n_213), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_78), .A2(n_147), .B(n_152), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_79), .A2(n_147), .B(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g204 ( .A(n_80), .B(n_159), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_81), .B(n_158), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_82), .B(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g123 ( .A(n_82), .Y(n_123) );
AND2x2_ASAP7_75t_L g501 ( .A(n_83), .B(n_185), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_84), .B(n_138), .Y(n_532) );
AND2x2_ASAP7_75t_L g162 ( .A(n_85), .B(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g542 ( .A(n_86), .B(n_195), .Y(n_542) );
AND2x2_ASAP7_75t_L g489 ( .A(n_88), .B(n_185), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_89), .B(n_156), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_91), .B(n_154), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_92), .B(n_156), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_93), .A2(n_147), .B(n_529), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_94), .A2(n_147), .B(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_96), .B(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_97), .B(n_154), .Y(n_506) );
BUFx2_ASAP7_75t_L g223 ( .A(n_98), .Y(n_223) );
BUFx2_ASAP7_75t_L g116 ( .A(n_99), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_100), .A2(n_147), .B(n_521), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_111), .B(n_762), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g765 ( .A(n_103), .Y(n_765) );
INVx3_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_SL g104 ( .A(n_105), .B(n_107), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_106), .B(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_110), .B(n_120), .Y(n_119) );
OR2x6_ASAP7_75t_SL g748 ( .A(n_110), .B(n_120), .Y(n_748) );
AND2x6_ASAP7_75t_SL g750 ( .A(n_110), .B(n_121), .Y(n_750) );
OR2x2_ASAP7_75t_L g759 ( .A(n_110), .B(n_121), .Y(n_759) );
OR2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_460), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_117), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx3_ASAP7_75t_L g761 ( .A(n_114), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_124), .B(n_458), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_118), .B(n_459), .Y(n_458) );
BUFx2_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
NAND2x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_455), .Y(n_124) );
NAND2x1p5_ASAP7_75t_L g125 ( .A(n_126), .B(n_129), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_126), .Y(n_457) );
INVx4_ASAP7_75t_L g456 ( .A(n_129), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_129), .A2(n_467), .B1(n_748), .B2(n_752), .Y(n_751) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_363), .Y(n_129) );
NOR3xp33_ASAP7_75t_SL g130 ( .A(n_131), .B(n_286), .C(n_321), .Y(n_130) );
OAI211xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_186), .B(n_238), .C(n_276), .Y(n_131) );
INVx1_ASAP7_75t_SL g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_165), .Y(n_133) );
AND2x2_ASAP7_75t_L g269 ( .A(n_134), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_134), .B(n_275), .Y(n_309) );
AND2x2_ASAP7_75t_L g334 ( .A(n_134), .B(n_289), .Y(n_334) );
INVx4_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx2_ASAP7_75t_L g241 ( .A(n_135), .Y(n_241) );
OR2x2_ASAP7_75t_L g272 ( .A(n_135), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g280 ( .A(n_135), .B(n_176), .Y(n_280) );
AND2x2_ASAP7_75t_L g288 ( .A(n_135), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g315 ( .A(n_135), .B(n_316), .Y(n_315) );
NOR2x1_ASAP7_75t_L g326 ( .A(n_135), .B(n_318), .Y(n_326) );
AND2x4_ASAP7_75t_L g343 ( .A(n_135), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g381 ( .A(n_135), .Y(n_381) );
AND2x4_ASAP7_75t_SL g386 ( .A(n_135), .B(n_166), .Y(n_386) );
OR2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_162), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_146), .B(n_158), .Y(n_136) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_144), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
AND2x6_ASAP7_75t_L g156 ( .A(n_140), .B(n_149), .Y(n_156) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g154 ( .A(n_142), .B(n_151), .Y(n_154) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx5_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
AND2x2_ASAP7_75t_L g150 ( .A(n_145), .B(n_151), .Y(n_150) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_145), .Y(n_251) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
BUFx3_ASAP7_75t_L g252 ( .A(n_148), .Y(n_252) );
INVx2_ASAP7_75t_L g258 ( .A(n_149), .Y(n_258) );
AND2x4_ASAP7_75t_L g254 ( .A(n_150), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g250 ( .A(n_151), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_155), .B(n_157), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_156), .B(n_223), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_157), .A2(n_172), .B(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_157), .A2(n_181), .B(n_182), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_157), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_157), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_157), .A2(n_214), .B(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_157), .A2(n_221), .B(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_157), .A2(n_478), .B(n_479), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_157), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_157), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_157), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_157), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_157), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_157), .A2(n_530), .B(n_531), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_157), .A2(n_545), .B(n_546), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_158), .Y(n_168) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_158), .A2(n_247), .B(n_253), .Y(n_246) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_158), .A2(n_476), .B(n_480), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_158), .A2(n_503), .B(n_504), .Y(n_502) );
OA21x2_ASAP7_75t_L g582 ( .A1(n_158), .A2(n_476), .B(n_480), .Y(n_582) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_160), .B(n_161), .Y(n_159) );
AND2x4_ASAP7_75t_L g195 ( .A(n_160), .B(n_161), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_163), .A2(n_218), .B(n_219), .Y(n_217) );
BUFx4f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx3_ASAP7_75t_L g177 ( .A(n_164), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_165), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_165), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_176), .Y(n_165) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_166), .Y(n_281) );
INVx2_ASAP7_75t_L g317 ( .A(n_166), .Y(n_317) );
INVx1_ASAP7_75t_L g344 ( .A(n_166), .Y(n_344) );
AND2x2_ASAP7_75t_L g443 ( .A(n_166), .B(n_353), .Y(n_443) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_167), .Y(n_275) );
AND2x2_ASAP7_75t_L g289 ( .A(n_167), .B(n_176), .Y(n_289) );
AOI21x1_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_175), .Y(n_167) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_168), .A2(n_509), .B(n_515), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_174), .Y(n_169) );
INVx2_ASAP7_75t_L g318 ( .A(n_176), .Y(n_318) );
INVx2_ASAP7_75t_L g353 ( .A(n_176), .Y(n_353) );
OR2x2_ASAP7_75t_L g438 ( .A(n_176), .B(n_270), .Y(n_438) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_184), .Y(n_176) );
INVx4_ASAP7_75t_L g185 ( .A(n_177), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_183), .Y(n_178) );
INVx3_ASAP7_75t_L g197 ( .A(n_185), .Y(n_197) );
AOI211xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_205), .B(n_225), .C(n_232), .Y(n_186) );
INVx2_ASAP7_75t_SL g327 ( .A(n_187), .Y(n_327) );
AND2x2_ASAP7_75t_L g333 ( .A(n_187), .B(n_206), .Y(n_333) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_196), .Y(n_187) );
INVx1_ASAP7_75t_L g229 ( .A(n_188), .Y(n_229) );
INVx1_ASAP7_75t_L g235 ( .A(n_188), .Y(n_235) );
INVx2_ASAP7_75t_L g260 ( .A(n_188), .Y(n_260) );
AND2x2_ASAP7_75t_L g284 ( .A(n_188), .B(n_208), .Y(n_284) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_188), .Y(n_313) );
OR2x2_ASAP7_75t_L g393 ( .A(n_188), .B(n_216), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_195), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_195), .A2(n_211), .B(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_195), .A2(n_519), .B(n_520), .Y(n_518) );
INVx1_ASAP7_75t_SL g526 ( .A(n_195), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_195), .B(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g259 ( .A(n_196), .B(n_260), .Y(n_259) );
NOR2x1_ASAP7_75t_SL g291 ( .A(n_196), .B(n_216), .Y(n_291) );
AO21x1_ASAP7_75t_SL g196 ( .A1(n_197), .A2(n_198), .B(n_204), .Y(n_196) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_197), .A2(n_198), .B(n_204), .Y(n_231) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_197), .A2(n_483), .B(n_489), .Y(n_482) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_197), .A2(n_491), .B(n_497), .Y(n_490) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_197), .A2(n_491), .B(n_497), .Y(n_549) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_197), .A2(n_483), .B(n_489), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_203), .Y(n_198) );
INVxp67_ASAP7_75t_SL g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g305 ( .A(n_206), .B(n_228), .Y(n_305) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_216), .Y(n_206) );
OR2x2_ASAP7_75t_L g237 ( .A(n_207), .B(n_216), .Y(n_237) );
BUFx2_ASAP7_75t_L g261 ( .A(n_207), .Y(n_261) );
NOR2xp67_ASAP7_75t_L g312 ( .A(n_207), .B(n_313), .Y(n_312) );
INVx4_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_208), .Y(n_264) );
AND2x2_ASAP7_75t_L g290 ( .A(n_208), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g300 ( .A(n_208), .Y(n_300) );
NAND2x1_ASAP7_75t_L g338 ( .A(n_208), .B(n_216), .Y(n_338) );
OR2x2_ASAP7_75t_L g413 ( .A(n_208), .B(n_230), .Y(n_413) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
INVx2_ASAP7_75t_SL g226 ( .A(n_216), .Y(n_226) );
AND2x2_ASAP7_75t_L g285 ( .A(n_216), .B(n_230), .Y(n_285) );
AND2x2_ASAP7_75t_L g356 ( .A(n_216), .B(n_357), .Y(n_356) );
BUFx2_ASAP7_75t_L g377 ( .A(n_216), .Y(n_377) );
OR2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_224), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
INVx1_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g299 ( .A(n_228), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
BUFx2_ASAP7_75t_L g294 ( .A(n_229), .Y(n_294) );
AND2x2_ASAP7_75t_L g266 ( .A(n_230), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g357 ( .A(n_230), .Y(n_357) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_236), .Y(n_233) );
OR2x2_ASAP7_75t_L g303 ( .A(n_234), .B(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_SL g345 ( .A(n_234), .B(n_346), .Y(n_345) );
AOI322xp5_ASAP7_75t_L g382 ( .A1(n_234), .A2(n_261), .A3(n_383), .B1(n_385), .B2(n_388), .C1(n_390), .C2(n_392), .Y(n_382) );
AND2x2_ASAP7_75t_L g447 ( .A(n_234), .B(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_235), .B(n_261), .Y(n_271) );
AOI322xp5_ASAP7_75t_L g322 ( .A1(n_236), .A2(n_323), .A3(n_327), .B1(n_328), .B2(n_331), .C1(n_333), .C2(n_334), .Y(n_322) );
INVx2_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g374 ( .A(n_237), .B(n_327), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_237), .A2(n_434), .B1(n_436), .B2(n_439), .Y(n_433) );
OR2x2_ASAP7_75t_L g451 ( .A(n_237), .B(n_400), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_261), .B(n_262), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
AOI221xp5_ASAP7_75t_SL g301 ( .A1(n_240), .A2(n_277), .B1(n_302), .B2(n_305), .C(n_306), .Y(n_301) );
AND2x2_ASAP7_75t_L g328 ( .A(n_240), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_241), .B(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g370 ( .A(n_241), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g399 ( .A(n_242), .Y(n_399) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_259), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_243), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g341 ( .A(n_243), .Y(n_341) );
OR2x2_ASAP7_75t_L g348 ( .A(n_243), .B(n_349), .Y(n_348) );
INVx3_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g391 ( .A(n_244), .B(n_353), .Y(n_391) );
AND2x4_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
AND2x4_ASAP7_75t_L g270 ( .A(n_245), .B(n_246), .Y(n_270) );
AND2x4_ASAP7_75t_L g248 ( .A(n_249), .B(n_252), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NOR2x1p5_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_259), .B(n_320), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_259), .B(n_300), .Y(n_396) );
INVx1_ASAP7_75t_L g400 ( .A(n_259), .Y(n_400) );
INVx1_ASAP7_75t_L g267 ( .A(n_260), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_268), .B1(n_271), .B2(n_272), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
BUFx2_ASAP7_75t_SL g378 ( .A(n_266), .Y(n_378) );
AND2x2_ASAP7_75t_L g435 ( .A(n_267), .B(n_291), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_269), .B(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_SL g307 ( .A(n_269), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_269), .B(n_428), .Y(n_427) );
BUFx3_ASAP7_75t_L g295 ( .A(n_270), .Y(n_295) );
INVx2_ASAP7_75t_L g325 ( .A(n_270), .Y(n_325) );
AND2x2_ASAP7_75t_L g368 ( .A(n_270), .B(n_352), .Y(n_368) );
INVx1_ASAP7_75t_L g282 ( .A(n_272), .Y(n_282) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OAI21xp5_ASAP7_75t_SL g276 ( .A1(n_277), .A2(n_282), .B(n_283), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g361 ( .A(n_280), .Y(n_361) );
INVx2_ASAP7_75t_L g349 ( .A(n_281), .Y(n_349) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x2_ASAP7_75t_L g346 ( .A(n_285), .B(n_300), .Y(n_346) );
OAI21xp5_ASAP7_75t_L g406 ( .A1(n_285), .A2(n_383), .B(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_287), .B(n_301), .Y(n_286) );
AOI32xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_290), .A3(n_292), .B1(n_296), .B2(n_299), .Y(n_287) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_288), .Y(n_362) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_288), .A2(n_377), .B1(n_395), .B2(n_397), .C(n_403), .Y(n_394) );
AND2x2_ASAP7_75t_L g414 ( .A(n_288), .B(n_295), .Y(n_414) );
BUFx2_ASAP7_75t_L g298 ( .A(n_289), .Y(n_298) );
INVx1_ASAP7_75t_L g423 ( .A(n_289), .Y(n_423) );
INVx1_ASAP7_75t_L g428 ( .A(n_289), .Y(n_428) );
INVx1_ASAP7_75t_SL g421 ( .A(n_290), .Y(n_421) );
INVx2_ASAP7_75t_L g304 ( .A(n_291), .Y(n_304) );
AND2x2_ASAP7_75t_L g416 ( .A(n_292), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x2_ASAP7_75t_L g388 ( .A(n_294), .B(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g360 ( .A(n_295), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_295), .B(n_386), .Y(n_408) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g320 ( .A(n_300), .Y(n_320) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g310 ( .A(n_304), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g319 ( .A(n_304), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g424 ( .A(n_305), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_310), .B1(n_314), .B2(n_319), .Y(n_306) );
INVx2_ASAP7_75t_SL g398 ( .A(n_308), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_308), .B(n_437), .Y(n_439) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_310), .A2(n_404), .B(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g355 ( .A(n_312), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g383 ( .A(n_315), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g330 ( .A(n_316), .Y(n_330) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g372 ( .A(n_318), .Y(n_372) );
INVx1_ASAP7_75t_L g417 ( .A(n_319), .Y(n_417) );
NAND3xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_335), .C(n_358), .Y(n_321) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
INVx2_ASAP7_75t_L g384 ( .A(n_324), .Y(n_384) );
AND2x2_ASAP7_75t_L g402 ( .A(n_324), .B(n_343), .Y(n_402) );
OR2x2_ASAP7_75t_L g441 ( .A(n_324), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_325), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g337 ( .A(n_327), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g404 ( .A(n_330), .B(n_341), .Y(n_404) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_333), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g445 ( .A(n_333), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_339), .B1(n_343), .B2(n_345), .C(n_347), .Y(n_335) );
OAI21xp5_ASAP7_75t_L g358 ( .A1(n_336), .A2(n_359), .B(n_362), .Y(n_358) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx3_ASAP7_75t_L g389 ( .A(n_338), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_338), .B(n_432), .Y(n_431) );
INVxp33_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g350 ( .A(n_346), .Y(n_350) );
OAI22xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_350), .B1(n_351), .B2(n_354), .Y(n_347) );
INVx2_ASAP7_75t_L g453 ( .A(n_349), .Y(n_453) );
BUFx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVxp67_ASAP7_75t_L g432 ( .A(n_357), .Y(n_432) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
NOR2x1_ASAP7_75t_L g363 ( .A(n_364), .B(n_409), .Y(n_363) );
NAND4xp25_ASAP7_75t_L g364 ( .A(n_365), .B(n_382), .C(n_394), .D(n_406), .Y(n_364) );
O2A1O1Ixp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_369), .B(n_373), .C(n_375), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g405 ( .A(n_368), .Y(n_405) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI21xp5_ASAP7_75t_L g375 ( .A1(n_370), .A2(n_376), .B(n_379), .Y(n_375) );
INVx2_ASAP7_75t_L g454 ( .A(n_371), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_372), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g387 ( .A(n_372), .Y(n_387) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
OR2x2_ASAP7_75t_L g449 ( .A(n_377), .B(n_413), .Y(n_449) );
INVxp67_ASAP7_75t_SL g420 ( .A(n_384), .Y(n_420) );
AND2x2_ASAP7_75t_SL g385 ( .A(n_386), .B(n_387), .Y(n_385) );
AND2x2_ASAP7_75t_L g390 ( .A(n_386), .B(n_391), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_386), .A2(n_416), .B(n_418), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_386), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_SL g444 ( .A(n_386), .Y(n_444) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI22xp33_ASAP7_75t_SL g397 ( .A1(n_398), .A2(n_399), .B1(n_400), .B2(n_401), .Y(n_397) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND4xp25_ASAP7_75t_L g409 ( .A(n_410), .B(n_415), .C(n_425), .D(n_446), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .B1(n_422), .B2(n_424), .Y(n_418) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI211xp5_ASAP7_75t_SL g425 ( .A1(n_426), .A2(n_429), .B(n_433), .C(n_440), .Y(n_425) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
AOI21xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_444), .B(n_445), .Y(n_440) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
OAI21xp5_ASAP7_75t_SL g446 ( .A1(n_447), .A2(n_450), .B(n_452), .Y(n_446) );
INVx1_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
OAI22x1_ASAP7_75t_L g465 ( .A1(n_456), .A2(n_466), .B1(n_746), .B2(n_749), .Y(n_465) );
INVxp33_ASAP7_75t_L g760 ( .A(n_458), .Y(n_760) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_760), .B(n_761), .Y(n_460) );
AOI221xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_465), .B1(n_751), .B2(n_754), .C(n_755), .Y(n_461) );
INVx1_ASAP7_75t_L g754 ( .A(n_462), .Y(n_754) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_658), .Y(n_467) );
AND4x1_ASAP7_75t_L g468 ( .A(n_469), .B(n_570), .C(n_597), .D(n_632), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_498), .B1(n_535), .B2(n_550), .C(n_554), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_481), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_472), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g611 ( .A(n_473), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g666 ( .A(n_473), .B(n_621), .Y(n_666) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g569 ( .A(n_474), .B(n_490), .Y(n_569) );
AND2x4_ASAP7_75t_L g605 ( .A(n_474), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g619 ( .A(n_474), .B(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g536 ( .A(n_475), .Y(n_536) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_475), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_SL g563 ( .A1(n_481), .A2(n_536), .B(n_564), .C(n_568), .Y(n_563) );
AND2x2_ASAP7_75t_L g584 ( .A(n_481), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_481), .B(n_536), .Y(n_724) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_490), .Y(n_481) );
INVx2_ASAP7_75t_L g604 ( .A(n_482), .Y(n_604) );
BUFx3_ASAP7_75t_L g620 ( .A(n_482), .Y(n_620) );
INVxp67_ASAP7_75t_L g624 ( .A(n_482), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_488), .Y(n_483) );
INVx2_ASAP7_75t_L g603 ( .A(n_490), .Y(n_603) );
AND2x2_ASAP7_75t_L g609 ( .A(n_490), .B(n_582), .Y(n_609) );
AND2x2_ASAP7_75t_L g635 ( .A(n_490), .B(n_604), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_492), .B(n_496), .Y(n_491) );
AOI211xp5_ASAP7_75t_L g632 ( .A1(n_498), .A2(n_633), .B(n_636), .C(n_646), .Y(n_632) );
AND2x2_ASAP7_75t_SL g498 ( .A(n_499), .B(n_516), .Y(n_498) );
OAI321xp33_ASAP7_75t_L g607 ( .A1(n_499), .A2(n_555), .A3(n_608), .B1(n_610), .B2(n_611), .C(n_613), .Y(n_607) );
AND2x2_ASAP7_75t_L g728 ( .A(n_499), .B(n_703), .Y(n_728) );
INVx1_ASAP7_75t_L g731 ( .A(n_499), .Y(n_731) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_508), .Y(n_499) );
INVx5_ASAP7_75t_L g553 ( .A(n_500), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_500), .B(n_567), .Y(n_566) );
NOR2x1_ASAP7_75t_SL g598 ( .A(n_500), .B(n_599), .Y(n_598) );
BUFx2_ASAP7_75t_L g643 ( .A(n_500), .Y(n_643) );
AND2x2_ASAP7_75t_L g745 ( .A(n_500), .B(n_517), .Y(n_745) );
OR2x6_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
AND2x2_ASAP7_75t_L g552 ( .A(n_508), .B(n_553), .Y(n_552) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_508), .Y(n_562) );
INVx4_ASAP7_75t_L g567 ( .A(n_508), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_514), .Y(n_509) );
INVx1_ASAP7_75t_L g610 ( .A(n_516), .Y(n_610) );
A2O1A1Ixp33_ASAP7_75t_R g713 ( .A1(n_516), .A2(n_552), .B(n_584), .C(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g733 ( .A(n_516), .B(n_558), .Y(n_733) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_524), .Y(n_516) );
INVx1_ASAP7_75t_L g551 ( .A(n_517), .Y(n_551) );
INVx2_ASAP7_75t_L g557 ( .A(n_517), .Y(n_557) );
OR2x2_ASAP7_75t_L g576 ( .A(n_517), .B(n_567), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_517), .B(n_599), .Y(n_645) );
BUFx3_ASAP7_75t_L g652 ( .A(n_517), .Y(n_652) );
INVx1_ASAP7_75t_L g615 ( .A(n_524), .Y(n_615) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_524), .Y(n_628) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g561 ( .A(n_525), .Y(n_561) );
INVx1_ASAP7_75t_L g670 ( .A(n_525), .Y(n_670) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B(n_533), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_526), .B(n_534), .Y(n_533) );
AO21x2_ASAP7_75t_L g599 ( .A1(n_526), .A2(n_527), .B(n_533), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_532), .Y(n_527) );
AND2x2_ASAP7_75t_L g571 ( .A(n_535), .B(n_572), .Y(n_571) );
OAI31xp33_ASAP7_75t_L g722 ( .A1(n_535), .A2(n_723), .A3(n_725), .B(n_728), .Y(n_722) );
INVx1_ASAP7_75t_SL g740 ( .A(n_535), .Y(n_740) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
AOI21xp33_ASAP7_75t_L g554 ( .A1(n_536), .A2(n_555), .B(n_563), .Y(n_554) );
NAND2x1_ASAP7_75t_L g634 ( .A(n_536), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g663 ( .A(n_536), .Y(n_663) );
INVx2_ASAP7_75t_L g612 ( .A(n_537), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_537), .B(n_595), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_537), .B(n_594), .Y(n_704) );
NOR2xp33_ASAP7_75t_SL g712 ( .A(n_537), .B(n_663), .Y(n_712) );
AND2x4_ASAP7_75t_L g537 ( .A(n_538), .B(n_549), .Y(n_537) );
AND2x2_ASAP7_75t_SL g581 ( .A(n_538), .B(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g592 ( .A(n_538), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g621 ( .A(n_538), .B(n_603), .Y(n_621) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g585 ( .A(n_539), .Y(n_585) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g606 ( .A(n_540), .Y(n_606) );
OAI21x1_ASAP7_75t_SL g540 ( .A1(n_541), .A2(n_543), .B(n_547), .Y(n_540) );
INVx1_ASAP7_75t_L g548 ( .A(n_542), .Y(n_548) );
INVx2_ASAP7_75t_L g593 ( .A(n_549), .Y(n_593) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_549), .Y(n_653) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g589 ( .A(n_551), .Y(n_589) );
AND2x2_ASAP7_75t_L g668 ( .A(n_551), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g579 ( .A(n_552), .B(n_573), .Y(n_579) );
INVx2_ASAP7_75t_SL g627 ( .A(n_552), .Y(n_627) );
INVx4_ASAP7_75t_L g558 ( .A(n_553), .Y(n_558) );
AND2x2_ASAP7_75t_L g656 ( .A(n_553), .B(n_599), .Y(n_656) );
AND2x2_ASAP7_75t_SL g674 ( .A(n_553), .B(n_669), .Y(n_674) );
NAND2x1p5_ASAP7_75t_L g691 ( .A(n_553), .B(n_567), .Y(n_691) );
INVx1_ASAP7_75t_L g697 ( .A(n_555), .Y(n_697) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_559), .Y(n_555) );
INVx1_ASAP7_75t_L g616 ( .A(n_556), .Y(n_616) );
OR2x2_ASAP7_75t_L g629 ( .A(n_556), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
OR2x2_ASAP7_75t_L g681 ( .A(n_557), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g711 ( .A(n_557), .B(n_599), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_558), .B(n_561), .Y(n_587) );
AND2x2_ASAP7_75t_L g679 ( .A(n_558), .B(n_669), .Y(n_679) );
AND2x4_ASAP7_75t_L g741 ( .A(n_558), .B(n_620), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
INVx2_ASAP7_75t_L g565 ( .A(n_560), .Y(n_565) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NOR2xp67_ASAP7_75t_SL g564 ( .A(n_565), .B(n_566), .Y(n_564) );
OAI322xp33_ASAP7_75t_SL g577 ( .A1(n_565), .A2(n_578), .A3(n_580), .B1(n_583), .B2(n_586), .C1(n_588), .C2(n_590), .Y(n_577) );
INVx1_ASAP7_75t_L g735 ( .A(n_565), .Y(n_735) );
OR2x2_ASAP7_75t_L g588 ( .A(n_566), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g614 ( .A(n_567), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_567), .B(n_615), .Y(n_630) );
INVx2_ASAP7_75t_L g657 ( .A(n_567), .Y(n_657) );
AND2x4_ASAP7_75t_L g669 ( .A(n_567), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_SL g672 ( .A(n_569), .B(n_585), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_575), .B(n_577), .Y(n_570) );
AND2x2_ASAP7_75t_L g638 ( .A(n_572), .B(n_605), .Y(n_638) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_573), .B(n_727), .Y(n_726) );
BUFx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g596 ( .A(n_574), .Y(n_596) );
AND2x4_ASAP7_75t_SL g678 ( .A(n_574), .B(n_593), .Y(n_678) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g586 ( .A(n_576), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_579), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g714 ( .A(n_581), .B(n_678), .Y(n_714) );
NOR4xp25_ASAP7_75t_L g718 ( .A(n_581), .B(n_595), .C(n_635), .D(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g595 ( .A(n_582), .B(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g631 ( .A(n_582), .B(n_606), .Y(n_631) );
AND2x4_ASAP7_75t_L g695 ( .A(n_582), .B(n_606), .Y(n_695) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_585), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_594), .Y(n_591) );
OR2x2_ASAP7_75t_L g684 ( .A(n_592), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g738 ( .A(n_592), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_593), .B(n_605), .Y(n_639) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
AOI211xp5_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_600), .B(n_607), .C(n_622), .Y(n_597) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_605), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_603), .B(n_606), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_604), .B(n_609), .Y(n_608) );
BUFx2_ASAP7_75t_L g686 ( .A(n_604), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_605), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g701 ( .A(n_605), .Y(n_701) );
OAI21xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .B(n_617), .Y(n_613) );
AND2x4_ASAP7_75t_L g650 ( .A(n_614), .B(n_651), .Y(n_650) );
AND2x4_ASAP7_75t_L g744 ( .A(n_614), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
INVx1_ASAP7_75t_SL g648 ( .A(n_620), .Y(n_648) );
AND2x2_ASAP7_75t_L g707 ( .A(n_621), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g721 ( .A(n_621), .Y(n_721) );
O2A1O1Ixp33_ASAP7_75t_SL g622 ( .A1(n_623), .A2(n_625), .B(n_629), .C(n_631), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_623), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g699 ( .A(n_624), .B(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g720 ( .A(n_624), .B(n_721), .Y(n_720) );
INVxp67_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
OR2x2_ASAP7_75t_L g709 ( .A(n_627), .B(n_651), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_630), .A2(n_637), .B1(n_639), .B2(n_640), .Y(n_636) );
INVx1_ASAP7_75t_SL g727 ( .A(n_631), .Y(n_727) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVxp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_642), .B(n_651), .Y(n_693) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVxp67_ASAP7_75t_SL g703 ( .A(n_645), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B1(n_653), .B2(n_654), .Y(n_646) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI21xp5_ASAP7_75t_SL g660 ( .A1(n_651), .A2(n_661), .B(n_664), .Y(n_660) );
AND2x2_ASAP7_75t_L g689 ( .A(n_651), .B(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND3x2_ASAP7_75t_L g655 ( .A(n_652), .B(n_656), .C(n_657), .Y(n_655) );
AND2x2_ASAP7_75t_L g717 ( .A(n_652), .B(n_674), .Y(n_717) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g702 ( .A(n_657), .B(n_703), .Y(n_702) );
NOR2xp67_ASAP7_75t_L g658 ( .A(n_659), .B(n_715), .Y(n_658) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_660), .B(n_675), .C(n_696), .D(n_713), .Y(n_659) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_667), .B1(n_671), .B2(n_673), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_667), .A2(n_681), .B1(n_701), .B2(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g682 ( .A(n_669), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g742 ( .A1(n_671), .A2(n_694), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx3_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_679), .B1(n_680), .B2(n_683), .C(n_687), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_692), .B1(n_693), .B2(n_694), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_690), .B(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_690), .B(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B1(n_702), .B2(n_704), .C(n_705), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_699), .B(n_701), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_709), .B1(n_710), .B2(n_712), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI211xp5_ASAP7_75t_SL g730 ( .A1(n_711), .A2(n_731), .B(n_732), .C(n_734), .Y(n_730) );
OAI211xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_718), .B(n_722), .C(n_729), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_736), .B1(n_739), .B2(n_741), .C(n_742), .Y(n_729) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
CKINVDCx5p33_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
CKINVDCx11_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
INVx3_ASAP7_75t_SL g753 ( .A(n_749), .Y(n_753) );
CKINVDCx5p33_ASAP7_75t_R g749 ( .A(n_750), .Y(n_749) );
CKINVDCx6p67_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx3_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
endmodule