module real_jpeg_32985_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_0),
.Y(n_116)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_0),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_1),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_87),
.Y(n_92)
);

AND2x4_ASAP7_75t_L g143 ( 
.A(n_1),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_2),
.B(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_3),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_5),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_6),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_6),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_7),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_7),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_7),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_7),
.B(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_7),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_8),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_8),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_8),
.B(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_9),
.Y(n_146)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_9),
.Y(n_190)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_10),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_11),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_11),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_11),
.B(n_121),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_11),
.B(n_187),
.Y(n_186)
);

NAND2x1_ASAP7_75t_L g201 ( 
.A(n_11),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_11),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_11),
.B(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_12),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_13),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_13),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_13),
.B(n_111),
.Y(n_110)
);

AND2x4_ASAP7_75t_SL g183 ( 
.A(n_13),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_13),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_13),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_13),
.B(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_14),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_14),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_15),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_15),
.B(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_15),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_15),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_15),
.B(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_169),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_167),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

NOR2xp67_ASAP7_75t_L g168 ( 
.A(n_19),
.B(n_106),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_68),
.C(n_89),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_20),
.B(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_40),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_22),
.B(n_41),
.C(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_29),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_24),
.B(n_30),
.C(n_39),
.Y(n_162)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_27),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_33),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_33),
.Y(n_204)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_36),
.Y(n_184)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_36),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_51),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_46),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_42),
.B(n_46),
.Y(n_160)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_58),
.C(n_62),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_52),
.B(n_58),
.C(n_62),
.Y(n_165)
);

XNOR2x1_ASAP7_75t_L g247 ( 
.A(n_52),
.B(n_62),
.Y(n_247)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

XNOR2x1_ASAP7_75t_L g246 ( 
.A(n_58),
.B(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_68),
.A2(n_69),
.B1(n_89),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_70),
.B(n_83),
.C(n_88),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_71),
.A2(n_73),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_71),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g182 ( 
.A(n_72),
.Y(n_182)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_75),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_83),
.B1(n_84),
.B2(n_88),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_89),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_97),
.C(n_103),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_90),
.B(n_97),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_92),
.B(n_93),
.Y(n_196)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_103),
.B(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_138),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_137),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_119),
.B1(n_135),
.B2(n_136),
.Y(n_108)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_114),
.B(n_117),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_114),
.Y(n_118)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_116),
.Y(n_216)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_126),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_138)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_158),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_153),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_147),
.B2(n_148),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_156),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_251),
.B(n_256),
.Y(n_170)
);

OAI21x1_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_239),
.B(n_250),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_207),
.B(n_238),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_191),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_174),
.B(n_191),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_183),
.C(n_185),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_175),
.A2(n_176),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_180),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_183),
.A2(n_185),
.B1(n_186),
.B2(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_183),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_197),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_196),
.C(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_201),
.C(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_231),
.B(n_237),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_220),
.B(n_230),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_217),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_217),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_214),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_225),
.Y(n_220)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_233),
.Y(n_237)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_242),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_248),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_246),
.C(n_248),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_255),
.Y(n_251)
);

NOR2xp67_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_255),
.Y(n_256)
);


endmodule