module fake_netlist_5_1035_n_2194 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2194);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2194;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_696;
wire n_550;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_604;
wire n_314;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_2033;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1982;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_2176;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2131;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1865;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_328;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_2135;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g219 ( 
.A(n_147),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_68),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_190),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_62),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_89),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_218),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_122),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_111),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_194),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_54),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_43),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_1),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_82),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_182),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_28),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_1),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_132),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_110),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_4),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_167),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_155),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_193),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_146),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_126),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_49),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_35),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_104),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_160),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_137),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_119),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_78),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_98),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_39),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_157),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_14),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_87),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_130),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_65),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_29),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_127),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_10),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_206),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_9),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_118),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_154),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_144),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_185),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_59),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_44),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_56),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_76),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_33),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_57),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_168),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_38),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_125),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_181),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_213),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_80),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_10),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_48),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_28),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_107),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_21),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_19),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_63),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_174),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_21),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_134),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_42),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_170),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_73),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_183),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_179),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_150),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_162),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_216),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_5),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_79),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_2),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_5),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_141),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_62),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_69),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_96),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_43),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_72),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_133),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_208),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_156),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_211),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_201),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_38),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_18),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_142),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_145),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_59),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_97),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_171),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_8),
.Y(n_319)
);

BUFx10_ASAP7_75t_L g320 ( 
.A(n_8),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_72),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_120),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_116),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_103),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_77),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_7),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_189),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_71),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_60),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_31),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_165),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_114),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_23),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_128),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_151),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_166),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_67),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_124),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_169),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_51),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_42),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_203),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_198),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_85),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_100),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_178),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_55),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_197),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_207),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_139),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_48),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_53),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_54),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_70),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_2),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_123),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_56),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_9),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_217),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_26),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_44),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_158),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_18),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_52),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_16),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_88),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_175),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_30),
.Y(n_368)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_209),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_101),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_94),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_52),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_64),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_192),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_200),
.Y(n_375)
);

INVx4_ASAP7_75t_R g376 ( 
.A(n_83),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_30),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_77),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_15),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_60),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_112),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_180),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_84),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_93),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_41),
.Y(n_385)
);

BUFx2_ASAP7_75t_SL g386 ( 
.A(n_41),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_26),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_65),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_34),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_131),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_176),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_74),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_66),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_91),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_163),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_53),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_69),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_105),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_129),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_108),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_14),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_204),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_64),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_68),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_0),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_49),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_58),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_57),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_109),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_22),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_81),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_73),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_32),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_149),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_29),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_136),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_50),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_115),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_16),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_24),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_95),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_47),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_195),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_143),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_212),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_33),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_35),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_76),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_23),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_117),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_22),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_71),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_7),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_12),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_223),
.B(n_3),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_264),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_221),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_234),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_234),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_224),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_263),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_234),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_234),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_234),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_227),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_265),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_307),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_268),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_310),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_228),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_362),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_233),
.Y(n_452)
);

NOR2xp67_ASAP7_75t_L g453 ( 
.A(n_389),
.B(n_3),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_268),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_223),
.B(n_4),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_287),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_268),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_414),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_236),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_389),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_424),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_237),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_264),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_268),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_239),
.Y(n_465)
);

NOR2xp67_ASAP7_75t_L g466 ( 
.A(n_389),
.B(n_6),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_369),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_268),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_410),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_313),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_382),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_397),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_243),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_L g474 ( 
.A(n_262),
.B(n_6),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_313),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_246),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_313),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_313),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_277),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_250),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_251),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_226),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_255),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_313),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_283),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_261),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_283),
.Y(n_487)
);

INVxp33_ASAP7_75t_L g488 ( 
.A(n_364),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_341),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_273),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_341),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_357),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_357),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_397),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_276),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_278),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_293),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_220),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_220),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_230),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_295),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_296),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g503 ( 
.A(n_297),
.B(n_11),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_230),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_320),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_238),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_308),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_284),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_238),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_309),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_311),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_258),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_258),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_318),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_272),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_272),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_274),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_323),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_334),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_229),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_274),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_231),
.Y(n_522)
);

CKINVDCx14_ASAP7_75t_R g523 ( 
.A(n_277),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_219),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_335),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_279),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_279),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_320),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_303),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_303),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_338),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_305),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_305),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_320),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_306),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_306),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_324),
.B(n_11),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_324),
.B(n_12),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_342),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_390),
.B(n_13),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_R g541 ( 
.A(n_343),
.B(n_86),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_329),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_R g543 ( 
.A(n_346),
.B(n_90),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_329),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_226),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_226),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_219),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_333),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_333),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_337),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_441),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_438),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_478),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_456),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_436),
.B(n_390),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_446),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_438),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_437),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_453),
.B(n_232),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_478),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_439),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_R g562 ( 
.A(n_465),
.B(n_348),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_439),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_510),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_435),
.A2(n_244),
.B1(n_270),
.B2(n_222),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_447),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_436),
.Y(n_567)
);

AND3x1_ASAP7_75t_L g568 ( 
.A(n_455),
.B(n_312),
.C(n_297),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_442),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_469),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_440),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_510),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_443),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_449),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_445),
.B(n_232),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_443),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_444),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_450),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_444),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_448),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_448),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_510),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_454),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_520),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_454),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_452),
.B(n_459),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_457),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_510),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_510),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_462),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_505),
.B(n_259),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_457),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_464),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_464),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_476),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_468),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_468),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_470),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_451),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_470),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_475),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_R g602 ( 
.A(n_467),
.B(n_349),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_475),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_477),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_477),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_484),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_458),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_480),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_484),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_489),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_460),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_463),
.B(n_479),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_463),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_489),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_498),
.Y(n_615)
);

CKINVDCx16_ASAP7_75t_R g616 ( 
.A(n_461),
.Y(n_616)
);

NAND2xp33_ASAP7_75t_R g617 ( 
.A(n_481),
.B(n_483),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_498),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_471),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_486),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_524),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_495),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_499),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_R g624 ( 
.A(n_523),
.B(n_356),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_473),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_496),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_490),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_508),
.B(n_284),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_499),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_500),
.Y(n_630)
);

AND2x6_ASAP7_75t_L g631 ( 
.A(n_460),
.B(n_309),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_500),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_524),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_497),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_501),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_R g636 ( 
.A(n_507),
.B(n_359),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_547),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_547),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_504),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_485),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_485),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_504),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_502),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_553),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_615),
.Y(n_645)
);

NOR2x1p5_ASAP7_75t_L g646 ( 
.A(n_558),
.B(n_482),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_567),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_559),
.B(n_511),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_553),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_567),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_615),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_559),
.B(n_538),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_559),
.B(n_514),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_618),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_559),
.B(n_518),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_575),
.B(n_568),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_564),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_618),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_631),
.B(n_309),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_625),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_564),
.Y(n_661)
);

AND2x6_ASAP7_75t_L g662 ( 
.A(n_555),
.B(n_225),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_560),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_612),
.B(n_519),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_623),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_564),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_612),
.B(n_525),
.Y(n_667)
);

BUFx10_ASAP7_75t_L g668 ( 
.A(n_571),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_560),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_624),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_564),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_586),
.B(n_531),
.Y(n_672)
);

OAI21xp33_ASAP7_75t_SL g673 ( 
.A1(n_555),
.A2(n_540),
.B(n_537),
.Y(n_673)
);

AND2x6_ASAP7_75t_SL g674 ( 
.A(n_628),
.B(n_337),
.Y(n_674)
);

AND2x2_ASAP7_75t_SL g675 ( 
.A(n_565),
.B(n_253),
.Y(n_675)
);

INVxp67_ASAP7_75t_L g676 ( 
.A(n_628),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_613),
.Y(n_677)
);

BUFx4f_ASAP7_75t_L g678 ( 
.A(n_637),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_613),
.B(n_253),
.Y(n_679)
);

AND2x2_ASAP7_75t_SL g680 ( 
.A(n_565),
.B(n_286),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_623),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_584),
.B(n_522),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_578),
.B(n_539),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_590),
.B(n_494),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_564),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_629),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_629),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_630),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_563),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_637),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_630),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_589),
.B(n_247),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_636),
.B(n_286),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_632),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_632),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_564),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_563),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_576),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_595),
.B(n_288),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_639),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_576),
.Y(n_701)
);

BUFx10_ASAP7_75t_L g702 ( 
.A(n_608),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_639),
.Y(n_703)
);

AND2x6_ASAP7_75t_L g704 ( 
.A(n_642),
.B(n_225),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_631),
.B(n_309),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_577),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_SL g707 ( 
.A(n_591),
.B(n_312),
.Y(n_707)
);

NOR3xp33_ASAP7_75t_L g708 ( 
.A(n_616),
.B(n_528),
.C(n_534),
.Y(n_708)
);

INVx4_ASAP7_75t_SL g709 ( 
.A(n_631),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_642),
.A2(n_466),
.B1(n_420),
.B2(n_352),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_577),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_611),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_551),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_620),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_622),
.B(n_482),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_552),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_552),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_585),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_556),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_640),
.B(n_240),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_585),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_637),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_557),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_589),
.B(n_545),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_589),
.B(n_545),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_557),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_572),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_597),
.Y(n_728)
);

INVx4_ASAP7_75t_SL g729 ( 
.A(n_631),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_597),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_561),
.B(n_569),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_561),
.B(n_546),
.Y(n_732)
);

INVx4_ASAP7_75t_SL g733 ( 
.A(n_631),
.Y(n_733)
);

INVx4_ASAP7_75t_SL g734 ( 
.A(n_631),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_569),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_554),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_570),
.B(n_472),
.Y(n_737)
);

AND2x6_ASAP7_75t_L g738 ( 
.A(n_611),
.B(n_240),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_637),
.Y(n_739)
);

NAND3xp33_ASAP7_75t_L g740 ( 
.A(n_617),
.B(n_474),
.C(n_508),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_626),
.B(n_288),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_634),
.B(n_546),
.Y(n_742)
);

INVx5_ASAP7_75t_L g743 ( 
.A(n_631),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_573),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_621),
.A2(n_420),
.B1(n_351),
.B2(n_360),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_572),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_SL g747 ( 
.A(n_635),
.B(n_300),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_637),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_643),
.A2(n_292),
.B1(n_331),
.B2(n_256),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_579),
.B(n_580),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_579),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_600),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_580),
.B(n_332),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_640),
.B(n_241),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_600),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_581),
.B(n_344),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_583),
.B(n_395),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_611),
.B(n_350),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_583),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_611),
.Y(n_760)
);

OR2x6_ASAP7_75t_L g761 ( 
.A(n_616),
.B(n_386),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_603),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_621),
.A2(n_351),
.B1(n_360),
.B2(n_352),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_587),
.B(n_488),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_587),
.B(n_409),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_592),
.B(n_366),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_603),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_592),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_611),
.B(n_350),
.Y(n_769)
);

NAND3xp33_ASAP7_75t_L g770 ( 
.A(n_593),
.B(n_503),
.C(n_245),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_637),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_605),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_611),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_605),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_593),
.B(n_367),
.Y(n_775)
);

AND2x2_ASAP7_75t_SL g776 ( 
.A(n_633),
.B(n_374),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_562),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_641),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_602),
.B(n_374),
.Y(n_779)
);

CKINVDCx14_ASAP7_75t_R g780 ( 
.A(n_619),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_594),
.B(n_370),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_594),
.B(n_506),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_610),
.B(n_431),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_596),
.B(n_371),
.Y(n_784)
);

CKINVDCx16_ASAP7_75t_R g785 ( 
.A(n_566),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_641),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_574),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_641),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_610),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_596),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_614),
.B(n_433),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_627),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_598),
.B(n_309),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_614),
.B(n_506),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_633),
.B(n_241),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_638),
.B(n_509),
.Y(n_796)
);

INVx4_ASAP7_75t_SL g797 ( 
.A(n_572),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_689),
.Y(n_798)
);

O2A1O1Ixp5_ASAP7_75t_L g799 ( 
.A1(n_652),
.A2(n_656),
.B(n_769),
.C(n_758),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_645),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_776),
.B(n_638),
.Y(n_801)
);

OAI221xp5_ASAP7_75t_L g802 ( 
.A1(n_673),
.A2(n_289),
.B1(n_429),
.B2(n_379),
.C(n_373),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_676),
.B(n_509),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_776),
.B(n_601),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_644),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_656),
.A2(n_249),
.B1(n_384),
.B2(n_383),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_652),
.B(n_601),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_699),
.A2(n_365),
.B(n_368),
.C(n_363),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_644),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_667),
.B(n_606),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_783),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_667),
.B(n_651),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_654),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_658),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_665),
.B(n_606),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_649),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_664),
.B(n_599),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_662),
.A2(n_394),
.B1(n_400),
.B2(n_399),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_L g819 ( 
.A(n_662),
.B(n_375),
.Y(n_819)
);

NAND3xp33_ASAP7_75t_L g820 ( 
.A(n_740),
.B(n_252),
.C(n_235),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_681),
.B(n_609),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_791),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_684),
.B(n_607),
.Y(n_823)
);

INVx4_ASAP7_75t_L g824 ( 
.A(n_678),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_648),
.B(n_375),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_686),
.B(n_609),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_649),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_662),
.A2(n_680),
.B1(n_675),
.B2(n_655),
.Y(n_828)
);

BUFx12f_ASAP7_75t_L g829 ( 
.A(n_668),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_684),
.B(n_254),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_737),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_683),
.B(n_257),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_662),
.A2(n_416),
.B1(n_430),
.B2(n_421),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_699),
.A2(n_388),
.B(n_373),
.C(n_368),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_687),
.B(n_604),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_688),
.B(n_604),
.Y(n_836)
);

INVxp33_ASAP7_75t_L g837 ( 
.A(n_764),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_691),
.Y(n_838)
);

AOI22x1_ASAP7_75t_L g839 ( 
.A1(n_694),
.A2(n_402),
.B1(n_345),
.B2(n_339),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_695),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_700),
.B(n_604),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_683),
.B(n_260),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_672),
.B(n_267),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_653),
.B(n_269),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_703),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_675),
.B(n_402),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_662),
.B(n_716),
.Y(n_847)
);

NOR2xp67_ASAP7_75t_L g848 ( 
.A(n_777),
.B(n_736),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_796),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_794),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_680),
.A2(n_322),
.B1(n_425),
.B2(n_418),
.Y(n_851)
);

XNOR2xp5_ASAP7_75t_L g852 ( 
.A(n_713),
.B(n_719),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_715),
.B(n_271),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_764),
.B(n_281),
.C(n_280),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_663),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_717),
.B(n_604),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_689),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_749),
.B(n_282),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_723),
.B(n_641),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_663),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_715),
.B(n_285),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_742),
.B(n_741),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_678),
.A2(n_582),
.B(n_572),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_742),
.B(n_299),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_726),
.B(n_641),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_735),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_669),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_657),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_677),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_743),
.B(n_423),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_677),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_R g872 ( 
.A(n_780),
.B(n_415),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_669),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_L g874 ( 
.A(n_765),
.B(n_741),
.C(n_693),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_704),
.A2(n_242),
.B1(n_248),
.B2(n_266),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_647),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_693),
.A2(n_294),
.B1(n_290),
.B2(n_275),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_704),
.A2(n_242),
.B1(n_248),
.B2(n_266),
.Y(n_878)
);

INVxp67_ASAP7_75t_L g879 ( 
.A(n_682),
.Y(n_879)
);

NAND3xp33_ASAP7_75t_L g880 ( 
.A(n_765),
.B(n_316),
.C(n_302),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_743),
.B(n_275),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_744),
.B(n_641),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_761),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_647),
.B(n_650),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_697),
.Y(n_885)
);

BUFx8_ASAP7_75t_L g886 ( 
.A(n_670),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_650),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_732),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_751),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_779),
.B(n_319),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_697),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_743),
.B(n_294),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_759),
.B(n_768),
.Y(n_893)
);

O2A1O1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_679),
.A2(n_365),
.B(n_363),
.C(n_379),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_779),
.B(n_321),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_747),
.B(n_325),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_790),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_698),
.Y(n_898)
);

AND2x6_ASAP7_75t_SL g899 ( 
.A(n_761),
.B(n_388),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_789),
.B(n_298),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_698),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_766),
.B(n_301),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_778),
.B(n_301),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_701),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_701),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_778),
.B(n_314),
.Y(n_906)
);

OAI22xp33_ASAP7_75t_L g907 ( 
.A1(n_753),
.A2(n_336),
.B1(n_327),
.B2(n_322),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_706),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_720),
.B(n_512),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_761),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_706),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_786),
.B(n_314),
.Y(n_912)
);

CKINVDCx11_ASAP7_75t_R g913 ( 
.A(n_668),
.Y(n_913)
);

OAI221xp5_ASAP7_75t_L g914 ( 
.A1(n_710),
.A2(n_745),
.B1(n_763),
.B2(n_756),
.C(n_757),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_775),
.B(n_315),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_711),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_711),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_704),
.A2(n_398),
.B1(n_327),
.B2(n_317),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_786),
.B(n_788),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_781),
.B(n_315),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_784),
.B(n_707),
.Y(n_921)
);

CKINVDCx16_ASAP7_75t_R g922 ( 
.A(n_785),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_718),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_704),
.A2(n_418),
.B1(n_317),
.B2(n_425),
.Y(n_924)
);

OAI21xp33_ASAP7_75t_L g925 ( 
.A1(n_710),
.A2(n_291),
.B(n_393),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_718),
.Y(n_926)
);

INVxp67_ASAP7_75t_L g927 ( 
.A(n_707),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_721),
.Y(n_928)
);

NOR2xp67_ASAP7_75t_L g929 ( 
.A(n_770),
.B(n_92),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_788),
.B(n_381),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_731),
.B(n_381),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_750),
.B(n_391),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_704),
.A2(n_411),
.B1(n_398),
.B2(n_391),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_720),
.A2(n_411),
.B1(n_386),
.B2(n_291),
.Y(n_934)
);

NAND3xp33_ASAP7_75t_SL g935 ( 
.A(n_708),
.B(n_419),
.C(n_328),
.Y(n_935)
);

AND2x6_ASAP7_75t_SL g936 ( 
.A(n_713),
.B(n_393),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_795),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_721),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_724),
.B(n_541),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_720),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_725),
.B(n_326),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_754),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_660),
.B(n_330),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_792),
.B(n_340),
.Y(n_944)
);

AND2x2_ASAP7_75t_SL g945 ( 
.A(n_659),
.B(n_405),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_679),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_754),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_754),
.B(n_512),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_690),
.B(n_572),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_690),
.B(n_572),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_722),
.B(n_582),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_722),
.B(n_582),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_782),
.B(n_513),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_787),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_739),
.B(n_582),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_728),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_739),
.B(n_582),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_748),
.B(n_582),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_748),
.B(n_588),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_728),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_674),
.B(n_347),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_771),
.B(n_588),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_646),
.A2(n_259),
.B1(n_304),
.B2(n_385),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_953),
.B(n_782),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_891),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_799),
.A2(n_769),
.B(n_758),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_953),
.B(n_730),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_819),
.A2(n_760),
.B(n_712),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_888),
.B(n_752),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_819),
.A2(n_847),
.B(n_949),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_950),
.A2(n_952),
.B(n_951),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_851),
.A2(n_763),
.B1(n_745),
.B2(n_417),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_955),
.A2(n_958),
.B(n_957),
.Y(n_973)
);

AO21x1_ASAP7_75t_L g974 ( 
.A1(n_846),
.A2(n_692),
.B(n_793),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_829),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_888),
.B(n_752),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_846),
.A2(n_762),
.B(n_755),
.C(n_774),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_811),
.B(n_513),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_802),
.A2(n_762),
.B1(n_755),
.B2(n_767),
.Y(n_979)
);

AND2x6_ASAP7_75t_SL g980 ( 
.A(n_961),
.B(n_405),
.Y(n_980)
);

CKINVDCx10_ASAP7_75t_R g981 ( 
.A(n_922),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_SL g982 ( 
.A1(n_862),
.A2(n_830),
.B1(n_842),
.B2(n_832),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_837),
.B(n_879),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_959),
.A2(n_760),
.B(n_712),
.Y(n_984)
);

AND2x4_ASAP7_75t_SL g985 ( 
.A(n_869),
.B(n_702),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_831),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_962),
.A2(n_773),
.B(n_771),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_837),
.B(n_702),
.Y(n_988)
);

CKINVDCx10_ASAP7_75t_R g989 ( 
.A(n_852),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_810),
.B(n_773),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_874),
.A2(n_772),
.B(n_767),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_868),
.A2(n_661),
.B(n_657),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_868),
.A2(n_824),
.B(n_807),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_812),
.B(n_772),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_L g995 ( 
.A1(n_914),
.A2(n_774),
.B1(n_738),
.B2(n_304),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_804),
.A2(n_877),
.B(n_858),
.C(n_907),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_843),
.B(n_671),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_868),
.A2(n_661),
.B(n_657),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_801),
.A2(n_696),
.B(n_671),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_853),
.B(n_696),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_861),
.B(n_746),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_824),
.A2(n_661),
.B(n_657),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_871),
.Y(n_1003)
);

O2A1O1Ixp5_ASAP7_75t_L g1004 ( 
.A1(n_825),
.A2(n_746),
.B(n_432),
.C(n_434),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_811),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_891),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_824),
.A2(n_666),
.B(n_661),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_822),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_946),
.A2(n_705),
.B(n_659),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_919),
.A2(n_685),
.B(n_666),
.Y(n_1010)
);

BUFx4f_ASAP7_75t_L g1011 ( 
.A(n_829),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_805),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_822),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_823),
.B(n_515),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_864),
.B(n_666),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_919),
.A2(n_685),
.B(n_666),
.Y(n_1016)
);

BUFx8_ASAP7_75t_L g1017 ( 
.A(n_803),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_954),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_800),
.B(n_727),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_893),
.A2(n_588),
.B(n_793),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_835),
.A2(n_841),
.B(n_836),
.Y(n_1021)
);

NAND3xp33_ASAP7_75t_L g1022 ( 
.A(n_896),
.B(n_780),
.C(n_361),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_828),
.B(n_714),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_937),
.A2(n_588),
.B(n_797),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_813),
.B(n_738),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_814),
.B(n_738),
.Y(n_1026)
);

AO21x1_ASAP7_75t_L g1027 ( 
.A1(n_890),
.A2(n_434),
.B(n_432),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_848),
.B(n_714),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_871),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_940),
.A2(n_738),
.B1(n_259),
.B2(n_304),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_817),
.B(n_719),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_809),
.Y(n_1032)
);

AO21x1_ASAP7_75t_L g1033 ( 
.A1(n_895),
.A2(n_428),
.B(n_412),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_942),
.A2(n_588),
.B(n_797),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_947),
.A2(n_738),
.B1(n_543),
.B2(n_417),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_859),
.A2(n_588),
.B(n_797),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_865),
.A2(n_376),
.B(n_733),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_798),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_850),
.B(n_709),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_876),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_844),
.B(n_709),
.Y(n_1041)
);

NAND3xp33_ASAP7_75t_L g1042 ( 
.A(n_943),
.B(n_380),
.C(n_378),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_856),
.A2(n_530),
.B(n_515),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_809),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_909),
.B(n_729),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_SL g1046 ( 
.A(n_954),
.B(n_353),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_798),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_921),
.B(n_849),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_882),
.A2(n_939),
.B(n_884),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_876),
.B(n_887),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_857),
.A2(n_426),
.B(n_517),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_939),
.A2(n_734),
.B(n_733),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_909),
.B(n_729),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_902),
.A2(n_354),
.B(n_355),
.C(n_358),
.Y(n_1054)
);

AND2x4_ASAP7_75t_SL g1055 ( 
.A(n_883),
.B(n_516),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_915),
.A2(n_734),
.B(n_733),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_948),
.B(n_729),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_R g1058 ( 
.A(n_852),
.B(n_372),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_887),
.B(n_941),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_820),
.A2(n_734),
.B1(n_377),
.B2(n_401),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_816),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_806),
.B(n_387),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_948),
.B(n_392),
.Y(n_1063)
);

INVxp67_ASAP7_75t_L g1064 ( 
.A(n_944),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_920),
.A2(n_396),
.B(n_403),
.C(n_404),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_857),
.A2(n_550),
.B(n_549),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_911),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_815),
.A2(n_548),
.B(n_544),
.Y(n_1068)
);

AOI21x1_ASAP7_75t_L g1069 ( 
.A1(n_863),
.A2(n_487),
.B(n_491),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_931),
.B(n_406),
.Y(n_1070)
);

AOI21x1_ASAP7_75t_L g1071 ( 
.A1(n_932),
.A2(n_487),
.B(n_491),
.Y(n_1071)
);

INVxp67_ASAP7_75t_L g1072 ( 
.A(n_854),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_SL g1073 ( 
.A(n_886),
.B(n_407),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_821),
.A2(n_544),
.B(n_542),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_838),
.B(n_840),
.Y(n_1075)
);

BUFx4f_ASAP7_75t_L g1076 ( 
.A(n_845),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_934),
.A2(n_408),
.B1(n_413),
.B2(n_422),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_826),
.A2(n_542),
.B(n_536),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_880),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_875),
.A2(n_427),
.B1(n_535),
.B2(n_533),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_911),
.A2(n_536),
.B(n_535),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_923),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_872),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_870),
.A2(n_533),
.B(n_532),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_866),
.B(n_516),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_870),
.A2(n_532),
.B(n_530),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_885),
.A2(n_529),
.B(n_527),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_878),
.A2(n_529),
.B1(n_527),
.B2(n_526),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_901),
.A2(n_521),
.B(n_517),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_808),
.A2(n_493),
.B(n_492),
.C(n_17),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_904),
.A2(n_113),
.B(n_214),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_904),
.A2(n_106),
.B(n_210),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_923),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_926),
.A2(n_102),
.B(n_205),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_889),
.B(n_99),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_891),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_R g1097 ( 
.A(n_913),
.B(n_202),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_827),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_897),
.B(n_199),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_928),
.B(n_164),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_918),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_905),
.A2(n_196),
.B(n_191),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_928),
.A2(n_188),
.B(n_187),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_927),
.B(n_19),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_905),
.A2(n_186),
.B(n_184),
.Y(n_1105)
);

OAI21xp33_ASAP7_75t_L g1106 ( 
.A1(n_925),
.A2(n_20),
.B(n_24),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_960),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_924),
.A2(n_20),
.B1(n_25),
.B2(n_27),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_834),
.A2(n_25),
.B(n_27),
.C(n_31),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_818),
.B(n_177),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_898),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_SL g1112 ( 
.A(n_886),
.B(n_173),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_908),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_898),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_908),
.B(n_152),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_910),
.B(n_172),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_916),
.A2(n_161),
.B(n_159),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_833),
.A2(n_929),
.B1(n_935),
.B2(n_930),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_916),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_898),
.Y(n_1120)
);

CKINVDCx8_ASAP7_75t_R g1121 ( 
.A(n_899),
.Y(n_1121)
);

NOR2x1p5_ASAP7_75t_SL g1122 ( 
.A(n_917),
.B(n_148),
.Y(n_1122)
);

BUFx12f_ASAP7_75t_L g1123 ( 
.A(n_913),
.Y(n_1123)
);

BUFx8_ASAP7_75t_L g1124 ( 
.A(n_886),
.Y(n_1124)
);

AOI21x1_ASAP7_75t_L g1125 ( 
.A1(n_881),
.A2(n_153),
.B(n_140),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_900),
.B(n_138),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_903),
.A2(n_32),
.B(n_34),
.C(n_36),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_894),
.A2(n_36),
.B(n_37),
.C(n_39),
.Y(n_1128)
);

NAND2xp33_ASAP7_75t_L g1129 ( 
.A(n_933),
.B(n_135),
.Y(n_1129)
);

AND2x2_ASAP7_75t_SL g1130 ( 
.A(n_945),
.B(n_37),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_917),
.B(n_121),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_938),
.Y(n_1132)
);

AO21x1_ASAP7_75t_L g1133 ( 
.A1(n_903),
.A2(n_40),
.B(n_45),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_938),
.A2(n_40),
.B(n_45),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_945),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_956),
.A2(n_46),
.B(n_47),
.Y(n_1136)
);

INVx1_ASAP7_75t_SL g1137 ( 
.A(n_936),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_956),
.A2(n_46),
.B(n_50),
.Y(n_1138)
);

AO21x1_ASAP7_75t_L g1139 ( 
.A1(n_906),
.A2(n_55),
.B(n_58),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_855),
.A2(n_61),
.B(n_63),
.Y(n_1140)
);

NAND2x1p5_ASAP7_75t_L g1141 ( 
.A(n_1040),
.B(n_860),
.Y(n_1141)
);

OAI22x1_ASAP7_75t_L g1142 ( 
.A1(n_1031),
.A2(n_963),
.B1(n_839),
.B2(n_912),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_1005),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1012),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_1014),
.B(n_855),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_971),
.A2(n_860),
.B(n_873),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_982),
.A2(n_966),
.B(n_970),
.Y(n_1147)
);

AO31x2_ASAP7_75t_L g1148 ( 
.A1(n_974),
.A2(n_873),
.A3(n_867),
.B(n_839),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1015),
.A2(n_892),
.B(n_867),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_964),
.A2(n_973),
.B(n_967),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_1018),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_964),
.B(n_930),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1064),
.B(n_912),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1038),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_967),
.B(n_906),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_1083),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1008),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1017),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_994),
.B(n_892),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1047),
.Y(n_1160)
);

AOI221xp5_ASAP7_75t_SL g1161 ( 
.A1(n_1106),
.A2(n_61),
.B1(n_66),
.B2(n_67),
.C(n_70),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_969),
.B(n_74),
.Y(n_1162)
);

OAI22x1_ASAP7_75t_L g1163 ( 
.A1(n_988),
.A2(n_75),
.B1(n_1104),
.B2(n_1116),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_1040),
.B(n_75),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_969),
.B(n_976),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_987),
.A2(n_984),
.B(n_968),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_L g1167 ( 
.A1(n_1077),
.A2(n_972),
.B1(n_983),
.B2(n_1101),
.C(n_1108),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1075),
.B(n_1070),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_991),
.A2(n_999),
.B(n_1021),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1067),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_978),
.B(n_1063),
.Y(n_1171)
);

AOI21x1_ASAP7_75t_SL g1172 ( 
.A1(n_1099),
.A2(n_1100),
.B(n_1115),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1043),
.A2(n_1016),
.B(n_1010),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_1017),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_993),
.A2(n_1049),
.B(n_1001),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1040),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1000),
.A2(n_997),
.B(n_990),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1055),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1130),
.A2(n_1135),
.B1(n_972),
.B2(n_1134),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_1111),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1063),
.B(n_1013),
.Y(n_1181)
);

AND2x6_ASAP7_75t_L g1182 ( 
.A(n_1135),
.B(n_1045),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1075),
.B(n_1070),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_SL g1184 ( 
.A1(n_1094),
.A2(n_1103),
.B(n_1110),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_986),
.B(n_1085),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1053),
.A2(n_1057),
.B(n_1120),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1082),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1057),
.A2(n_1120),
.B(n_1041),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1027),
.A2(n_1033),
.A3(n_1139),
.B(n_1133),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_976),
.B(n_1048),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1050),
.A2(n_998),
.B(n_992),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1093),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1079),
.B(n_1072),
.Y(n_1193)
);

NOR2x1_ASAP7_75t_L g1194 ( 
.A(n_1022),
.B(n_1028),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1002),
.A2(n_1007),
.B(n_1037),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1085),
.B(n_1135),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1032),
.Y(n_1197)
);

AOI21xp33_ASAP7_75t_L g1198 ( 
.A1(n_996),
.A2(n_1140),
.B(n_1062),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1076),
.A2(n_1023),
.B1(n_1118),
.B2(n_1108),
.Y(n_1199)
);

INVx5_ASAP7_75t_L g1200 ( 
.A(n_1111),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1107),
.B(n_1113),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_1046),
.Y(n_1202)
);

AOI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1100),
.A2(n_1131),
.B(n_1115),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1124),
.Y(n_1204)
);

NAND2x1_ASAP7_75t_L g1205 ( 
.A(n_965),
.B(n_1006),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_985),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1076),
.A2(n_1099),
.B(n_1065),
.C(n_1054),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1101),
.A2(n_995),
.B1(n_979),
.B2(n_1009),
.Y(n_1208)
);

NOR2xp67_ASAP7_75t_L g1209 ( 
.A(n_1042),
.B(n_1060),
.Y(n_1209)
);

AOI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1131),
.A2(n_1069),
.B(n_1036),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1119),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_1003),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_SL g1213 ( 
.A(n_1112),
.B(n_1073),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1003),
.B(n_1029),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1003),
.B(n_1029),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1052),
.A2(n_1019),
.B(n_1039),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1124),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1128),
.A2(n_1138),
.A3(n_1020),
.B(n_1026),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1051),
.B(n_1044),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1132),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1039),
.A2(n_1129),
.B(n_1056),
.Y(n_1221)
);

NOR2x1_ASAP7_75t_SL g1222 ( 
.A(n_1111),
.B(n_1114),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_SL g1223 ( 
.A1(n_977),
.A2(n_1066),
.B(n_1081),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1004),
.A2(n_1061),
.B(n_1098),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1025),
.A2(n_1024),
.B(n_1034),
.Y(n_1225)
);

OAI22x1_ASAP7_75t_L g1226 ( 
.A1(n_1116),
.A2(n_1137),
.B1(n_989),
.B2(n_980),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1029),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_965),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1084),
.A2(n_1086),
.B(n_1136),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1006),
.A2(n_1096),
.B(n_1125),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1058),
.B(n_1077),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1096),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1114),
.A2(n_1095),
.B(n_1035),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1114),
.B(n_1030),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_975),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1011),
.B(n_1068),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1011),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_981),
.B(n_1121),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1122),
.B(n_1126),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1071),
.A2(n_1092),
.B(n_1091),
.Y(n_1240)
);

O2A1O1Ixp5_ASAP7_75t_L g1241 ( 
.A1(n_1102),
.A2(n_1105),
.B(n_1117),
.C(n_1078),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1097),
.B(n_1080),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1088),
.A2(n_1074),
.B(n_1089),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1127),
.A2(n_1090),
.B(n_1087),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_SL g1245 ( 
.A1(n_1109),
.A2(n_1088),
.B(n_1080),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1123),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1015),
.A2(n_824),
.B(n_968),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1015),
.A2(n_824),
.B(n_968),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_982),
.A2(n_799),
.B(n_966),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1003),
.B(n_871),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_982),
.A2(n_862),
.B(n_874),
.C(n_996),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_971),
.A2(n_973),
.B(n_970),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_982),
.B(n_964),
.Y(n_1253)
);

AOI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1015),
.A2(n_1049),
.B(n_1041),
.Y(n_1254)
);

AO21x2_ASAP7_75t_L g1255 ( 
.A1(n_999),
.A2(n_966),
.B(n_1049),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1005),
.Y(n_1256)
);

INVxp67_ASAP7_75t_SL g1257 ( 
.A(n_1040),
.Y(n_1257)
);

NAND2x1_ASAP7_75t_L g1258 ( 
.A(n_1120),
.B(n_868),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_971),
.A2(n_973),
.B(n_970),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1015),
.A2(n_824),
.B(n_968),
.Y(n_1260)
);

OAI21xp33_ASAP7_75t_SL g1261 ( 
.A1(n_964),
.A2(n_1048),
.B(n_1130),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_982),
.B(n_964),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1040),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_971),
.A2(n_973),
.B(n_970),
.Y(n_1264)
);

AOI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1015),
.A2(n_1049),
.B(n_1041),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_982),
.A2(n_799),
.B(n_966),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1015),
.A2(n_824),
.B(n_968),
.Y(n_1267)
);

NAND3xp33_ASAP7_75t_L g1268 ( 
.A(n_982),
.B(n_830),
.C(n_832),
.Y(n_1268)
);

AND2x2_ASAP7_75t_SL g1269 ( 
.A(n_1130),
.B(n_1112),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_982),
.B(n_964),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1017),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_982),
.A2(n_862),
.B1(n_832),
.B2(n_842),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1005),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1040),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1014),
.B(n_660),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_982),
.B(n_964),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1015),
.A2(n_824),
.B(n_968),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_982),
.B(n_964),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1038),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_982),
.B(n_1064),
.Y(n_1280)
);

INVx3_ASAP7_75t_SL g1281 ( 
.A(n_1018),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1003),
.B(n_871),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_982),
.A2(n_964),
.B1(n_851),
.B2(n_1130),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1015),
.A2(n_824),
.B(n_968),
.Y(n_1284)
);

OAI21xp33_ASAP7_75t_L g1285 ( 
.A1(n_982),
.A2(n_830),
.B(n_565),
.Y(n_1285)
);

O2A1O1Ixp5_ASAP7_75t_L g1286 ( 
.A1(n_1059),
.A2(n_862),
.B(n_832),
.C(n_842),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_982),
.B(n_964),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1040),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1014),
.B(n_837),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_971),
.A2(n_973),
.B(n_970),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1015),
.A2(n_824),
.B(n_968),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_983),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_971),
.A2(n_973),
.B(n_970),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_971),
.A2(n_973),
.B(n_970),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_983),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1215),
.B(n_1250),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1154),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1180),
.Y(n_1298)
);

NOR2xp67_ASAP7_75t_L g1299 ( 
.A(n_1202),
.B(n_1275),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1143),
.Y(n_1300)
);

AOI21xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1226),
.A2(n_1285),
.B(n_1163),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1171),
.B(n_1289),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1160),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1215),
.B(n_1250),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1168),
.B(n_1183),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1281),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1253),
.B(n_1270),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_1157),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1272),
.B(n_1193),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1256),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1268),
.A2(n_1269),
.B1(n_1231),
.B2(n_1280),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1170),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1282),
.B(n_1212),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1292),
.B(n_1295),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1187),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1192),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1253),
.B(n_1270),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1273),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1180),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1151),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1227),
.Y(n_1321)
);

INVx3_ASAP7_75t_SL g1322 ( 
.A(n_1237),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1282),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1287),
.B(n_1262),
.Y(n_1324)
);

BUFx8_ASAP7_75t_SL g1325 ( 
.A(n_1217),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1176),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1184),
.A2(n_1260),
.B(n_1267),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1251),
.A2(n_1249),
.B(n_1266),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1287),
.B(n_1276),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1279),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1181),
.B(n_1242),
.Y(n_1331)
);

NAND3xp33_ASAP7_75t_L g1332 ( 
.A(n_1286),
.B(n_1167),
.C(n_1283),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1213),
.B(n_1185),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_1227),
.Y(n_1334)
);

AOI21xp33_ASAP7_75t_L g1335 ( 
.A1(n_1283),
.A2(n_1199),
.B(n_1278),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1277),
.A2(n_1284),
.B(n_1291),
.Y(n_1336)
);

NAND2x1p5_ASAP7_75t_L g1337 ( 
.A(n_1200),
.B(n_1176),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1227),
.Y(n_1338)
);

AOI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1210),
.A2(n_1265),
.B(n_1254),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1198),
.A2(n_1261),
.B(n_1199),
.C(n_1208),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1198),
.A2(n_1208),
.B(n_1179),
.C(n_1209),
.Y(n_1341)
);

OR2x6_ASAP7_75t_L g1342 ( 
.A(n_1237),
.B(n_1196),
.Y(n_1342)
);

O2A1O1Ixp5_ASAP7_75t_L g1343 ( 
.A1(n_1147),
.A2(n_1249),
.B(n_1266),
.C(n_1175),
.Y(n_1343)
);

O2A1O1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1179),
.A2(n_1207),
.B(n_1213),
.C(n_1236),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1153),
.A2(n_1147),
.B(n_1162),
.C(n_1190),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1165),
.A2(n_1145),
.B1(n_1245),
.B2(n_1152),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1177),
.A2(n_1150),
.B(n_1223),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1165),
.A2(n_1190),
.B1(n_1201),
.B2(n_1162),
.Y(n_1348)
);

INVxp67_ASAP7_75t_SL g1349 ( 
.A(n_1263),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1164),
.B(n_1257),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1233),
.A2(n_1244),
.B(n_1243),
.C(n_1169),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1155),
.B(n_1182),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1263),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1263),
.B(n_1274),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1178),
.B(n_1206),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1274),
.Y(n_1356)
);

BUFx12f_ASAP7_75t_L g1357 ( 
.A(n_1237),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1201),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1156),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1252),
.A2(n_1294),
.B(n_1264),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1274),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1211),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1155),
.A2(n_1220),
.B1(n_1219),
.B2(n_1159),
.Y(n_1363)
);

NOR3xp33_ASAP7_75t_L g1364 ( 
.A(n_1194),
.B(n_1238),
.C(n_1234),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1164),
.B(n_1288),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1144),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1206),
.Y(n_1367)
);

AND2x2_ASAP7_75t_SL g1368 ( 
.A(n_1158),
.B(n_1174),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1288),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1214),
.B(n_1200),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1235),
.Y(n_1371)
);

NAND2xp33_ASAP7_75t_L g1372 ( 
.A(n_1182),
.B(n_1142),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1197),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1228),
.Y(n_1374)
);

OAI221xp5_ASAP7_75t_L g1375 ( 
.A1(n_1161),
.A2(n_1159),
.B1(n_1229),
.B2(n_1225),
.C(n_1271),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1232),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1230),
.A2(n_1146),
.B(n_1195),
.Y(n_1377)
);

NAND2x1p5_ASAP7_75t_L g1378 ( 
.A(n_1200),
.B(n_1258),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1182),
.B(n_1186),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1259),
.A2(n_1293),
.B(n_1290),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1141),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1200),
.B(n_1222),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1255),
.A2(n_1221),
.B(n_1191),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1182),
.A2(n_1239),
.B1(n_1141),
.B2(n_1225),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_SL g1385 ( 
.A1(n_1229),
.A2(n_1216),
.B(n_1224),
.C(n_1188),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1239),
.A2(n_1161),
.B1(n_1203),
.B2(n_1224),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1246),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1205),
.B(n_1204),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1149),
.A2(n_1189),
.B1(n_1172),
.B2(n_1218),
.Y(n_1389)
);

AND2x4_ASAP7_75t_SL g1390 ( 
.A(n_1218),
.B(n_1189),
.Y(n_1390)
);

AO22x1_ASAP7_75t_L g1391 ( 
.A1(n_1189),
.A2(n_1218),
.B1(n_1241),
.B2(n_1148),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1148),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1148),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1166),
.A2(n_1173),
.B(n_1240),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1227),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1154),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1215),
.B(n_1250),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1143),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1272),
.A2(n_982),
.B1(n_1283),
.B2(n_1268),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1143),
.Y(n_1400)
);

INVx1_ASAP7_75t_SL g1401 ( 
.A(n_1143),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1230),
.A2(n_1146),
.B(n_1195),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1168),
.B(n_1183),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1176),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1184),
.A2(n_1248),
.B(n_1247),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1285),
.A2(n_982),
.B1(n_1268),
.B2(n_1272),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1143),
.Y(n_1407)
);

INVxp67_ASAP7_75t_SL g1408 ( 
.A(n_1143),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1285),
.A2(n_982),
.B1(n_1272),
.B2(n_1268),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1180),
.Y(n_1410)
);

INVxp67_ASAP7_75t_SL g1411 ( 
.A(n_1143),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1285),
.A2(n_1280),
.B(n_1251),
.C(n_1268),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1289),
.B(n_837),
.Y(n_1413)
);

NAND3xp33_ASAP7_75t_L g1414 ( 
.A(n_1272),
.B(n_982),
.C(n_1268),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1168),
.B(n_1183),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1168),
.B(n_1183),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1215),
.B(n_1250),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1143),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1143),
.Y(n_1419)
);

INVx5_ASAP7_75t_L g1420 ( 
.A(n_1176),
.Y(n_1420)
);

HAxp5_ASAP7_75t_L g1421 ( 
.A(n_1226),
.B(n_646),
.CON(n_1421),
.SN(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1215),
.B(n_1250),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1289),
.B(n_837),
.Y(n_1423)
);

NAND2x1p5_ASAP7_75t_L g1424 ( 
.A(n_1200),
.B(n_1215),
.Y(n_1424)
);

O2A1O1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1285),
.A2(n_1280),
.B(n_1251),
.C(n_1268),
.Y(n_1425)
);

AOI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1285),
.A2(n_982),
.B1(n_1272),
.B2(n_1268),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1151),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1143),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1168),
.B(n_1183),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1227),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1272),
.A2(n_1285),
.B(n_1268),
.C(n_982),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1227),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1143),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_SL g1434 ( 
.A(n_1204),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1285),
.B(n_837),
.Y(n_1435)
);

OAI21xp33_ASAP7_75t_L g1436 ( 
.A1(n_1285),
.A2(n_982),
.B(n_1272),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1143),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1275),
.B(n_1014),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1215),
.B(n_1250),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1285),
.B(n_837),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1147),
.A2(n_1266),
.B(n_1249),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1289),
.B(n_837),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1154),
.Y(n_1443)
);

NOR2xp67_ASAP7_75t_L g1444 ( 
.A(n_1202),
.B(n_1018),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_SL g1445 ( 
.A1(n_1251),
.A2(n_1208),
.B(n_1272),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1289),
.B(n_837),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1285),
.A2(n_982),
.B1(n_1272),
.B2(n_1268),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1143),
.Y(n_1448)
);

NAND2x1p5_ASAP7_75t_L g1449 ( 
.A(n_1200),
.B(n_1215),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1289),
.B(n_837),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1151),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1289),
.B(n_837),
.Y(n_1452)
);

BUFx2_ASAP7_75t_L g1453 ( 
.A(n_1143),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1227),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1227),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1215),
.B(n_1250),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1168),
.B(n_1183),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1143),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1154),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1143),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1184),
.A2(n_1175),
.B(n_1247),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1419),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1318),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1323),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1343),
.A2(n_1328),
.B(n_1351),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1436),
.A2(n_1399),
.B1(n_1335),
.B2(n_1309),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1297),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1399),
.A2(n_1335),
.B1(n_1414),
.B2(n_1332),
.Y(n_1468)
);

AO21x1_ASAP7_75t_L g1469 ( 
.A1(n_1412),
.A2(n_1425),
.B(n_1409),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1382),
.Y(n_1470)
);

OAI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1426),
.A2(n_1447),
.B1(n_1311),
.B2(n_1414),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1382),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1303),
.Y(n_1473)
);

AO21x2_ASAP7_75t_L g1474 ( 
.A1(n_1394),
.A2(n_1380),
.B(n_1461),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1328),
.A2(n_1347),
.B(n_1383),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1315),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1302),
.B(n_1438),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1420),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1330),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1406),
.A2(n_1301),
.B(n_1431),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1396),
.Y(n_1481)
);

INVx5_ASAP7_75t_L g1482 ( 
.A(n_1342),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1435),
.A2(n_1440),
.B1(n_1364),
.B2(n_1299),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1325),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1437),
.Y(n_1485)
);

AOI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1391),
.A2(n_1386),
.B(n_1339),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1332),
.A2(n_1324),
.B1(n_1329),
.B2(n_1307),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1443),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1461),
.A2(n_1405),
.B(n_1327),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1305),
.B(n_1403),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1448),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1427),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1337),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1300),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1459),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1312),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_SL g1497 ( 
.A1(n_1344),
.A2(n_1345),
.B(n_1348),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1316),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1324),
.A2(n_1329),
.B1(n_1333),
.B2(n_1317),
.Y(n_1499)
);

INVx6_ASAP7_75t_L g1500 ( 
.A(n_1420),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1362),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1366),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1373),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1337),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1424),
.Y(n_1505)
);

BUFx2_ASAP7_75t_SL g1506 ( 
.A(n_1451),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1424),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_SL g1508 ( 
.A1(n_1307),
.A2(n_1317),
.B1(n_1331),
.B2(n_1416),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1376),
.Y(n_1509)
);

CKINVDCx11_ASAP7_75t_R g1510 ( 
.A(n_1322),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1420),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1305),
.A2(n_1416),
.B1(n_1429),
.B2(n_1415),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1403),
.A2(n_1429),
.B1(n_1415),
.B2(n_1457),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1453),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1458),
.Y(n_1515)
);

OAI21xp5_ASAP7_75t_SL g1516 ( 
.A1(n_1341),
.A2(n_1340),
.B(n_1423),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1457),
.B(n_1358),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1357),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1413),
.B(n_1442),
.Y(n_1519)
);

AO21x1_ASAP7_75t_SL g1520 ( 
.A1(n_1379),
.A2(n_1393),
.B(n_1352),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_SL g1521 ( 
.A1(n_1368),
.A2(n_1372),
.B1(n_1375),
.B2(n_1445),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1407),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1446),
.B(n_1450),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_SL g1524 ( 
.A1(n_1375),
.A2(n_1452),
.B1(n_1411),
.B2(n_1308),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1390),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1374),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1352),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1298),
.Y(n_1528)
);

INVx1_ASAP7_75t_SL g1529 ( 
.A(n_1300),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1398),
.B(n_1401),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1360),
.A2(n_1336),
.B(n_1389),
.Y(n_1531)
);

NAND2x1p5_ASAP7_75t_L g1532 ( 
.A(n_1420),
.B(n_1350),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1449),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1389),
.A2(n_1379),
.B(n_1386),
.Y(n_1534)
);

BUFx5_ASAP7_75t_L g1535 ( 
.A(n_1381),
.Y(n_1535)
);

BUFx10_ASAP7_75t_L g1536 ( 
.A(n_1306),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1384),
.A2(n_1346),
.B(n_1363),
.Y(n_1537)
);

AO21x2_ASAP7_75t_L g1538 ( 
.A1(n_1385),
.A2(n_1370),
.B(n_1365),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_1359),
.Y(n_1539)
);

INVxp33_ASAP7_75t_L g1540 ( 
.A(n_1433),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1321),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1441),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1319),
.Y(n_1543)
);

AO21x2_ASAP7_75t_L g1544 ( 
.A1(n_1392),
.A2(n_1370),
.B(n_1349),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1319),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1434),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1410),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1342),
.B(n_1296),
.Y(n_1548)
);

BUFx4f_ASAP7_75t_SL g1549 ( 
.A(n_1367),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1342),
.A2(n_1401),
.B1(n_1398),
.B2(n_1408),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1410),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1310),
.Y(n_1552)
);

INVx4_ASAP7_75t_L g1553 ( 
.A(n_1321),
.Y(n_1553)
);

OAI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1444),
.A2(n_1367),
.B1(n_1355),
.B2(n_1400),
.Y(n_1554)
);

INVx8_ASAP7_75t_L g1555 ( 
.A(n_1354),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1314),
.A2(n_1460),
.B(n_1418),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1378),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1356),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1321),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1428),
.A2(n_1434),
.B1(n_1304),
.B2(n_1397),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1449),
.A2(n_1388),
.B(n_1369),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1296),
.B(n_1304),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1334),
.Y(n_1563)
);

BUFx12f_ASAP7_75t_L g1564 ( 
.A(n_1371),
.Y(n_1564)
);

CKINVDCx6p67_ASAP7_75t_R g1565 ( 
.A(n_1354),
.Y(n_1565)
);

BUFx2_ASAP7_75t_SL g1566 ( 
.A(n_1320),
.Y(n_1566)
);

BUFx10_ASAP7_75t_L g1567 ( 
.A(n_1397),
.Y(n_1567)
);

CKINVDCx11_ASAP7_75t_R g1568 ( 
.A(n_1334),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1313),
.Y(n_1569)
);

AO21x1_ASAP7_75t_L g1570 ( 
.A1(n_1326),
.A2(n_1404),
.B(n_1313),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1417),
.Y(n_1571)
);

CKINVDCx11_ASAP7_75t_R g1572 ( 
.A(n_1361),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1417),
.B(n_1456),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_1361),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1361),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1338),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1353),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1395),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1395),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1395),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1430),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1430),
.Y(n_1582)
);

OAI21x1_ASAP7_75t_L g1583 ( 
.A1(n_1421),
.A2(n_1326),
.B(n_1404),
.Y(n_1583)
);

AO21x2_ASAP7_75t_L g1584 ( 
.A1(n_1422),
.A2(n_1439),
.B(n_1456),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1387),
.Y(n_1585)
);

OAI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1432),
.A2(n_1454),
.B(n_1455),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1432),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1432),
.A2(n_1454),
.B(n_1455),
.Y(n_1588)
);

AO21x1_ASAP7_75t_L g1589 ( 
.A1(n_1422),
.A2(n_1439),
.B(n_1455),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1454),
.A2(n_1339),
.B(n_1377),
.Y(n_1590)
);

NAND2x1p5_ASAP7_75t_L g1591 ( 
.A(n_1420),
.B(n_1200),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1297),
.Y(n_1592)
);

INVx5_ASAP7_75t_L g1593 ( 
.A(n_1382),
.Y(n_1593)
);

NAND2x1p5_ASAP7_75t_L g1594 ( 
.A(n_1420),
.B(n_1200),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1297),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1323),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1307),
.B(n_1317),
.Y(n_1597)
);

BUFx4f_ASAP7_75t_SL g1598 ( 
.A(n_1357),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1307),
.B(n_1317),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1419),
.Y(n_1600)
);

INVx4_ASAP7_75t_SL g1601 ( 
.A(n_1382),
.Y(n_1601)
);

CKINVDCx12_ASAP7_75t_R g1602 ( 
.A(n_1342),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1297),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1297),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1325),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1307),
.B(n_1317),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1297),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1419),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1406),
.A2(n_1272),
.B1(n_982),
.B2(n_1269),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1297),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1297),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1436),
.A2(n_1285),
.B1(n_1399),
.B2(n_1335),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1297),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1307),
.B(n_1317),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1339),
.A2(n_1402),
.B(n_1377),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1297),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1300),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1297),
.Y(n_1618)
);

BUFx10_ASAP7_75t_L g1619 ( 
.A(n_1306),
.Y(n_1619)
);

INVx6_ASAP7_75t_L g1620 ( 
.A(n_1420),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1300),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1297),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1297),
.Y(n_1623)
);

OR2x6_ASAP7_75t_L g1624 ( 
.A(n_1445),
.B(n_1344),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1297),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1297),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1342),
.B(n_1365),
.Y(n_1627)
);

AO21x1_ASAP7_75t_SL g1628 ( 
.A1(n_1335),
.A2(n_1406),
.B(n_1409),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1436),
.A2(n_1285),
.B1(n_1399),
.B2(n_1335),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1323),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_SL g1631 ( 
.A1(n_1609),
.A2(n_1624),
.B1(n_1497),
.B2(n_1480),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1527),
.Y(n_1632)
);

BUFx6f_ASAP7_75t_L g1633 ( 
.A(n_1482),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1527),
.B(n_1542),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1597),
.B(n_1599),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1482),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1597),
.B(n_1599),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1606),
.B(n_1614),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1468),
.B(n_1517),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1470),
.B(n_1472),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1496),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1498),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1522),
.Y(n_1643)
);

OA21x2_ASAP7_75t_L g1644 ( 
.A1(n_1531),
.A2(n_1534),
.B(n_1489),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1534),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1470),
.B(n_1472),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1530),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1490),
.B(n_1512),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1544),
.B(n_1465),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1471),
.A2(n_1469),
.B1(n_1629),
.B2(n_1612),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1482),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1537),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1486),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1468),
.B(n_1517),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1544),
.B(n_1465),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1501),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1544),
.B(n_1465),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1612),
.A2(n_1629),
.B1(n_1483),
.B2(n_1466),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1482),
.Y(n_1659)
);

AO21x1_ASAP7_75t_SL g1660 ( 
.A1(n_1466),
.A2(n_1487),
.B(n_1499),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1615),
.A2(n_1590),
.B(n_1475),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1487),
.B(n_1520),
.Y(n_1662)
);

AOI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1624),
.A2(n_1475),
.B(n_1513),
.Y(n_1663)
);

BUFx2_ASAP7_75t_L g1664 ( 
.A(n_1538),
.Y(n_1664)
);

OAI21x1_ASAP7_75t_L g1665 ( 
.A1(n_1525),
.A2(n_1583),
.B(n_1557),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1482),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1502),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1512),
.B(n_1477),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1503),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1601),
.B(n_1627),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1628),
.A2(n_1624),
.B1(n_1521),
.B2(n_1508),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1538),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1467),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1473),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1624),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1601),
.B(n_1627),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1476),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1516),
.B(n_1523),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1535),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1535),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1535),
.Y(n_1681)
);

AO21x2_ASAP7_75t_L g1682 ( 
.A1(n_1474),
.A2(n_1543),
.B(n_1545),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1462),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1479),
.B(n_1481),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1488),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1535),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1564),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1495),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1592),
.Y(n_1689)
);

INVxp67_ASAP7_75t_L g1690 ( 
.A(n_1485),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1519),
.B(n_1550),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1478),
.Y(n_1692)
);

BUFx4f_ASAP7_75t_SL g1693 ( 
.A(n_1539),
.Y(n_1693)
);

AO21x2_ASAP7_75t_L g1694 ( 
.A1(n_1528),
.A2(n_1547),
.B(n_1551),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1595),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1535),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1535),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_1556),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1603),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1601),
.B(n_1548),
.Y(n_1700)
);

BUFx6f_ASAP7_75t_L g1701 ( 
.A(n_1478),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1491),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1604),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1607),
.B(n_1610),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1611),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1613),
.Y(n_1706)
);

OAI21x1_ASAP7_75t_L g1707 ( 
.A1(n_1561),
.A2(n_1588),
.B(n_1586),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1616),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1618),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1622),
.Y(n_1710)
);

INVx4_ASAP7_75t_L g1711 ( 
.A(n_1478),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1623),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1625),
.B(n_1626),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1600),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1509),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1526),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1589),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1550),
.B(n_1556),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1602),
.Y(n_1719)
);

OR2x6_ASAP7_75t_L g1720 ( 
.A(n_1532),
.B(n_1506),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1608),
.Y(n_1721)
);

OAI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1554),
.A2(n_1524),
.B(n_1540),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1602),
.Y(n_1723)
);

OAI21x1_ASAP7_75t_L g1724 ( 
.A1(n_1586),
.A2(n_1532),
.B(n_1533),
.Y(n_1724)
);

INVx1_ASAP7_75t_SL g1725 ( 
.A(n_1549),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1494),
.B(n_1529),
.Y(n_1726)
);

AO21x2_ASAP7_75t_L g1727 ( 
.A1(n_1558),
.A2(n_1570),
.B(n_1580),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1593),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1593),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1593),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1548),
.B(n_1584),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1617),
.B(n_1621),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1556),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1505),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1514),
.Y(n_1735)
);

OR2x6_ASAP7_75t_L g1736 ( 
.A(n_1566),
.B(n_1548),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1505),
.Y(n_1737)
);

INVxp67_ASAP7_75t_L g1738 ( 
.A(n_1552),
.Y(n_1738)
);

INVx8_ASAP7_75t_L g1739 ( 
.A(n_1555),
.Y(n_1739)
);

OAI21x1_ASAP7_75t_L g1740 ( 
.A1(n_1507),
.A2(n_1533),
.B(n_1504),
.Y(n_1740)
);

OA21x2_ASAP7_75t_L g1741 ( 
.A1(n_1576),
.A2(n_1577),
.B(n_1560),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1569),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1493),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1515),
.Y(n_1744)
);

OA21x2_ASAP7_75t_L g1745 ( 
.A1(n_1560),
.A2(n_1563),
.B(n_1575),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1578),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1584),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1581),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1584),
.Y(n_1749)
);

OR2x6_ASAP7_75t_L g1750 ( 
.A(n_1500),
.B(n_1620),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1500),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1463),
.B(n_1540),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1656),
.Y(n_1753)
);

INVxp67_ASAP7_75t_SL g1754 ( 
.A(n_1733),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1648),
.B(n_1515),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1733),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1731),
.Y(n_1757)
);

AOI222xp33_ASAP7_75t_L g1758 ( 
.A1(n_1650),
.A2(n_1678),
.B1(n_1671),
.B2(n_1722),
.C1(n_1668),
.C2(n_1639),
.Y(n_1758)
);

BUFx3_ASAP7_75t_L g1759 ( 
.A(n_1720),
.Y(n_1759)
);

AO21x2_ASAP7_75t_L g1760 ( 
.A1(n_1653),
.A2(n_1582),
.B(n_1587),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1652),
.B(n_1645),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1698),
.Y(n_1762)
);

NAND2x1_ASAP7_75t_L g1763 ( 
.A(n_1675),
.B(n_1620),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1707),
.Y(n_1764)
);

INVxp67_ASAP7_75t_L g1765 ( 
.A(n_1718),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1731),
.B(n_1571),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1639),
.B(n_1464),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1731),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1698),
.Y(n_1769)
);

INVx1_ASAP7_75t_SL g1770 ( 
.A(n_1643),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1635),
.B(n_1630),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1635),
.B(n_1596),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1631),
.A2(n_1539),
.B1(n_1571),
.B2(n_1510),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1637),
.B(n_1579),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1637),
.B(n_1638),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1638),
.B(n_1562),
.Y(n_1776)
);

INVxp67_ASAP7_75t_L g1777 ( 
.A(n_1718),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1634),
.Y(n_1778)
);

AO21x2_ASAP7_75t_L g1779 ( 
.A1(n_1653),
.A2(n_1573),
.B(n_1500),
.Y(n_1779)
);

BUFx2_ASAP7_75t_SL g1780 ( 
.A(n_1687),
.Y(n_1780)
);

INVxp67_ASAP7_75t_SL g1781 ( 
.A(n_1649),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1654),
.B(n_1559),
.Y(n_1782)
);

AND2x4_ASAP7_75t_SL g1783 ( 
.A(n_1633),
.B(n_1567),
.Y(n_1783)
);

INVx4_ASAP7_75t_L g1784 ( 
.A(n_1720),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1694),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1747),
.B(n_1559),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1654),
.B(n_1565),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1749),
.B(n_1559),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1649),
.B(n_1492),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1655),
.B(n_1492),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1655),
.B(n_1559),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1694),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1657),
.B(n_1541),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1657),
.B(n_1565),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1662),
.B(n_1541),
.Y(n_1795)
);

BUFx3_ASAP7_75t_L g1796 ( 
.A(n_1720),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1682),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1691),
.B(n_1574),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1693),
.B(n_1725),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1632),
.B(n_1541),
.Y(n_1800)
);

OAI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1658),
.A2(n_1585),
.B1(n_1546),
.B2(n_1478),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1665),
.B(n_1553),
.Y(n_1802)
);

BUFx2_ASAP7_75t_L g1803 ( 
.A(n_1665),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1664),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1691),
.B(n_1574),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1663),
.B(n_1541),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1641),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1664),
.Y(n_1808)
);

HB1xp67_ASAP7_75t_L g1809 ( 
.A(n_1672),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1642),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1660),
.A2(n_1510),
.B1(n_1564),
.B2(n_1518),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1667),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1669),
.Y(n_1813)
);

BUFx2_ASAP7_75t_L g1814 ( 
.A(n_1675),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1753),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1755),
.B(n_1647),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1755),
.B(n_1683),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_R g1818 ( 
.A(n_1811),
.B(n_1484),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1758),
.B(n_1640),
.Y(n_1819)
);

NAND3xp33_ASAP7_75t_L g1820 ( 
.A(n_1758),
.B(n_1717),
.C(n_1741),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1791),
.B(n_1679),
.Y(n_1821)
);

NOR3xp33_ASAP7_75t_L g1822 ( 
.A(n_1801),
.B(n_1719),
.C(n_1723),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1770),
.B(n_1702),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1770),
.B(n_1714),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1767),
.B(n_1721),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1791),
.B(n_1680),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1801),
.B(n_1640),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1767),
.B(n_1716),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1775),
.B(n_1716),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1753),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1773),
.A2(n_1660),
.B1(n_1719),
.B2(n_1723),
.Y(n_1831)
);

OAI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1763),
.A2(n_1752),
.B1(n_1690),
.B2(n_1738),
.C(n_1735),
.Y(n_1832)
);

OA21x2_ASAP7_75t_L g1833 ( 
.A1(n_1785),
.A2(n_1661),
.B(n_1707),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1780),
.A2(n_1720),
.B1(n_1736),
.B2(n_1750),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1791),
.B(n_1793),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1787),
.A2(n_1717),
.B1(n_1640),
.B2(n_1646),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1793),
.B(n_1680),
.Y(n_1837)
);

NAND3xp33_ASAP7_75t_L g1838 ( 
.A(n_1789),
.B(n_1741),
.C(n_1742),
.Y(n_1838)
);

OAI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1763),
.A2(n_1736),
.B1(n_1750),
.B2(n_1666),
.Y(n_1839)
);

OAI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1789),
.A2(n_1744),
.B1(n_1732),
.B2(n_1726),
.C(n_1736),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1775),
.B(n_1688),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1776),
.B(n_1782),
.Y(n_1842)
);

NAND3xp33_ASAP7_75t_L g1843 ( 
.A(n_1790),
.B(n_1741),
.C(n_1745),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1757),
.B(n_1681),
.Y(n_1844)
);

INVx4_ASAP7_75t_L g1845 ( 
.A(n_1784),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1768),
.B(n_1686),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1776),
.B(n_1688),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1768),
.B(n_1696),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1782),
.B(n_1689),
.Y(n_1849)
);

INVxp67_ASAP7_75t_L g1850 ( 
.A(n_1790),
.Y(n_1850)
);

AOI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1779),
.A2(n_1750),
.B(n_1644),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1765),
.B(n_1696),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1771),
.B(n_1772),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1765),
.B(n_1697),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1771),
.B(n_1689),
.Y(n_1855)
);

OAI221xp5_ASAP7_75t_L g1856 ( 
.A1(n_1799),
.A2(n_1736),
.B1(n_1687),
.B2(n_1518),
.C(n_1546),
.Y(n_1856)
);

OA21x2_ASAP7_75t_L g1857 ( 
.A1(n_1785),
.A2(n_1661),
.B(n_1724),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1780),
.A2(n_1750),
.B1(n_1585),
.B2(n_1700),
.Y(n_1858)
);

OA211x2_ASAP7_75t_L g1859 ( 
.A1(n_1777),
.A2(n_1727),
.B(n_1745),
.C(n_1724),
.Y(n_1859)
);

OAI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1798),
.A2(n_1700),
.B1(n_1670),
.B2(n_1676),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1772),
.B(n_1712),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_L g1862 ( 
.A(n_1795),
.B(n_1536),
.Y(n_1862)
);

OAI221xp5_ASAP7_75t_SL g1863 ( 
.A1(n_1798),
.A2(n_1685),
.B1(n_1673),
.B2(n_1674),
.C(n_1677),
.Y(n_1863)
);

OAI21xp5_ASAP7_75t_SL g1864 ( 
.A1(n_1783),
.A2(n_1700),
.B(n_1676),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1786),
.B(n_1788),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1805),
.B(n_1712),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1805),
.B(n_1715),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1807),
.B(n_1715),
.Y(n_1868)
);

OAI221xp5_ASAP7_75t_SL g1869 ( 
.A1(n_1794),
.A2(n_1806),
.B1(n_1814),
.B2(n_1781),
.C(n_1796),
.Y(n_1869)
);

OA21x2_ASAP7_75t_L g1870 ( 
.A1(n_1792),
.A2(n_1740),
.B(n_1730),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1807),
.B(n_1695),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_SL g1872 ( 
.A1(n_1783),
.A2(n_1670),
.B(n_1730),
.Y(n_1872)
);

OAI21xp33_ASAP7_75t_L g1873 ( 
.A1(n_1781),
.A2(n_1709),
.B(n_1710),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1774),
.B(n_1536),
.Y(n_1874)
);

OAI221xp5_ASAP7_75t_L g1875 ( 
.A1(n_1784),
.A2(n_1751),
.B1(n_1705),
.B2(n_1699),
.C(n_1703),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1810),
.B(n_1706),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1810),
.B(n_1708),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1784),
.A2(n_1751),
.B1(n_1666),
.B2(n_1633),
.Y(n_1878)
);

NAND4xp25_ASAP7_75t_L g1879 ( 
.A(n_1800),
.B(n_1746),
.C(n_1748),
.D(n_1713),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1812),
.B(n_1684),
.Y(n_1880)
);

AOI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1766),
.A2(n_1636),
.B1(n_1659),
.B2(n_1651),
.Y(n_1881)
);

OAI21xp5_ASAP7_75t_SL g1882 ( 
.A1(n_1783),
.A2(n_1728),
.B(n_1729),
.Y(n_1882)
);

NAND3xp33_ASAP7_75t_L g1883 ( 
.A(n_1797),
.B(n_1745),
.C(n_1734),
.Y(n_1883)
);

OAI221xp5_ASAP7_75t_L g1884 ( 
.A1(n_1784),
.A2(n_1729),
.B1(n_1728),
.B2(n_1484),
.C(n_1605),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1813),
.B(n_1713),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1766),
.A2(n_1743),
.B1(n_1739),
.B2(n_1737),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1815),
.Y(n_1887)
);

BUFx6f_ASAP7_75t_L g1888 ( 
.A(n_1845),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1849),
.B(n_1762),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1815),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1835),
.B(n_1806),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1845),
.B(n_1806),
.Y(n_1892)
);

NAND2x1p5_ASAP7_75t_L g1893 ( 
.A(n_1845),
.B(n_1759),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1850),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1835),
.B(n_1865),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1830),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1865),
.B(n_1802),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1830),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1828),
.B(n_1769),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1816),
.B(n_1769),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1847),
.B(n_1756),
.Y(n_1901)
);

INVxp33_ASAP7_75t_L g1902 ( 
.A(n_1862),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1871),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1876),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1825),
.B(n_1804),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1842),
.B(n_1804),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1870),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1852),
.B(n_1756),
.Y(n_1908)
);

HB1xp67_ASAP7_75t_L g1909 ( 
.A(n_1870),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1870),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1877),
.Y(n_1911)
);

OAI21xp33_ASAP7_75t_L g1912 ( 
.A1(n_1820),
.A2(n_1704),
.B(n_1759),
.Y(n_1912)
);

INVxp67_ASAP7_75t_L g1913 ( 
.A(n_1819),
.Y(n_1913)
);

INVx2_ASAP7_75t_SL g1914 ( 
.A(n_1854),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1833),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1854),
.B(n_1754),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1833),
.Y(n_1917)
);

INVx3_ASAP7_75t_L g1918 ( 
.A(n_1857),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1866),
.B(n_1808),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1833),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1867),
.B(n_1754),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1841),
.B(n_1809),
.Y(n_1922)
);

AND2x2_ASAP7_75t_SL g1923 ( 
.A(n_1822),
.B(n_1766),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1821),
.B(n_1786),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1817),
.B(n_1760),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1821),
.B(n_1786),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1856),
.B(n_1536),
.Y(n_1927)
);

INVx2_ASAP7_75t_SL g1928 ( 
.A(n_1844),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1868),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1826),
.B(n_1788),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1826),
.B(n_1788),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1857),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1837),
.B(n_1761),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1880),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1885),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1873),
.B(n_1778),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1857),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1829),
.B(n_1778),
.Y(n_1938)
);

OR2x2_ASAP7_75t_L g1939 ( 
.A(n_1925),
.B(n_1823),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1925),
.B(n_1824),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1908),
.B(n_1855),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1890),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1890),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1887),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1923),
.B(n_1913),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1897),
.B(n_1846),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1887),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1890),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1896),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1908),
.B(n_1869),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1905),
.B(n_1861),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1913),
.B(n_1853),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1897),
.B(n_1848),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1896),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1897),
.B(n_1923),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1896),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1897),
.B(n_1848),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1903),
.B(n_1879),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1905),
.B(n_1838),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1898),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1898),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1923),
.B(n_1881),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1891),
.B(n_1766),
.Y(n_1963)
);

OR2x2_ASAP7_75t_L g1964 ( 
.A(n_1916),
.B(n_1843),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1898),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1907),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1903),
.B(n_1774),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1907),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1929),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1916),
.B(n_1883),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1904),
.B(n_1874),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1929),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1904),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1891),
.B(n_1759),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1911),
.B(n_1840),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1895),
.B(n_1796),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1895),
.B(n_1796),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1911),
.B(n_1819),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1919),
.B(n_1760),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1900),
.B(n_1882),
.Y(n_1980)
);

NAND2x1_ASAP7_75t_L g1981 ( 
.A(n_1892),
.B(n_1803),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1894),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1907),
.Y(n_1983)
);

NOR2xp33_ASAP7_75t_R g1984 ( 
.A(n_1927),
.B(n_1605),
.Y(n_1984)
);

NOR2x1_ASAP7_75t_L g1985 ( 
.A(n_1900),
.B(n_1832),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1919),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1906),
.B(n_1760),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1906),
.B(n_1922),
.Y(n_1988)
);

O2A1O1Ixp5_ASAP7_75t_L g1989 ( 
.A1(n_1892),
.A2(n_1827),
.B(n_1839),
.C(n_1834),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1944),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1966),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1947),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1973),
.Y(n_1993)
);

INVx1_ASAP7_75t_SL g1994 ( 
.A(n_1984),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1955),
.B(n_1892),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1966),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1978),
.B(n_1938),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1985),
.B(n_1934),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1969),
.Y(n_1999)
);

NAND2x1p5_ASAP7_75t_L g2000 ( 
.A(n_1981),
.B(n_1888),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1975),
.B(n_1934),
.Y(n_2001)
);

AND2x2_ASAP7_75t_SL g2002 ( 
.A(n_1962),
.B(n_1831),
.Y(n_2002)
);

AO22x1_ASAP7_75t_L g2003 ( 
.A1(n_1962),
.A2(n_1902),
.B1(n_1888),
.B2(n_1892),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1972),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1958),
.B(n_1935),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1955),
.B(n_1924),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1982),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_1976),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1986),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1942),
.Y(n_2010)
);

OAI31xp33_ASAP7_75t_L g2011 ( 
.A1(n_1945),
.A2(n_1912),
.A3(n_1884),
.B(n_1893),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1942),
.Y(n_2012)
);

NOR2x1_ASAP7_75t_L g2013 ( 
.A(n_1980),
.B(n_1959),
.Y(n_2013)
);

AND2x4_ASAP7_75t_L g2014 ( 
.A(n_1946),
.B(n_1953),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1943),
.Y(n_2015)
);

OR2x2_ASAP7_75t_L g2016 ( 
.A(n_1988),
.B(n_1938),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1946),
.B(n_1924),
.Y(n_2017)
);

INVx3_ASAP7_75t_SL g2018 ( 
.A(n_1959),
.Y(n_2018)
);

INVx1_ASAP7_75t_SL g2019 ( 
.A(n_1971),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1952),
.B(n_1935),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1943),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1964),
.B(n_1901),
.Y(n_2022)
);

AND2x4_ASAP7_75t_L g2023 ( 
.A(n_1953),
.B(n_1957),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1960),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1950),
.B(n_1912),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1950),
.B(n_1926),
.Y(n_2026)
);

AOI31xp33_ASAP7_75t_L g2027 ( 
.A1(n_1964),
.A2(n_1893),
.A3(n_1858),
.B(n_1827),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1968),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1960),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1957),
.B(n_1926),
.Y(n_2030)
);

OR2x2_ASAP7_75t_L g2031 ( 
.A(n_1988),
.B(n_1970),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1963),
.B(n_1930),
.Y(n_2032)
);

HB1xp67_ASAP7_75t_L g2033 ( 
.A(n_1948),
.Y(n_2033)
);

NAND2xp33_ASAP7_75t_L g2034 ( 
.A(n_1970),
.B(n_1818),
.Y(n_2034)
);

AO32x1_ASAP7_75t_L g2035 ( 
.A1(n_1968),
.A2(n_1878),
.A3(n_1764),
.B1(n_1983),
.B2(n_1711),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1941),
.B(n_1930),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1941),
.B(n_1931),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1961),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1951),
.B(n_1931),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1951),
.B(n_1889),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_2018),
.B(n_1963),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_2031),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2019),
.B(n_1939),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1991),
.Y(n_2044)
);

INVx3_ASAP7_75t_L g2045 ( 
.A(n_2000),
.Y(n_2045)
);

NOR2xp33_ASAP7_75t_L g2046 ( 
.A(n_1994),
.B(n_1619),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2018),
.B(n_1976),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1992),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_R g2049 ( 
.A(n_2034),
.B(n_1598),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1992),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_2006),
.B(n_1977),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_2031),
.B(n_1939),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1990),
.Y(n_2053)
);

INVx1_ASAP7_75t_SL g2054 ( 
.A(n_2034),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2006),
.B(n_1977),
.Y(n_2055)
);

INVxp67_ASAP7_75t_L g2056 ( 
.A(n_2013),
.Y(n_2056)
);

OR2x2_ASAP7_75t_L g2057 ( 
.A(n_2022),
.B(n_1940),
.Y(n_2057)
);

AND2x2_ASAP7_75t_SL g2058 ( 
.A(n_2002),
.B(n_1888),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_2002),
.B(n_1619),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2033),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2033),
.Y(n_2061)
);

INVxp33_ASAP7_75t_L g2062 ( 
.A(n_2026),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1991),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1995),
.B(n_1989),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1993),
.Y(n_2065)
);

OAI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_2011),
.A2(n_1940),
.B(n_1981),
.Y(n_2066)
);

NOR2x1_ASAP7_75t_L g2067 ( 
.A(n_1998),
.B(n_1983),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2001),
.B(n_1967),
.Y(n_2068)
);

INVx3_ASAP7_75t_L g2069 ( 
.A(n_2000),
.Y(n_2069)
);

INVx1_ASAP7_75t_SL g2070 ( 
.A(n_2008),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_2025),
.B(n_2005),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2007),
.B(n_1974),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1999),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1996),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_1995),
.B(n_1974),
.Y(n_2075)
);

INVx1_ASAP7_75t_SL g2076 ( 
.A(n_2003),
.Y(n_2076)
);

OR2x2_ASAP7_75t_L g2077 ( 
.A(n_2022),
.B(n_1987),
.Y(n_2077)
);

INVx1_ASAP7_75t_SL g2078 ( 
.A(n_1997),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_2014),
.B(n_1933),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2004),
.Y(n_2080)
);

AOI22xp33_ASAP7_75t_SL g2081 ( 
.A1(n_2027),
.A2(n_1818),
.B1(n_1888),
.B2(n_1860),
.Y(n_2081)
);

AOI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_2058),
.A2(n_2035),
.B(n_2009),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2042),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2056),
.B(n_2071),
.Y(n_2084)
);

XOR2x2_ASAP7_75t_L g2085 ( 
.A(n_2058),
.B(n_2059),
.Y(n_2085)
);

AOI332xp33_ASAP7_75t_L g2086 ( 
.A1(n_2048),
.A2(n_2015),
.A3(n_2024),
.B1(n_2038),
.B2(n_2010),
.B3(n_2012),
.C1(n_2021),
.C2(n_2029),
.Y(n_2086)
);

OAI21xp33_ASAP7_75t_SL g2087 ( 
.A1(n_2058),
.A2(n_2030),
.B(n_2017),
.Y(n_2087)
);

OAI21xp33_ASAP7_75t_L g2088 ( 
.A1(n_2062),
.A2(n_2064),
.B(n_2081),
.Y(n_2088)
);

OAI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_2076),
.A2(n_1859),
.B1(n_1893),
.B2(n_2014),
.Y(n_2089)
);

OAI221xp5_ASAP7_75t_L g2090 ( 
.A1(n_2066),
.A2(n_2020),
.B1(n_2040),
.B2(n_2016),
.C(n_2036),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2048),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_2047),
.Y(n_2092)
);

OAI32xp33_ASAP7_75t_L g2093 ( 
.A1(n_2054),
.A2(n_1909),
.A3(n_2037),
.B1(n_1987),
.B2(n_1979),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2070),
.B(n_2039),
.Y(n_2094)
);

AOI31xp33_ASAP7_75t_L g2095 ( 
.A1(n_2070),
.A2(n_2014),
.A3(n_2023),
.B(n_2030),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2047),
.B(n_2023),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_2078),
.B(n_2050),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2050),
.Y(n_2098)
);

AOI211xp5_ASAP7_75t_L g2099 ( 
.A1(n_2049),
.A2(n_1888),
.B(n_1996),
.C(n_2028),
.Y(n_2099)
);

AOI22xp33_ASAP7_75t_L g2100 ( 
.A1(n_2064),
.A2(n_2023),
.B1(n_1888),
.B2(n_1836),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2053),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2041),
.B(n_2017),
.Y(n_2102)
);

AOI211xp5_ASAP7_75t_L g2103 ( 
.A1(n_2041),
.A2(n_2028),
.B(n_1875),
.C(n_1872),
.Y(n_2103)
);

NAND2x1p5_ASAP7_75t_L g2104 ( 
.A(n_2045),
.B(n_1511),
.Y(n_2104)
);

INVx2_ASAP7_75t_SL g2105 ( 
.A(n_2045),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2053),
.Y(n_2106)
);

AOI222xp33_ASAP7_75t_L g2107 ( 
.A1(n_2043),
.A2(n_1909),
.B1(n_1936),
.B2(n_2032),
.C1(n_1921),
.C2(n_1910),
.Y(n_2107)
);

AOI21xp5_ASAP7_75t_L g2108 ( 
.A1(n_2046),
.A2(n_2035),
.B(n_1936),
.Y(n_2108)
);

AOI22xp5_ASAP7_75t_L g2109 ( 
.A1(n_2072),
.A2(n_1864),
.B1(n_2032),
.B2(n_1886),
.Y(n_2109)
);

A2O1A1Ixp33_ASAP7_75t_L g2110 ( 
.A1(n_2067),
.A2(n_1979),
.B(n_1863),
.C(n_1851),
.Y(n_2110)
);

CKINVDCx5p33_ASAP7_75t_R g2111 ( 
.A(n_2084),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2083),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2092),
.B(n_2051),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2096),
.B(n_2075),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2097),
.Y(n_2115)
);

NOR2x1p5_ASAP7_75t_L g2116 ( 
.A(n_2084),
.B(n_2045),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2097),
.Y(n_2117)
);

OR2x2_ASAP7_75t_L g2118 ( 
.A(n_2094),
.B(n_2052),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2088),
.B(n_2102),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2101),
.Y(n_2120)
);

OR2x2_ASAP7_75t_L g2121 ( 
.A(n_2094),
.B(n_2052),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2095),
.B(n_2051),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2091),
.B(n_2055),
.Y(n_2123)
);

NOR3xp33_ASAP7_75t_L g2124 ( 
.A(n_2099),
.B(n_2087),
.C(n_2098),
.Y(n_2124)
);

NOR2xp33_ASAP7_75t_L g2125 ( 
.A(n_2090),
.B(n_2068),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2105),
.B(n_2055),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2100),
.B(n_2075),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2106),
.Y(n_2128)
);

AOI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_2085),
.A2(n_2045),
.B1(n_2069),
.B2(n_2067),
.Y(n_2129)
);

NOR2x1p5_ASAP7_75t_L g2130 ( 
.A(n_2086),
.B(n_2069),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2108),
.B(n_2079),
.Y(n_2131)
);

HB1xp67_ASAP7_75t_L g2132 ( 
.A(n_2104),
.Y(n_2132)
);

INVx1_ASAP7_75t_SL g2133 ( 
.A(n_2104),
.Y(n_2133)
);

INVx1_ASAP7_75t_SL g2134 ( 
.A(n_2089),
.Y(n_2134)
);

NOR3xp33_ASAP7_75t_L g2135 ( 
.A(n_2119),
.B(n_2089),
.C(n_2110),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_L g2136 ( 
.A(n_2111),
.B(n_2109),
.Y(n_2136)
);

OAI21xp33_ASAP7_75t_L g2137 ( 
.A1(n_2122),
.A2(n_2107),
.B(n_2103),
.Y(n_2137)
);

AOI21xp5_ASAP7_75t_L g2138 ( 
.A1(n_2125),
.A2(n_2082),
.B(n_2093),
.Y(n_2138)
);

NAND3xp33_ASAP7_75t_L g2139 ( 
.A(n_2124),
.B(n_2111),
.C(n_2129),
.Y(n_2139)
);

AOI221x1_ASAP7_75t_L g2140 ( 
.A1(n_2115),
.A2(n_2061),
.B1(n_2060),
.B2(n_2069),
.C(n_2073),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2123),
.Y(n_2141)
);

NAND3xp33_ASAP7_75t_L g2142 ( 
.A(n_2117),
.B(n_2061),
.C(n_2060),
.Y(n_2142)
);

AOI211xp5_ASAP7_75t_L g2143 ( 
.A1(n_2125),
.A2(n_2134),
.B(n_2131),
.C(n_2127),
.Y(n_2143)
);

NOR2xp33_ASAP7_75t_R g2144 ( 
.A(n_2112),
.B(n_1619),
.Y(n_2144)
);

NAND4xp25_ASAP7_75t_SL g2145 ( 
.A(n_2127),
.B(n_2057),
.C(n_2079),
.D(n_2077),
.Y(n_2145)
);

NOR3xp33_ASAP7_75t_SL g2146 ( 
.A(n_2113),
.B(n_2073),
.C(n_2065),
.Y(n_2146)
);

AOI221xp5_ASAP7_75t_L g2147 ( 
.A1(n_2126),
.A2(n_2080),
.B1(n_2065),
.B2(n_2069),
.C(n_2074),
.Y(n_2147)
);

AOI21xp5_ASAP7_75t_L g2148 ( 
.A1(n_2121),
.A2(n_2080),
.B(n_2057),
.Y(n_2148)
);

OAI21xp5_ASAP7_75t_L g2149 ( 
.A1(n_2121),
.A2(n_2063),
.B(n_2044),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2142),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2149),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2143),
.B(n_2130),
.Y(n_2152)
);

NAND4xp25_ASAP7_75t_L g2153 ( 
.A(n_2139),
.B(n_2118),
.C(n_2128),
.D(n_2120),
.Y(n_2153)
);

NOR3xp33_ASAP7_75t_L g2154 ( 
.A(n_2136),
.B(n_2114),
.C(n_2133),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2140),
.Y(n_2155)
);

NOR4xp25_ASAP7_75t_L g2156 ( 
.A(n_2137),
.B(n_2114),
.C(n_2063),
.D(n_2044),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2148),
.B(n_2138),
.Y(n_2157)
);

AOI211x1_ASAP7_75t_L g2158 ( 
.A1(n_2145),
.A2(n_2116),
.B(n_2132),
.C(n_1961),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2141),
.Y(n_2159)
);

OAI21xp33_ASAP7_75t_L g2160 ( 
.A1(n_2135),
.A2(n_2063),
.B(n_2044),
.Y(n_2160)
);

NAND3xp33_ASAP7_75t_SL g2161 ( 
.A(n_2157),
.B(n_2152),
.C(n_2154),
.Y(n_2161)
);

NAND4xp25_ASAP7_75t_L g2162 ( 
.A(n_2153),
.B(n_2147),
.C(n_2144),
.D(n_2146),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2156),
.B(n_2074),
.Y(n_2163)
);

AOI211xp5_ASAP7_75t_L g2164 ( 
.A1(n_2150),
.A2(n_2074),
.B(n_2077),
.C(n_1910),
.Y(n_2164)
);

NAND2x1_ASAP7_75t_L g2165 ( 
.A(n_2158),
.B(n_1948),
.Y(n_2165)
);

BUFx3_ASAP7_75t_L g2166 ( 
.A(n_2159),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_2165),
.Y(n_2167)
);

AOI22xp5_ASAP7_75t_L g2168 ( 
.A1(n_2161),
.A2(n_2155),
.B1(n_2162),
.B2(n_2151),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2163),
.Y(n_2169)
);

AOI22xp5_ASAP7_75t_L g2170 ( 
.A1(n_2166),
.A2(n_2160),
.B1(n_1568),
.B2(n_1572),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2164),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2166),
.B(n_1949),
.Y(n_2172)
);

NOR2x2_ASAP7_75t_L g2173 ( 
.A(n_2161),
.B(n_1568),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2167),
.Y(n_2174)
);

AOI21xp33_ASAP7_75t_L g2175 ( 
.A1(n_2169),
.A2(n_2168),
.B(n_2170),
.Y(n_2175)
);

OAI211xp5_ASAP7_75t_SL g2176 ( 
.A1(n_2171),
.A2(n_2172),
.B(n_2173),
.C(n_1572),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_L g2177 ( 
.A(n_2168),
.B(n_1956),
.Y(n_2177)
);

INVx3_ASAP7_75t_L g2178 ( 
.A(n_2167),
.Y(n_2178)
);

NAND4xp75_ASAP7_75t_L g2179 ( 
.A(n_2168),
.B(n_2035),
.C(n_1954),
.D(n_1910),
.Y(n_2179)
);

AOI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_2176),
.A2(n_1918),
.B1(n_1965),
.B2(n_1956),
.Y(n_2180)
);

NOR3xp33_ASAP7_75t_SL g2181 ( 
.A(n_2175),
.B(n_1921),
.C(n_1889),
.Y(n_2181)
);

BUFx2_ASAP7_75t_L g2182 ( 
.A(n_2178),
.Y(n_2182)
);

XNOR2xp5_ASAP7_75t_SL g2183 ( 
.A(n_2182),
.B(n_2174),
.Y(n_2183)
);

OAI22xp5_ASAP7_75t_SL g2184 ( 
.A1(n_2183),
.A2(n_2177),
.B1(n_2180),
.B2(n_2181),
.Y(n_2184)
);

AOI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_2184),
.A2(n_2179),
.B1(n_1965),
.B2(n_1918),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2184),
.Y(n_2186)
);

OAI22xp5_ASAP7_75t_L g2187 ( 
.A1(n_2185),
.A2(n_1918),
.B1(n_1932),
.B2(n_1937),
.Y(n_2187)
);

AOI31xp33_ASAP7_75t_L g2188 ( 
.A1(n_2186),
.A2(n_1594),
.A3(n_1591),
.B(n_1651),
.Y(n_2188)
);

AOI22xp33_ASAP7_75t_L g2189 ( 
.A1(n_2187),
.A2(n_1918),
.B1(n_1932),
.B2(n_1937),
.Y(n_2189)
);

AOI22xp33_ASAP7_75t_L g2190 ( 
.A1(n_2188),
.A2(n_1932),
.B1(n_1937),
.B2(n_1915),
.Y(n_2190)
);

OAI21xp5_ASAP7_75t_L g2191 ( 
.A1(n_2189),
.A2(n_1899),
.B(n_1901),
.Y(n_2191)
);

AOI322xp5_ASAP7_75t_L g2192 ( 
.A1(n_2191),
.A2(n_2190),
.A3(n_1920),
.B1(n_1917),
.B2(n_1915),
.C1(n_1928),
.C2(n_1914),
.Y(n_2192)
);

AOI221xp5_ASAP7_75t_L g2193 ( 
.A1(n_2192),
.A2(n_1511),
.B1(n_1920),
.B2(n_1915),
.C(n_1917),
.Y(n_2193)
);

AOI211xp5_ASAP7_75t_L g2194 ( 
.A1(n_2193),
.A2(n_1511),
.B(n_1692),
.C(n_1701),
.Y(n_2194)
);


endmodule