module fake_netlist_6_4486_n_1852 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1852);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1852;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g175 ( 
.A(n_77),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_35),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_38),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_44),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_7),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_108),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_85),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_29),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_81),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_68),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_79),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_152),
.Y(n_186)
);

BUFx2_ASAP7_75t_SL g187 ( 
.A(n_173),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_35),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_133),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_43),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_115),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_74),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_48),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_86),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_70),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_37),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_23),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_32),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_136),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_146),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_142),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_127),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_143),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_52),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_83),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_18),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_116),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_75),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_56),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_125),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_3),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_94),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_43),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_90),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_129),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_154),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_46),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_8),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_88),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_145),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_165),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_119),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_84),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_113),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_42),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_150),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_14),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_172),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_103),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_7),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_47),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_56),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_156),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_128),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_149),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_139),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_109),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_121),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_50),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_38),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_137),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_37),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_162),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_41),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_163),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_122),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_170),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_31),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_91),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_147),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_76),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_36),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_134),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_63),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g259 ( 
.A(n_57),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_1),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_82),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_87),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_53),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_59),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_120),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_135),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_47),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_97),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_61),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_15),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_27),
.Y(n_271)
);

BUFx8_ASAP7_75t_SL g272 ( 
.A(n_63),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_144),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_42),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_99),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_30),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_27),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_48),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_52),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_101),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_19),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_12),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_21),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_167),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_57),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_11),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_18),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_67),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_45),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_118),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_26),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_50),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_36),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_39),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_104),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_106),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_98),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_2),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_11),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_117),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_26),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_16),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_161),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_5),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_140),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_66),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_51),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_16),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_8),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_89),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_164),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_72),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_126),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_153),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_54),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_49),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_138),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_23),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_62),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_9),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_132),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_0),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_54),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_114),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_102),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_3),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_168),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_49),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_15),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_69),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_40),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_55),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_21),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_59),
.Y(n_334)
);

BUFx10_ASAP7_75t_L g335 ( 
.A(n_5),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_95),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_112),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_158),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_25),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_105),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_39),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_0),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_141),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_171),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_148),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_13),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_80),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_32),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_205),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_259),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_284),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_259),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_299),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_259),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_259),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_259),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_259),
.B(n_1),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_259),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_259),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_237),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_196),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_196),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_272),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_196),
.Y(n_364)
);

INVxp33_ASAP7_75t_SL g365 ( 
.A(n_236),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_225),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_196),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_230),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_296),
.Y(n_369)
);

INVxp33_ASAP7_75t_SL g370 ( 
.A(n_182),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g371 ( 
.A(n_256),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_310),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_232),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_196),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_326),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_300),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_194),
.B(n_2),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_233),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_337),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_326),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_326),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_326),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_177),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_239),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_309),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_177),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_240),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_269),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_269),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_178),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_178),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_279),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_254),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_176),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_241),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_335),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_245),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_247),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_250),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_279),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_301),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_335),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_253),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_181),
.B(n_4),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_301),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_179),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_255),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_182),
.Y(n_409)
);

INVxp33_ASAP7_75t_SL g410 ( 
.A(n_193),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_321),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_266),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_188),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_190),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_335),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_305),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_200),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_213),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_220),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_180),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_228),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_180),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_231),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_194),
.B(n_4),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_305),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_234),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_244),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_258),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_243),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_271),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_248),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_252),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_260),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_235),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_274),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_183),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_R g437 ( 
.A(n_394),
.B(n_426),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_366),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_368),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_361),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_361),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_215),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_R g443 ( 
.A(n_429),
.B(n_183),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_362),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_362),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_373),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_364),
.B(n_184),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_378),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_385),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_416),
.B(n_215),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_349),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_353),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_374),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_380),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_364),
.B(n_184),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_380),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_431),
.B(n_432),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_388),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_396),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_367),
.B(n_189),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_409),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_367),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_350),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_400),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_412),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_398),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_351),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_375),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_399),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_375),
.Y(n_471)
);

NAND2xp33_ASAP7_75t_R g472 ( 
.A(n_433),
.B(n_370),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_381),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_381),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_386),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_404),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_350),
.Y(n_477)
);

AND3x2_ASAP7_75t_L g478 ( 
.A(n_405),
.B(n_285),
.C(n_199),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_411),
.B(n_185),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_416),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_408),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_416),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_434),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_382),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_R g485 ( 
.A(n_410),
.B(n_189),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_420),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_382),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_383),
.B(n_191),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_422),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_383),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_369),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_352),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_352),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_354),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_354),
.B(n_175),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_436),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_355),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_355),
.B(n_191),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_356),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_356),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_358),
.B(n_175),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_358),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_359),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_363),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_391),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_376),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_359),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_360),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_395),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_384),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_357),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_397),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_379),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_384),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_482),
.B(n_395),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_511),
.B(n_377),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_372),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_508),
.B(n_372),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_483),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_492),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_445),
.Y(n_521)
);

INVxp33_ASAP7_75t_L g522 ( 
.A(n_475),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_492),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_482),
.B(n_407),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_494),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_500),
.Y(n_526)
);

INVx4_ASAP7_75t_L g527 ( 
.A(n_494),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_500),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_511),
.B(n_199),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_511),
.B(n_424),
.Y(n_530)
);

AOI22x1_ASAP7_75t_L g531 ( 
.A1(n_451),
.A2(n_207),
.B1(n_343),
.B2(n_345),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_445),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_507),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_494),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_458),
.B(n_365),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_507),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_451),
.B(n_435),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_445),
.Y(n_538)
);

AND2x6_ASAP7_75t_L g539 ( 
.A(n_511),
.B(n_207),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_511),
.B(n_186),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_479),
.A2(n_403),
.B1(n_415),
.B2(n_201),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_511),
.A2(n_315),
.B1(n_371),
.B2(n_316),
.Y(n_542)
);

BUFx4f_ASAP7_75t_L g543 ( 
.A(n_494),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_442),
.A2(n_315),
.B1(n_281),
.B2(n_329),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_498),
.B(n_343),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_504),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_L g547 ( 
.A(n_498),
.B(n_392),
.C(n_391),
.Y(n_547)
);

OAI21xp33_ASAP7_75t_SL g548 ( 
.A1(n_442),
.A2(n_286),
.B(n_282),
.Y(n_548)
);

BUFx10_ASAP7_75t_L g549 ( 
.A(n_438),
.Y(n_549)
);

INVxp33_ASAP7_75t_L g550 ( 
.A(n_475),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_480),
.B(n_392),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_454),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_502),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_494),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_480),
.B(n_187),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_454),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_502),
.B(n_345),
.Y(n_557)
);

AO22x2_ASAP7_75t_L g558 ( 
.A1(n_462),
.A2(n_287),
.B1(n_341),
.B2(n_291),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_505),
.B(n_407),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_494),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_495),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_437),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_462),
.B(n_505),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_503),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_505),
.B(n_393),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_502),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_502),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_448),
.B(n_192),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_448),
.B(n_195),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_495),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_464),
.Y(n_571)
);

BUFx4f_ASAP7_75t_L g572 ( 
.A(n_503),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_467),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_478),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_464),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_439),
.B(n_393),
.Y(n_576)
);

OAI22xp33_ASAP7_75t_L g577 ( 
.A1(n_512),
.A2(n_304),
.B1(n_289),
.B2(n_348),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_456),
.B(n_197),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_464),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_509),
.B(n_401),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_477),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_503),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_503),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_495),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_454),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_503),
.Y(n_586)
);

BUFx4f_ASAP7_75t_L g587 ( 
.A(n_503),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_455),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_512),
.A2(n_298),
.B1(n_246),
.B2(n_283),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_495),
.A2(n_203),
.B1(n_317),
.B2(n_401),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_453),
.B(n_402),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_501),
.B(n_203),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_447),
.B(n_402),
.Y(n_593)
);

OR2x6_ASAP7_75t_L g594 ( 
.A(n_453),
.B(n_406),
.Y(n_594)
);

INVx6_ASAP7_75t_L g595 ( 
.A(n_501),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_456),
.B(n_204),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_477),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_461),
.B(n_209),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_501),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_461),
.B(n_216),
.Y(n_600)
);

INVxp33_ASAP7_75t_L g601 ( 
.A(n_443),
.Y(n_601)
);

INVx6_ASAP7_75t_L g602 ( 
.A(n_501),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_477),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_488),
.B(n_203),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_488),
.B(n_203),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_455),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_509),
.B(n_406),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_463),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_449),
.B(n_201),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_463),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_493),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_SL g612 ( 
.A(n_485),
.B(n_318),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_478),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_455),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_457),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_493),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_493),
.B(n_497),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_497),
.A2(n_203),
.B1(n_317),
.B2(n_428),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_497),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_457),
.Y(n_620)
);

INVxp33_ASAP7_75t_L g621 ( 
.A(n_510),
.Y(n_621)
);

INVx6_ASAP7_75t_L g622 ( 
.A(n_463),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_463),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_450),
.B(n_323),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_486),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_457),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_499),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_499),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_499),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_463),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_440),
.B(n_221),
.Y(n_631)
);

AND2x6_ASAP7_75t_L g632 ( 
.A(n_440),
.B(n_317),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_441),
.B(n_222),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_441),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_444),
.Y(n_635)
);

NOR2x1p5_ASAP7_75t_L g636 ( 
.A(n_459),
.B(n_193),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_460),
.B(n_317),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_470),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_463),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_444),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_446),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_446),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_513),
.Y(n_643)
);

NAND3xp33_ASAP7_75t_L g644 ( 
.A(n_472),
.B(n_264),
.C(n_263),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_469),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_465),
.B(n_317),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_469),
.Y(n_647)
);

AND2x2_ASAP7_75t_SL g648 ( 
.A(n_510),
.B(n_224),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_471),
.Y(n_649)
);

INVxp33_ASAP7_75t_L g650 ( 
.A(n_510),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_471),
.B(n_226),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_466),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_473),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_473),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_SL g655 ( 
.A(n_474),
.B(n_333),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_474),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_484),
.Y(n_657)
);

OA22x2_ASAP7_75t_L g658 ( 
.A1(n_514),
.A2(n_435),
.B1(n_430),
.B2(n_428),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_484),
.Y(n_659)
);

INVx4_ASAP7_75t_SL g660 ( 
.A(n_487),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_487),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_489),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_496),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_476),
.Y(n_664)
);

AO21x2_ASAP7_75t_L g665 ( 
.A1(n_490),
.A2(n_227),
.B(n_347),
.Y(n_665)
);

AND3x2_ASAP7_75t_L g666 ( 
.A(n_514),
.B(n_288),
.C(n_280),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_490),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_561),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_640),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_540),
.B(n_229),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_516),
.A2(n_514),
.B(n_242),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_530),
.B(n_238),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_519),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_524),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_621),
.B(n_249),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_621),
.B(n_251),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_640),
.Y(n_677)
);

O2A1O1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_545),
.A2(n_419),
.B(n_413),
.C(n_414),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_591),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_650),
.B(n_257),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_601),
.B(n_481),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_535),
.B(n_202),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_517),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_518),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_586),
.A2(n_261),
.B(n_344),
.Y(n_685)
);

NOR3xp33_ASAP7_75t_L g686 ( 
.A(n_612),
.B(n_419),
.C(n_430),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_561),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_562),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_574),
.A2(n_214),
.B1(n_210),
.B2(n_340),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_656),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_650),
.B(n_520),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_584),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_523),
.B(n_265),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_526),
.B(n_268),
.Y(n_694)
);

NOR3x1_ASAP7_75t_L g695 ( 
.A(n_574),
.B(n_418),
.C(n_423),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_584),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_537),
.B(n_413),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_524),
.Y(n_698)
);

O2A1O1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_545),
.A2(n_414),
.B(n_417),
.C(n_418),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_524),
.Y(n_700)
);

INVx5_ASAP7_75t_L g701 ( 
.A(n_539),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_601),
.B(n_202),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_515),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_599),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_599),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_576),
.B(n_210),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_528),
.B(n_533),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_536),
.B(n_303),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_568),
.B(n_569),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_648),
.B(n_314),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_648),
.B(n_324),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_578),
.B(n_212),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_580),
.Y(n_713)
);

NOR2xp67_ASAP7_75t_SL g714 ( 
.A(n_595),
.B(n_212),
.Y(n_714)
);

OR2x6_ASAP7_75t_L g715 ( 
.A(n_652),
.B(n_417),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_596),
.B(n_214),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_598),
.B(n_217),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_600),
.B(n_217),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_593),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_580),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_629),
.B(n_218),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_629),
.B(n_218),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_641),
.B(n_654),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_656),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_591),
.B(n_421),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_537),
.B(n_421),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_607),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_607),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_628),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_537),
.B(n_223),
.Y(n_730)
);

NOR3xp33_ASAP7_75t_L g731 ( 
.A(n_612),
.B(n_423),
.C(n_427),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_595),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_641),
.B(n_223),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_555),
.B(n_262),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_628),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_L g736 ( 
.A(n_539),
.B(n_262),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_609),
.B(n_273),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_641),
.B(n_273),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_654),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_563),
.B(n_290),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_522),
.B(n_427),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_525),
.Y(n_742)
);

XNOR2xp5_ASAP7_75t_L g743 ( 
.A(n_573),
.B(n_452),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_654),
.B(n_290),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_659),
.B(n_295),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_659),
.B(n_295),
.Y(n_746)
);

OR2x6_ASAP7_75t_L g747 ( 
.A(n_652),
.B(n_468),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_591),
.B(n_198),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_563),
.B(n_297),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_L g750 ( 
.A(n_539),
.B(n_297),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_563),
.B(n_644),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_665),
.A2(n_339),
.B1(n_342),
.B2(n_198),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_659),
.B(n_634),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_595),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_635),
.B(n_306),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_595),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_602),
.Y(n_757)
);

NOR3xp33_ASAP7_75t_L g758 ( 
.A(n_589),
.B(n_267),
.C(n_206),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_642),
.B(n_306),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_563),
.B(n_311),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_613),
.B(n_311),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_613),
.B(n_591),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_594),
.B(n_312),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_594),
.B(n_312),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_602),
.Y(n_765)
);

A2O1A1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_548),
.A2(n_313),
.B(n_325),
.C(n_338),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_521),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_532),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_602),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_602),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_645),
.B(n_313),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_532),
.Y(n_772)
);

NOR2xp67_ASAP7_75t_L g773 ( 
.A(n_562),
.B(n_325),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_538),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_515),
.B(n_327),
.Y(n_775)
);

AND2x6_ASAP7_75t_L g776 ( 
.A(n_553),
.B(n_566),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_647),
.B(n_327),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_594),
.B(n_336),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_567),
.A2(n_336),
.B(n_338),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_637),
.A2(n_340),
.B1(n_275),
.B2(n_330),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_522),
.B(n_491),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_573),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_538),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_515),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_SL g785 ( 
.A(n_549),
.B(n_506),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_541),
.B(n_275),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_542),
.B(n_275),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_665),
.A2(n_319),
.B1(n_208),
.B2(n_211),
.Y(n_788)
);

AOI221xp5_ASAP7_75t_L g789 ( 
.A1(n_577),
.A2(n_319),
.B1(n_208),
.B2(n_211),
.C(n_346),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_559),
.B(n_387),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_649),
.B(n_330),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_637),
.A2(n_646),
.B1(n_655),
.B2(n_636),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_653),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_594),
.B(n_206),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_649),
.B(n_330),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_657),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_646),
.B(n_219),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_667),
.B(n_387),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_551),
.B(n_219),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_649),
.B(n_389),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_565),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_649),
.B(n_661),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_552),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_661),
.B(n_389),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_638),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_661),
.B(n_390),
.Y(n_806)
);

INVxp67_ASAP7_75t_SL g807 ( 
.A(n_525),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_661),
.B(n_390),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_665),
.A2(n_346),
.B1(n_334),
.B2(n_332),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_655),
.A2(n_334),
.B1(n_332),
.B2(n_331),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_539),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_565),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_550),
.B(n_331),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_559),
.B(n_328),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_559),
.Y(n_815)
);

NOR2x1_ASAP7_75t_L g816 ( 
.A(n_547),
.B(n_328),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_552),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_590),
.A2(n_322),
.B1(n_320),
.B2(n_308),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_534),
.B(n_322),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_534),
.B(n_320),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_643),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_SL g822 ( 
.A1(n_638),
.A2(n_308),
.B1(n_307),
.B2(n_302),
.Y(n_822)
);

A2O1A1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_529),
.A2(n_307),
.B(n_302),
.C(n_278),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_556),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_529),
.A2(n_278),
.B(n_277),
.C(n_276),
.Y(n_825)
);

OR2x2_ASAP7_75t_L g826 ( 
.A(n_550),
.B(n_277),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_605),
.B(n_276),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_658),
.Y(n_828)
);

INVxp67_ASAP7_75t_SL g829 ( 
.A(n_525),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_544),
.A2(n_270),
.B1(n_169),
.B2(n_160),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_664),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_534),
.B(n_583),
.Y(n_832)
);

OAI221xp5_ASAP7_75t_L g833 ( 
.A1(n_570),
.A2(n_270),
.B1(n_9),
.B2(n_10),
.C(n_12),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_605),
.B(n_6),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_556),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_546),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_583),
.B(n_157),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_631),
.B(n_6),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_673),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_709),
.B(n_583),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_710),
.A2(n_633),
.B(n_651),
.C(n_592),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_710),
.A2(n_592),
.B(n_557),
.C(n_604),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_815),
.B(n_571),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_781),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_815),
.B(n_812),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_719),
.B(n_624),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_L g847 ( 
.A(n_682),
.B(n_663),
.C(n_662),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_802),
.A2(n_543),
.B(n_572),
.Y(n_848)
);

AO21x1_ASAP7_75t_L g849 ( 
.A1(n_834),
.A2(n_604),
.B(n_575),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_723),
.A2(n_543),
.B(n_587),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_683),
.B(n_625),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_742),
.A2(n_572),
.B(n_543),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_741),
.B(n_549),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_807),
.A2(n_572),
.B(n_587),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_801),
.B(n_579),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_684),
.B(n_549),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_829),
.A2(n_587),
.B(n_527),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_739),
.Y(n_858)
);

O2A1O1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_711),
.A2(n_617),
.B(n_603),
.C(n_581),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_792),
.B(n_546),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_674),
.B(n_660),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_784),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_832),
.A2(n_560),
.B(n_527),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_834),
.A2(n_531),
.B1(n_539),
.B2(n_597),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_698),
.B(n_546),
.Y(n_865)
);

OAI21xp33_ASAP7_75t_L g866 ( 
.A1(n_682),
.A2(n_558),
.B(n_658),
.Y(n_866)
);

BUFx4f_ASAP7_75t_L g867 ( 
.A(n_747),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_706),
.B(n_527),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_821),
.Y(n_869)
);

O2A1O1Ixp5_ASAP7_75t_L g870 ( 
.A1(n_672),
.A2(n_711),
.B(n_706),
.C(n_670),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_705),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_691),
.B(n_611),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_833),
.A2(n_619),
.B(n_616),
.C(n_627),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_669),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_832),
.A2(n_560),
.B(n_564),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_762),
.B(n_560),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_751),
.A2(n_539),
.B1(n_582),
.B2(n_564),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_799),
.B(n_813),
.Y(n_878)
);

OAI321xp33_ASAP7_75t_L g879 ( 
.A1(n_752),
.A2(n_558),
.A3(n_618),
.B1(n_588),
.B2(n_606),
.C(n_614),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_705),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_751),
.A2(n_582),
.B1(n_564),
.B2(n_639),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_753),
.A2(n_582),
.B(n_554),
.Y(n_882)
);

AOI21x1_ASAP7_75t_L g883 ( 
.A1(n_672),
.A2(n_615),
.B(n_614),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_821),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_705),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_831),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_754),
.A2(n_525),
.B(n_554),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_734),
.B(n_639),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_734),
.B(n_639),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_799),
.B(n_630),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_757),
.A2(n_525),
.B(n_554),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_828),
.B(n_558),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_SL g893 ( 
.A(n_782),
.B(n_666),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_797),
.A2(n_630),
.B(n_615),
.C(n_626),
.Y(n_894)
);

INVx4_ASAP7_75t_L g895 ( 
.A(n_705),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_765),
.A2(n_554),
.B(n_623),
.Y(n_896)
);

AOI221xp5_ASAP7_75t_L g897 ( 
.A1(n_752),
.A2(n_558),
.B1(n_606),
.B2(n_585),
.C(n_588),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_700),
.A2(n_630),
.B1(n_622),
.B2(n_554),
.Y(n_898)
);

O2A1O1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_823),
.A2(n_626),
.B(n_620),
.C(n_585),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_L g900 ( 
.A(n_702),
.B(n_623),
.C(n_620),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_769),
.A2(n_623),
.B(n_608),
.Y(n_901)
);

OA22x2_ASAP7_75t_L g902 ( 
.A1(n_810),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_R g903 ( 
.A(n_688),
.B(n_110),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_713),
.B(n_610),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_770),
.A2(n_608),
.B(n_610),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_SL g906 ( 
.A1(n_837),
.A2(n_766),
.B(n_825),
.C(n_786),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_669),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_677),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_756),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_838),
.A2(n_660),
.B(n_19),
.C(n_20),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_756),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_720),
.B(n_610),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_727),
.B(n_610),
.Y(n_913)
);

O2A1O1Ixp5_ASAP7_75t_L g914 ( 
.A1(n_707),
.A2(n_660),
.B(n_632),
.C(n_622),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_826),
.B(n_17),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_728),
.B(n_610),
.Y(n_916)
);

BUFx8_ASAP7_75t_L g917 ( 
.A(n_836),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_788),
.A2(n_622),
.B1(n_608),
.B2(n_22),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_732),
.A2(n_608),
.B(n_622),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_788),
.A2(n_17),
.B1(n_20),
.B2(n_22),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_690),
.Y(n_921)
);

NOR2x1_ASAP7_75t_L g922 ( 
.A(n_836),
.B(n_660),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_690),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_SL g924 ( 
.A1(n_837),
.A2(n_632),
.B(n_25),
.C(n_28),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_793),
.B(n_632),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_732),
.A2(n_632),
.B(n_151),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_762),
.B(n_24),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_701),
.A2(n_632),
.B(n_131),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_724),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_809),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_701),
.A2(n_632),
.B(n_130),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_701),
.A2(n_124),
.B(n_123),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_838),
.A2(n_30),
.B(n_31),
.C(n_33),
.Y(n_933)
);

INVx1_ASAP7_75t_SL g934 ( 
.A(n_831),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_701),
.A2(n_111),
.B(n_107),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_721),
.A2(n_100),
.B(n_96),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_SL g937 ( 
.A(n_805),
.B(n_93),
.Y(n_937)
);

NOR2xp67_ASAP7_75t_L g938 ( 
.A(n_773),
.B(n_92),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_722),
.A2(n_78),
.B(n_73),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_697),
.B(n_65),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_827),
.A2(n_33),
.B1(n_34),
.B2(n_40),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_733),
.A2(n_71),
.B(n_41),
.Y(n_942)
);

NOR2x1_ASAP7_75t_L g943 ( 
.A(n_681),
.B(n_34),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_796),
.Y(n_944)
);

NOR2x1_ASAP7_75t_L g945 ( 
.A(n_715),
.B(n_44),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_671),
.A2(n_45),
.B(n_46),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_729),
.A2(n_735),
.B(n_768),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_738),
.A2(n_51),
.B(n_53),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_747),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_814),
.A2(n_55),
.B(n_58),
.C(n_60),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_761),
.B(n_58),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_715),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_729),
.A2(n_735),
.B(n_803),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_811),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_744),
.A2(n_60),
.B(n_61),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_726),
.B(n_62),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_745),
.A2(n_64),
.B(n_746),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_675),
.A2(n_64),
.B(n_676),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_668),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_703),
.B(n_790),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_813),
.B(n_715),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_779),
.A2(n_680),
.B(n_827),
.C(n_686),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_747),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_731),
.A2(n_717),
.B(n_716),
.C(n_712),
.Y(n_964)
);

NAND3xp33_ASAP7_75t_L g965 ( 
.A(n_797),
.B(n_761),
.C(n_809),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_687),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_819),
.A2(n_820),
.B(n_704),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_692),
.A2(n_696),
.B(n_800),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_804),
.A2(n_806),
.B(n_808),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_718),
.B(n_790),
.Y(n_970)
);

NOR2xp67_ASAP7_75t_L g971 ( 
.A(n_743),
.B(n_780),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_689),
.A2(n_725),
.B1(n_679),
.B2(n_749),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_767),
.A2(n_772),
.B(n_817),
.Y(n_973)
);

AOI21x1_ASAP7_75t_L g974 ( 
.A1(n_767),
.A2(n_772),
.B(n_817),
.Y(n_974)
);

AO32x1_ASAP7_75t_L g975 ( 
.A1(n_830),
.A2(n_768),
.A3(n_803),
.B1(n_783),
.B2(n_774),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_774),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_783),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_835),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_693),
.B(n_694),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_835),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_708),
.B(n_824),
.Y(n_981)
);

BUFx4f_ASAP7_75t_L g982 ( 
.A(n_748),
.Y(n_982)
);

AOI22x1_ASAP7_75t_L g983 ( 
.A1(n_811),
.A2(n_824),
.B1(n_685),
.B2(n_794),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_798),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_776),
.B(n_740),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_736),
.A2(n_750),
.B(n_771),
.Y(n_986)
);

AOI21x1_ASAP7_75t_L g987 ( 
.A1(n_714),
.A2(n_777),
.B(n_759),
.Y(n_987)
);

CKINVDCx8_ASAP7_75t_R g988 ( 
.A(n_763),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_SL g989 ( 
.A1(n_791),
.A2(n_795),
.B(n_737),
.C(n_730),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_755),
.A2(n_791),
.B(n_795),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_740),
.B(n_760),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_775),
.A2(n_811),
.B(n_787),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_749),
.B(n_760),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_776),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_811),
.A2(n_678),
.B(n_699),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_776),
.Y(n_996)
);

AO21x1_ASAP7_75t_L g997 ( 
.A1(n_763),
.A2(n_764),
.B(n_778),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_776),
.B(n_764),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_778),
.A2(n_816),
.B(n_776),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_822),
.B(n_785),
.Y(n_1000)
);

NAND2x1_ASAP7_75t_L g1001 ( 
.A(n_758),
.B(n_818),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_695),
.Y(n_1002)
);

OR2x6_ASAP7_75t_L g1003 ( 
.A(n_789),
.B(n_821),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_802),
.A2(n_572),
.B(n_543),
.Y(n_1004)
);

NOR2xp67_ASAP7_75t_L g1005 ( 
.A(n_688),
.B(n_652),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_828),
.A2(n_752),
.B1(n_809),
.B2(n_788),
.Y(n_1006)
);

AND2x6_ASAP7_75t_L g1007 ( 
.A(n_811),
.B(n_828),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_802),
.A2(n_572),
.B(n_543),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_815),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_802),
.A2(n_572),
.B(n_543),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_815),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_705),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_709),
.B(n_815),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_802),
.A2(n_572),
.B(n_543),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_673),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_709),
.B(n_815),
.Y(n_1016)
);

AND2x2_ASAP7_75t_SL g1017 ( 
.A(n_785),
.B(n_664),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_828),
.A2(n_709),
.B(n_723),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_709),
.B(n_815),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_802),
.A2(n_572),
.B(n_543),
.Y(n_1020)
);

NOR2xp67_ASAP7_75t_L g1021 ( 
.A(n_688),
.B(n_652),
.Y(n_1021)
);

NOR2xp67_ASAP7_75t_L g1022 ( 
.A(n_688),
.B(n_652),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_710),
.A2(n_711),
.B(n_834),
.C(n_709),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_705),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_802),
.A2(n_572),
.B(n_543),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_739),
.Y(n_1026)
);

AOI21x1_ASAP7_75t_L g1027 ( 
.A1(n_974),
.A2(n_1004),
.B(n_848),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_944),
.Y(n_1028)
);

AND2x2_ASAP7_75t_SL g1029 ( 
.A(n_878),
.B(n_1017),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_839),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_874),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1013),
.B(n_1016),
.Y(n_1032)
);

AOI21x1_ASAP7_75t_L g1033 ( 
.A1(n_1008),
.A2(n_1014),
.B(n_1010),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_929),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1013),
.B(n_1016),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_869),
.Y(n_1036)
);

AO31x2_ASAP7_75t_L g1037 ( 
.A1(n_849),
.A2(n_997),
.A3(n_894),
.B(n_918),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_1019),
.A2(n_840),
.B(n_986),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_984),
.B(n_868),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_969),
.A2(n_979),
.B(n_1023),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_993),
.A2(n_961),
.B1(n_846),
.B2(n_853),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_857),
.A2(n_850),
.B(n_1020),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_970),
.B(n_872),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_1025),
.A2(n_854),
.B(n_852),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_851),
.B(n_951),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_1015),
.Y(n_1046)
);

AOI21x1_ASAP7_75t_SL g1047 ( 
.A1(n_985),
.A2(n_998),
.B(n_940),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_888),
.A2(n_889),
.B(n_882),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_844),
.B(n_886),
.Y(n_1049)
);

NOR2x1_ASAP7_75t_L g1050 ( 
.A(n_1005),
.B(n_1021),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_967),
.A2(n_981),
.B(n_990),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1018),
.B(n_845),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_934),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1018),
.B(n_845),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_907),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_908),
.Y(n_1056)
);

AOI21xp33_ASAP7_75t_L g1057 ( 
.A1(n_962),
.A2(n_1006),
.B(n_1001),
.Y(n_1057)
);

NAND2x1p5_ASAP7_75t_L g1058 ( 
.A(n_895),
.B(n_880),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_SL g1059 ( 
.A1(n_1000),
.A2(n_1006),
.B(n_847),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_883),
.A2(n_983),
.B(n_953),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_927),
.A2(n_930),
.B(n_920),
.C(n_866),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_947),
.A2(n_953),
.B(n_987),
.Y(n_1062)
);

AOI21x1_ASAP7_75t_L g1063 ( 
.A1(n_890),
.A2(n_999),
.B(n_968),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_863),
.A2(n_875),
.B(n_876),
.Y(n_1064)
);

XNOR2xp5_ASAP7_75t_L g1065 ( 
.A(n_971),
.B(n_1022),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_SL g1066 ( 
.A1(n_920),
.A2(n_930),
.B(n_941),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_842),
.A2(n_940),
.B(n_843),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_880),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_956),
.B(n_855),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_985),
.A2(n_860),
.B1(n_909),
.B2(n_1011),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_964),
.B(n_870),
.Y(n_1071)
);

AOI21x1_ASAP7_75t_L g1072 ( 
.A1(n_887),
.A2(n_891),
.B(n_896),
.Y(n_1072)
);

BUFx2_ASAP7_75t_SL g1073 ( 
.A(n_884),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_956),
.B(n_855),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_947),
.A2(n_973),
.B(n_899),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_841),
.A2(n_995),
.B(n_859),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_856),
.B(n_982),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_880),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_914),
.A2(n_892),
.B(n_877),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_946),
.A2(n_918),
.B(n_933),
.C(n_892),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_905),
.A2(n_901),
.B(n_992),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_989),
.A2(n_904),
.B(n_912),
.Y(n_1082)
);

INVx2_ASAP7_75t_SL g1083 ( 
.A(n_1002),
.Y(n_1083)
);

AOI21xp33_ASAP7_75t_L g1084 ( 
.A1(n_972),
.A2(n_1003),
.B(n_952),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_862),
.B(n_959),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_SL g1086 ( 
.A1(n_895),
.A2(n_885),
.B(n_954),
.Y(n_1086)
);

AO31x2_ASAP7_75t_L g1087 ( 
.A1(n_957),
.A2(n_958),
.A3(n_948),
.B(n_955),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_929),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_904),
.A2(n_916),
.B(n_913),
.Y(n_1089)
);

AO31x2_ASAP7_75t_L g1090 ( 
.A1(n_942),
.A2(n_975),
.A3(n_923),
.B(n_921),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_994),
.A2(n_996),
.B(n_919),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_966),
.B(n_912),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_913),
.A2(n_916),
.B(n_909),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_871),
.B(n_1024),
.Y(n_1094)
);

AOI21x1_ASAP7_75t_SL g1095 ( 
.A1(n_925),
.A2(n_975),
.B(n_906),
.Y(n_1095)
);

NOR2xp67_ASAP7_75t_SL g1096 ( 
.A(n_988),
.B(n_885),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_917),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_864),
.A2(n_858),
.B(n_1026),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_879),
.A2(n_881),
.B(n_1009),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_960),
.A2(n_1024),
.B(n_1012),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_871),
.A2(n_1012),
.B(n_900),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_911),
.B(n_897),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_976),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_977),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_978),
.A2(n_980),
.B(n_939),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_873),
.A2(n_898),
.B(n_946),
.Y(n_1106)
);

AOI221xp5_ASAP7_75t_L g1107 ( 
.A1(n_972),
.A2(n_950),
.B1(n_915),
.B2(n_963),
.C(n_910),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1007),
.Y(n_1108)
);

NAND2x1p5_ASAP7_75t_L g1109 ( 
.A(n_885),
.B(n_954),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_SL g1110 ( 
.A1(n_954),
.A2(n_861),
.B(n_911),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_982),
.B(n_1003),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_936),
.A2(n_922),
.B(n_932),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_935),
.A2(n_926),
.B(n_928),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1007),
.A2(n_938),
.B(n_861),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_911),
.A2(n_975),
.B(n_865),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_931),
.A2(n_943),
.B(n_945),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1007),
.B(n_1003),
.Y(n_1117)
);

NOR3xp33_ASAP7_75t_L g1118 ( 
.A(n_949),
.B(n_924),
.C(n_867),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_902),
.A2(n_1007),
.B(n_867),
.Y(n_1119)
);

NAND2x1p5_ASAP7_75t_L g1120 ( 
.A(n_1007),
.B(n_917),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_902),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_903),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_937),
.A2(n_883),
.B(n_974),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_893),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_974),
.Y(n_1125)
);

BUFx10_ASAP7_75t_L g1126 ( 
.A(n_851),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1013),
.A2(n_1019),
.B(n_1016),
.Y(n_1127)
);

OAI22x1_ASAP7_75t_L g1128 ( 
.A1(n_1000),
.A2(n_965),
.B1(n_792),
.B2(n_878),
.Y(n_1128)
);

AOI21x1_ASAP7_75t_SL g1129 ( 
.A1(n_985),
.A2(n_998),
.B(n_940),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1013),
.A2(n_1019),
.B(n_1016),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_965),
.A2(n_1013),
.B1(n_1019),
.B2(n_1016),
.Y(n_1131)
);

INVx2_ASAP7_75t_SL g1132 ( 
.A(n_839),
.Y(n_1132)
);

NAND2x1p5_ASAP7_75t_L g1133 ( 
.A(n_895),
.B(n_880),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_974),
.A2(n_883),
.B(n_848),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_974),
.A2(n_883),
.B(n_848),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_SL g1136 ( 
.A1(n_1023),
.A2(n_1016),
.B(n_1013),
.Y(n_1136)
);

NAND2x1_ASAP7_75t_L g1137 ( 
.A(n_1007),
.B(n_895),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_974),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_878),
.B(n_853),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_954),
.Y(n_1140)
);

AND2x6_ASAP7_75t_L g1141 ( 
.A(n_994),
.B(n_996),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_878),
.B(n_1013),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_965),
.A2(n_1023),
.B(n_951),
.C(n_878),
.Y(n_1143)
);

AOI21xp33_ASAP7_75t_L g1144 ( 
.A1(n_965),
.A2(n_682),
.B(n_535),
.Y(n_1144)
);

AOI21x1_ASAP7_75t_L g1145 ( 
.A1(n_974),
.A2(n_1004),
.B(n_848),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1023),
.A2(n_870),
.B(n_1018),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1023),
.A2(n_870),
.B(n_1018),
.Y(n_1147)
);

AOI221xp5_ASAP7_75t_SL g1148 ( 
.A1(n_1006),
.A2(n_930),
.B1(n_920),
.B2(n_866),
.C(n_951),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_911),
.B(n_862),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_944),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1023),
.A2(n_870),
.B(n_1018),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_849),
.A2(n_997),
.A3(n_894),
.B(n_918),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_883),
.A2(n_974),
.B(n_953),
.Y(n_1153)
);

NAND2xp33_ASAP7_75t_SL g1154 ( 
.A(n_991),
.B(n_878),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1013),
.A2(n_1019),
.B(n_1016),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_965),
.A2(n_1023),
.B(n_951),
.C(n_878),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_878),
.B(n_1013),
.Y(n_1157)
);

AOI21x1_ASAP7_75t_SL g1158 ( 
.A1(n_985),
.A2(n_998),
.B(n_940),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_878),
.B(n_1013),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_883),
.A2(n_974),
.B(n_953),
.Y(n_1160)
);

AOI221x1_ASAP7_75t_L g1161 ( 
.A1(n_965),
.A2(n_951),
.B1(n_991),
.B2(n_918),
.C(n_946),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_880),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_880),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_869),
.Y(n_1164)
);

INVx2_ASAP7_75t_SL g1165 ( 
.A(n_839),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_993),
.A2(n_878),
.B1(n_682),
.B2(n_991),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_944),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_944),
.Y(n_1168)
);

AO21x1_ASAP7_75t_L g1169 ( 
.A1(n_1023),
.A2(n_951),
.B(n_918),
.Y(n_1169)
);

NAND2x1p5_ASAP7_75t_L g1170 ( 
.A(n_895),
.B(n_880),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_974),
.A2(n_883),
.B(n_848),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_839),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_839),
.Y(n_1173)
);

AOI21x1_ASAP7_75t_L g1174 ( 
.A1(n_974),
.A2(n_1004),
.B(n_848),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_878),
.B(n_683),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_878),
.B(n_853),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_878),
.B(n_1013),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_993),
.A2(n_878),
.B1(n_682),
.B2(n_991),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1040),
.A2(n_1064),
.B(n_1051),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1028),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1045),
.A2(n_1144),
.B(n_1059),
.C(n_1143),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1128),
.A2(n_1084),
.B1(n_1169),
.B2(n_1176),
.Y(n_1182)
);

OAI21xp33_ASAP7_75t_L g1183 ( 
.A1(n_1166),
.A2(n_1178),
.B(n_1175),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1067),
.A2(n_1136),
.B(n_1038),
.Y(n_1184)
);

BUFx4_ASAP7_75t_SL g1185 ( 
.A(n_1097),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1140),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1142),
.B(n_1157),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1048),
.A2(n_1076),
.B(n_1071),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1083),
.B(n_1149),
.Y(n_1189)
);

CKINVDCx20_ASAP7_75t_R g1190 ( 
.A(n_1065),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1149),
.B(n_1111),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1149),
.B(n_1050),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1159),
.B(n_1177),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1069),
.B(n_1074),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1043),
.B(n_1032),
.Y(n_1195)
);

AOI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1071),
.A2(n_1145),
.B(n_1027),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1035),
.B(n_1175),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_1097),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1164),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1127),
.A2(n_1155),
.B(n_1130),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1139),
.A2(n_1029),
.B1(n_1057),
.B2(n_1107),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1143),
.A2(n_1156),
.B(n_1061),
.C(n_1066),
.Y(n_1202)
);

NAND2x1p5_ASAP7_75t_L g1203 ( 
.A(n_1163),
.B(n_1096),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1147),
.A2(n_1151),
.B(n_1042),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1029),
.B(n_1077),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1041),
.B(n_1126),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1156),
.A2(n_1061),
.B(n_1080),
.C(n_1124),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1150),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1039),
.A2(n_1044),
.B(n_1106),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1126),
.B(n_1053),
.Y(n_1210)
);

NAND2xp33_ASAP7_75t_L g1211 ( 
.A(n_1120),
.B(n_1117),
.Y(n_1211)
);

INVx4_ASAP7_75t_L g1212 ( 
.A(n_1140),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1030),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1148),
.B(n_1052),
.Y(n_1214)
);

BUFx10_ASAP7_75t_L g1215 ( 
.A(n_1122),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1062),
.A2(n_1060),
.B(n_1075),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1049),
.B(n_1173),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1132),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1154),
.A2(n_1118),
.B1(n_1172),
.B2(n_1165),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1036),
.Y(n_1220)
);

AND2x2_ASAP7_75t_SL g1221 ( 
.A(n_1121),
.B(n_1118),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1073),
.Y(n_1222)
);

BUFx4_ASAP7_75t_SL g1223 ( 
.A(n_1167),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1168),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1036),
.Y(n_1225)
);

INVxp67_ASAP7_75t_L g1226 ( 
.A(n_1046),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1046),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1054),
.B(n_1131),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1154),
.A2(n_1173),
.B1(n_1102),
.B2(n_1085),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1082),
.A2(n_1114),
.B(n_1093),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1068),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1120),
.Y(n_1232)
);

AOI21xp33_ASAP7_75t_L g1233 ( 
.A1(n_1080),
.A2(n_1070),
.B(n_1099),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1089),
.A2(n_1079),
.B(n_1086),
.Y(n_1234)
);

NAND2x1p5_ASAP7_75t_L g1235 ( 
.A(n_1163),
.B(n_1140),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1121),
.A2(n_1119),
.B1(n_1104),
.B2(n_1031),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1161),
.A2(n_1081),
.B(n_1110),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1068),
.B(n_1078),
.Y(n_1238)
);

INVx3_ASAP7_75t_SL g1239 ( 
.A(n_1078),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1092),
.B(n_1103),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1162),
.B(n_1108),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1141),
.A2(n_1055),
.B1(n_1056),
.B2(n_1116),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1034),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1088),
.A2(n_1141),
.B1(n_1162),
.B2(n_1094),
.Y(n_1244)
);

BUFx10_ASAP7_75t_L g1245 ( 
.A(n_1141),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1125),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1141),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1087),
.B(n_1170),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1100),
.B(n_1091),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1109),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1141),
.Y(n_1251)
);

OR2x6_ASAP7_75t_L g1252 ( 
.A(n_1058),
.B(n_1133),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1081),
.A2(n_1060),
.B(n_1112),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1109),
.Y(n_1254)
);

AND2x6_ASAP7_75t_SL g1255 ( 
.A(n_1058),
.B(n_1170),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1087),
.B(n_1133),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1101),
.A2(n_1062),
.B(n_1105),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1087),
.Y(n_1258)
);

AOI21x1_ASAP7_75t_SL g1259 ( 
.A1(n_1047),
.A2(n_1129),
.B(n_1158),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1037),
.B(n_1152),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1087),
.B(n_1037),
.Y(n_1261)
);

NOR2x1p5_ASAP7_75t_SL g1262 ( 
.A(n_1174),
.B(n_1033),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1037),
.B(n_1152),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1105),
.A2(n_1123),
.B(n_1138),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1091),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1037),
.B(n_1152),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1098),
.B(n_1152),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1115),
.B(n_1098),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1090),
.B(n_1160),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1090),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1090),
.Y(n_1271)
);

INVxp67_ASAP7_75t_SL g1272 ( 
.A(n_1153),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1063),
.B(n_1171),
.Y(n_1273)
);

BUFx4_ASAP7_75t_SL g1274 ( 
.A(n_1047),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1134),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1113),
.A2(n_1135),
.B(n_1171),
.Y(n_1276)
);

BUFx8_ASAP7_75t_SL g1277 ( 
.A(n_1072),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1113),
.A2(n_1129),
.B(n_1158),
.Y(n_1278)
);

BUFx5_ASAP7_75t_L g1279 ( 
.A(n_1095),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1095),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1142),
.B(n_1157),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1142),
.B(n_1157),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1137),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1083),
.B(n_1149),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1045),
.B(n_719),
.Y(n_1285)
);

AOI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1045),
.A2(n_535),
.B1(n_682),
.B2(n_351),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1144),
.A2(n_965),
.B1(n_682),
.B2(n_1045),
.Y(n_1287)
);

INVx3_ASAP7_75t_SL g1288 ( 
.A(n_1097),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1045),
.A2(n_1144),
.B(n_682),
.C(n_1059),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1139),
.B(n_1176),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1142),
.B(n_1157),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1040),
.A2(n_1064),
.B(n_1067),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1061),
.A2(n_1045),
.B1(n_1066),
.B2(n_965),
.Y(n_1293)
);

CKINVDCx8_ASAP7_75t_R g1294 ( 
.A(n_1073),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1144),
.A2(n_965),
.B1(n_682),
.B2(n_1045),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1137),
.B(n_895),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1083),
.B(n_1149),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1097),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1142),
.B(n_1157),
.Y(n_1299)
);

INVx2_ASAP7_75t_SL g1300 ( 
.A(n_1049),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1142),
.B(n_1157),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1083),
.B(n_1149),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1061),
.A2(n_1045),
.B1(n_1066),
.B2(n_965),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1164),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1083),
.B(n_1149),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1083),
.B(n_1149),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1137),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1040),
.A2(n_1064),
.B(n_1051),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1028),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1040),
.A2(n_1064),
.B(n_1051),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1061),
.A2(n_1045),
.B1(n_1066),
.B2(n_965),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1040),
.A2(n_1064),
.B(n_1051),
.Y(n_1312)
);

AO21x1_ASAP7_75t_L g1313 ( 
.A1(n_1144),
.A2(n_1154),
.B(n_1057),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1083),
.B(n_1149),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1046),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1164),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1028),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1028),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1061),
.A2(n_1045),
.B1(n_1066),
.B2(n_965),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1028),
.Y(n_1320)
);

BUFx10_ASAP7_75t_L g1321 ( 
.A(n_1124),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1040),
.A2(n_1064),
.B(n_1051),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1140),
.Y(n_1323)
);

AO21x2_ASAP7_75t_L g1324 ( 
.A1(n_1076),
.A2(n_1071),
.B(n_1146),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1142),
.B(n_1157),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1142),
.B(n_1157),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1185),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1246),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1286),
.A2(n_1285),
.B1(n_1195),
.B2(n_1201),
.Y(n_1329)
);

BUFx12f_ASAP7_75t_L g1330 ( 
.A(n_1198),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1188),
.A2(n_1292),
.B(n_1179),
.Y(n_1331)
);

INVx6_ASAP7_75t_L g1332 ( 
.A(n_1255),
.Y(n_1332)
);

BUFx4f_ASAP7_75t_L g1333 ( 
.A(n_1203),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1298),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1195),
.A2(n_1287),
.B1(n_1295),
.B2(n_1194),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1187),
.B(n_1193),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1293),
.A2(n_1303),
.B1(n_1311),
.B2(n_1319),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1180),
.Y(n_1338)
);

AO21x1_ASAP7_75t_SL g1339 ( 
.A1(n_1233),
.A2(n_1263),
.B(n_1260),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1208),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1247),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1227),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_1190),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1220),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1293),
.A2(n_1319),
.B1(n_1303),
.B2(n_1311),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1183),
.A2(n_1206),
.B1(n_1290),
.B2(n_1205),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1315),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1248),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1194),
.B(n_1197),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1247),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1224),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1191),
.A2(n_1210),
.B1(n_1197),
.B2(n_1192),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1264),
.A2(n_1276),
.B(n_1253),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1240),
.A2(n_1219),
.B1(n_1229),
.B2(n_1182),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1300),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1199),
.Y(n_1356)
);

AO21x1_ASAP7_75t_L g1357 ( 
.A1(n_1289),
.A2(n_1181),
.B(n_1233),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1191),
.A2(n_1192),
.B1(n_1221),
.B2(n_1211),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1187),
.A2(n_1326),
.B1(n_1282),
.B2(n_1291),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1193),
.B(n_1281),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1309),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1317),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1318),
.Y(n_1363)
);

CKINVDCx6p67_ASAP7_75t_R g1364 ( 
.A(n_1288),
.Y(n_1364)
);

BUFx4f_ASAP7_75t_L g1365 ( 
.A(n_1203),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1281),
.A2(n_1326),
.B1(n_1282),
.B2(n_1299),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1291),
.B(n_1299),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1247),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_SL g1369 ( 
.A1(n_1321),
.A2(n_1234),
.B1(n_1247),
.B2(n_1325),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1320),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1243),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1179),
.A2(n_1312),
.B(n_1310),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1275),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1241),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1241),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1257),
.A2(n_1259),
.B(n_1196),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1232),
.B(n_1189),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1207),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1225),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1308),
.A2(n_1322),
.B(n_1310),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1294),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1308),
.A2(n_1322),
.B(n_1312),
.Y(n_1382)
);

INVx4_ASAP7_75t_L g1383 ( 
.A(n_1252),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1245),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1301),
.B(n_1325),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1186),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1186),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1321),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1213),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1313),
.A2(n_1301),
.B1(n_1277),
.B2(n_1324),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1324),
.A2(n_1256),
.B1(n_1217),
.B2(n_1214),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1214),
.A2(n_1316),
.B1(n_1304),
.B2(n_1228),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1184),
.A2(n_1230),
.B(n_1237),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1200),
.A2(n_1204),
.B(n_1209),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1254),
.Y(n_1395)
);

NAND2x1p5_ASAP7_75t_L g1396 ( 
.A(n_1242),
.B(n_1265),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1251),
.A2(n_1228),
.B1(n_1305),
.B2(n_1297),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1226),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1284),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1297),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1261),
.A2(n_1302),
.B1(n_1314),
.B2(n_1306),
.Y(n_1401)
);

BUFx12f_ASAP7_75t_L g1402 ( 
.A(n_1215),
.Y(n_1402)
);

BUFx10_ASAP7_75t_L g1403 ( 
.A(n_1222),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1302),
.A2(n_1305),
.B1(n_1314),
.B2(n_1306),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1258),
.A2(n_1236),
.B1(n_1267),
.B2(n_1218),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1202),
.A2(n_1231),
.B1(n_1250),
.B2(n_1215),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1267),
.Y(n_1407)
);

AO21x2_ASAP7_75t_L g1408 ( 
.A1(n_1268),
.A2(n_1273),
.B(n_1269),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1280),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1244),
.A2(n_1238),
.B1(n_1250),
.B2(n_1252),
.Y(n_1410)
);

AO21x1_ASAP7_75t_L g1411 ( 
.A1(n_1260),
.A2(n_1266),
.B(n_1263),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1238),
.B(n_1239),
.Y(n_1412)
);

BUFx10_ASAP7_75t_L g1413 ( 
.A(n_1252),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1283),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1272),
.Y(n_1415)
);

BUFx2_ASAP7_75t_SL g1416 ( 
.A(n_1212),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1323),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1266),
.A2(n_1279),
.B1(n_1249),
.B2(n_1270),
.Y(n_1418)
);

OAI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1223),
.A2(n_1307),
.B1(n_1283),
.B2(n_1296),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_1323),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1212),
.B(n_1235),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1279),
.A2(n_1249),
.B1(n_1268),
.B2(n_1307),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1278),
.A2(n_1269),
.B(n_1296),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1235),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1216),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1274),
.Y(n_1426)
);

OAI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1271),
.A2(n_1216),
.B1(n_1262),
.B2(n_1279),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1279),
.A2(n_1017),
.B1(n_1029),
.B2(n_1045),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1293),
.A2(n_1144),
.B1(n_965),
.B2(n_682),
.Y(n_1429)
);

CKINVDCx6p67_ASAP7_75t_R g1430 ( 
.A(n_1288),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_SL g1431 ( 
.A1(n_1286),
.A2(n_1000),
.B1(n_1017),
.B2(n_988),
.Y(n_1431)
);

AOI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1276),
.A2(n_1071),
.B(n_1196),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_SL g1433 ( 
.A1(n_1286),
.A2(n_1000),
.B1(n_1017),
.B2(n_988),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1191),
.B(n_1192),
.Y(n_1434)
);

NAND2x1p5_ASAP7_75t_L g1435 ( 
.A(n_1247),
.B(n_1248),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1247),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1180),
.Y(n_1437)
);

BUFx8_ASAP7_75t_SL g1438 ( 
.A(n_1198),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1286),
.A2(n_535),
.B1(n_682),
.B2(n_489),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1187),
.B(n_1325),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1286),
.A2(n_1045),
.B1(n_1285),
.B2(n_682),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1180),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1191),
.B(n_1192),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1247),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1227),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1180),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1247),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1187),
.B(n_1325),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1373),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1348),
.B(n_1337),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1344),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1344),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1408),
.B(n_1348),
.Y(n_1453)
);

AO21x1_ASAP7_75t_SL g1454 ( 
.A1(n_1345),
.A2(n_1390),
.B(n_1429),
.Y(n_1454)
);

OR2x6_ASAP7_75t_L g1455 ( 
.A(n_1393),
.B(n_1435),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1425),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1408),
.B(n_1391),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1411),
.Y(n_1458)
);

CKINVDCx16_ASAP7_75t_R g1459 ( 
.A(n_1330),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1336),
.B(n_1367),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1425),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_1355),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1411),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1407),
.B(n_1383),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1380),
.A2(n_1382),
.B(n_1394),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1440),
.B(n_1448),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1440),
.B(n_1448),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1408),
.B(n_1396),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1413),
.Y(n_1469)
);

INVxp67_ASAP7_75t_SL g1470 ( 
.A(n_1347),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1441),
.A2(n_1439),
.B(n_1329),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1435),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1342),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1339),
.B(n_1418),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1353),
.A2(n_1432),
.B(n_1376),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1328),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1415),
.Y(n_1477)
);

INVx2_ASAP7_75t_SL g1478 ( 
.A(n_1413),
.Y(n_1478)
);

OR2x6_ASAP7_75t_L g1479 ( 
.A(n_1435),
.B(n_1396),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1360),
.B(n_1385),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1423),
.A2(n_1372),
.B(n_1331),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1409),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1332),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1371),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1338),
.Y(n_1485)
);

BUFx2_ASAP7_75t_SL g1486 ( 
.A(n_1388),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1340),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1351),
.Y(n_1488)
);

INVx2_ASAP7_75t_SL g1489 ( 
.A(n_1413),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1341),
.A2(n_1447),
.B(n_1444),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1383),
.B(n_1436),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1389),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1361),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1445),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1362),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1363),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1378),
.B(n_1357),
.Y(n_1497)
);

OA21x2_ASAP7_75t_L g1498 ( 
.A1(n_1422),
.A2(n_1405),
.B(n_1354),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1370),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1359),
.B(n_1366),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1437),
.B(n_1442),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1350),
.B(n_1368),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1350),
.B(n_1368),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1446),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1431),
.A2(n_1433),
.B1(n_1335),
.B2(n_1332),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1346),
.B(n_1349),
.Y(n_1506)
);

BUFx4f_ASAP7_75t_SL g1507 ( 
.A(n_1330),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1398),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1343),
.B(n_1443),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1392),
.B(n_1352),
.Y(n_1510)
);

OR2x6_ASAP7_75t_L g1511 ( 
.A(n_1368),
.B(n_1332),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1428),
.A2(n_1397),
.B1(n_1406),
.B2(n_1332),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1427),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1398),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1460),
.B(n_1401),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1453),
.B(n_1395),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1460),
.B(n_1369),
.Y(n_1517)
);

INVxp67_ASAP7_75t_L g1518 ( 
.A(n_1473),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1453),
.B(n_1388),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1466),
.B(n_1358),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1449),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1466),
.B(n_1443),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1449),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1467),
.B(n_1379),
.Y(n_1524)
);

INVxp67_ASAP7_75t_R g1525 ( 
.A(n_1490),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1457),
.B(n_1426),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1474),
.B(n_1434),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1474),
.B(n_1434),
.Y(n_1528)
);

OAI321xp33_ASAP7_75t_L g1529 ( 
.A1(n_1471),
.A2(n_1419),
.A3(n_1410),
.B1(n_1404),
.B2(n_1375),
.C(n_1374),
.Y(n_1529)
);

INVx4_ASAP7_75t_L g1530 ( 
.A(n_1511),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1472),
.B(n_1414),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1480),
.B(n_1399),
.Y(n_1532)
);

OAI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1505),
.A2(n_1333),
.B1(n_1365),
.B2(n_1356),
.C(n_1412),
.Y(n_1533)
);

AND2x4_ASAP7_75t_SL g1534 ( 
.A(n_1479),
.B(n_1384),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1456),
.Y(n_1535)
);

AO31x2_ASAP7_75t_L g1536 ( 
.A1(n_1458),
.A2(n_1387),
.A3(n_1386),
.B(n_1400),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1468),
.B(n_1356),
.Y(n_1537)
);

INVx5_ASAP7_75t_L g1538 ( 
.A(n_1455),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1506),
.B(n_1377),
.Y(n_1539)
);

NAND3xp33_ASAP7_75t_SL g1540 ( 
.A(n_1512),
.B(n_1334),
.C(n_1420),
.Y(n_1540)
);

OAI221xp5_ASAP7_75t_L g1541 ( 
.A1(n_1500),
.A2(n_1333),
.B1(n_1365),
.B2(n_1381),
.C(n_1389),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1461),
.Y(n_1542)
);

INVx4_ASAP7_75t_L g1543 ( 
.A(n_1511),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1484),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1484),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1485),
.B(n_1377),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1487),
.B(n_1377),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1468),
.B(n_1417),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1477),
.Y(n_1549)
);

NOR3xp33_ASAP7_75t_L g1550 ( 
.A(n_1459),
.B(n_1421),
.C(n_1424),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1488),
.B(n_1384),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1500),
.A2(n_1479),
.B(n_1465),
.Y(n_1552)
);

NOR2x1_ASAP7_75t_L g1553 ( 
.A(n_1486),
.B(n_1416),
.Y(n_1553)
);

OAI211xp5_ASAP7_75t_SL g1554 ( 
.A1(n_1462),
.A2(n_1364),
.B(n_1430),
.C(n_1402),
.Y(n_1554)
);

NOR2x1_ASAP7_75t_L g1555 ( 
.A(n_1486),
.B(n_1416),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1493),
.B(n_1384),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1544),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1518),
.B(n_1470),
.Y(n_1558)
);

NAND3xp33_ASAP7_75t_L g1559 ( 
.A(n_1550),
.B(n_1497),
.C(n_1506),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1539),
.B(n_1497),
.Y(n_1560)
);

AOI221xp5_ASAP7_75t_L g1561 ( 
.A1(n_1540),
.A2(n_1494),
.B1(n_1451),
.B2(n_1452),
.C(n_1508),
.Y(n_1561)
);

NAND4xp25_ASAP7_75t_L g1562 ( 
.A(n_1526),
.B(n_1508),
.C(n_1483),
.D(n_1492),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1527),
.B(n_1458),
.Y(n_1563)
);

AOI221xp5_ASAP7_75t_L g1564 ( 
.A1(n_1529),
.A2(n_1533),
.B1(n_1514),
.B2(n_1517),
.C(n_1520),
.Y(n_1564)
);

NAND3xp33_ASAP7_75t_L g1565 ( 
.A(n_1526),
.B(n_1510),
.C(n_1498),
.Y(n_1565)
);

AOI221xp5_ASAP7_75t_L g1566 ( 
.A1(n_1517),
.A2(n_1520),
.B1(n_1515),
.B2(n_1524),
.C(n_1532),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1537),
.B(n_1495),
.Y(n_1567)
);

NAND3xp33_ASAP7_75t_L g1568 ( 
.A(n_1541),
.B(n_1510),
.C(n_1498),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1537),
.B(n_1495),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1527),
.A2(n_1483),
.B1(n_1511),
.B2(n_1479),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1535),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1544),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1546),
.B(n_1496),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1546),
.B(n_1496),
.Y(n_1574)
);

NAND3xp33_ASAP7_75t_L g1575 ( 
.A(n_1554),
.B(n_1498),
.C(n_1463),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1547),
.B(n_1519),
.Y(n_1576)
);

NAND3xp33_ASAP7_75t_L g1577 ( 
.A(n_1552),
.B(n_1498),
.C(n_1463),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_SL g1578 ( 
.A1(n_1534),
.A2(n_1450),
.B(n_1509),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1528),
.A2(n_1511),
.B1(n_1479),
.B2(n_1450),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1528),
.A2(n_1454),
.B1(n_1479),
.B2(n_1513),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1519),
.B(n_1499),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1531),
.B(n_1459),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1549),
.Y(n_1583)
);

NOR2xp67_ASAP7_75t_L g1584 ( 
.A(n_1538),
.B(n_1469),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1515),
.A2(n_1454),
.B1(n_1513),
.B2(n_1464),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1522),
.B(n_1507),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1521),
.B(n_1523),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1551),
.B(n_1504),
.Y(n_1588)
);

OAI21xp5_ASAP7_75t_SL g1589 ( 
.A1(n_1534),
.A2(n_1502),
.B(n_1503),
.Y(n_1589)
);

OA21x2_ASAP7_75t_L g1590 ( 
.A1(n_1545),
.A2(n_1481),
.B(n_1475),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1531),
.B(n_1469),
.Y(n_1591)
);

NAND3xp33_ASAP7_75t_L g1592 ( 
.A(n_1553),
.B(n_1482),
.C(n_1478),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1551),
.B(n_1501),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1556),
.B(n_1476),
.Y(n_1594)
);

NAND3xp33_ASAP7_75t_L g1595 ( 
.A(n_1553),
.B(n_1482),
.C(n_1489),
.Y(n_1595)
);

NAND3xp33_ASAP7_75t_SL g1596 ( 
.A(n_1516),
.B(n_1420),
.C(n_1334),
.Y(n_1596)
);

NAND3xp33_ASAP7_75t_L g1597 ( 
.A(n_1548),
.B(n_1489),
.C(n_1478),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1530),
.A2(n_1464),
.B1(n_1511),
.B2(n_1491),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1521),
.B(n_1523),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1556),
.B(n_1476),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1563),
.B(n_1587),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1571),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1583),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1557),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1584),
.B(n_1538),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1560),
.B(n_1549),
.Y(n_1606)
);

INVxp67_ASAP7_75t_SL g1607 ( 
.A(n_1557),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1572),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1572),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1581),
.B(n_1536),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1567),
.B(n_1536),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1599),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1569),
.B(n_1536),
.Y(n_1613)
);

OR2x6_ASAP7_75t_L g1614 ( 
.A(n_1584),
.B(n_1455),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1577),
.B(n_1516),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1577),
.B(n_1565),
.Y(n_1616)
);

INVxp67_ASAP7_75t_SL g1617 ( 
.A(n_1592),
.Y(n_1617)
);

INVx1_ASAP7_75t_SL g1618 ( 
.A(n_1591),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1590),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1590),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1590),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1593),
.B(n_1525),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1573),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1588),
.B(n_1536),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1594),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1600),
.B(n_1536),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1576),
.B(n_1525),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1598),
.B(n_1530),
.Y(n_1628)
);

BUFx2_ASAP7_75t_SL g1629 ( 
.A(n_1582),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1574),
.B(n_1542),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1592),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1604),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1623),
.B(n_1566),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1623),
.B(n_1559),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1627),
.B(n_1589),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1627),
.B(n_1530),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1605),
.B(n_1597),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1604),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1604),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1616),
.B(n_1559),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1624),
.B(n_1565),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1627),
.B(n_1530),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1609),
.Y(n_1643)
);

NOR2x1_ASAP7_75t_L g1644 ( 
.A(n_1616),
.B(n_1595),
.Y(n_1644)
);

NAND4xp75_ASAP7_75t_L g1645 ( 
.A(n_1616),
.B(n_1561),
.C(n_1555),
.D(n_1564),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1609),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1609),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1607),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1607),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1624),
.B(n_1558),
.Y(n_1650)
);

INVxp67_ASAP7_75t_SL g1651 ( 
.A(n_1631),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1608),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1608),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1622),
.B(n_1543),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1608),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1626),
.B(n_1610),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1622),
.B(n_1543),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1608),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1626),
.B(n_1548),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1602),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1601),
.Y(n_1661)
);

NAND2xp33_ASAP7_75t_L g1662 ( 
.A(n_1631),
.B(n_1575),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1617),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1623),
.B(n_1575),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1622),
.B(n_1543),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1611),
.B(n_1562),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1606),
.B(n_1630),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1612),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1612),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1640),
.A2(n_1617),
.B(n_1578),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1643),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1643),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1646),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1633),
.B(n_1364),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1634),
.B(n_1618),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1664),
.B(n_1611),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1663),
.B(n_1618),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1651),
.B(n_1641),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1644),
.B(n_1625),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1635),
.B(n_1629),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1662),
.A2(n_1628),
.B1(n_1629),
.B2(n_1568),
.Y(n_1681)
);

INVx2_ASAP7_75t_SL g1682 ( 
.A(n_1637),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1637),
.B(n_1605),
.Y(n_1683)
);

NOR5xp2_ASAP7_75t_L g1684 ( 
.A(n_1648),
.B(n_1603),
.C(n_1595),
.D(n_1568),
.E(n_1621),
.Y(n_1684)
);

INVxp33_ASAP7_75t_SL g1685 ( 
.A(n_1645),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1653),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1637),
.B(n_1635),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1646),
.Y(n_1688)
);

INVxp67_ASAP7_75t_SL g1689 ( 
.A(n_1662),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1636),
.B(n_1629),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1645),
.B(n_1430),
.Y(n_1691)
);

NOR5xp2_ASAP7_75t_L g1692 ( 
.A(n_1648),
.B(n_1603),
.C(n_1621),
.D(n_1620),
.E(n_1612),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1666),
.B(n_1625),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1653),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1666),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1647),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1647),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1660),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1632),
.Y(n_1699)
);

INVx1_ASAP7_75t_SL g1700 ( 
.A(n_1650),
.Y(n_1700)
);

NOR3xp33_ASAP7_75t_L g1701 ( 
.A(n_1641),
.B(n_1596),
.C(n_1615),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1650),
.B(n_1613),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1667),
.B(n_1625),
.Y(n_1703)
);

INVx3_ASAP7_75t_L g1704 ( 
.A(n_1660),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1636),
.B(n_1601),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1649),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1642),
.B(n_1654),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1654),
.B(n_1625),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1657),
.B(n_1606),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1642),
.B(n_1601),
.Y(n_1710)
);

NAND2x1p5_ASAP7_75t_L g1711 ( 
.A(n_1649),
.B(n_1555),
.Y(n_1711)
);

INVxp67_ASAP7_75t_L g1712 ( 
.A(n_1657),
.Y(n_1712)
);

OAI21xp33_ASAP7_75t_L g1713 ( 
.A1(n_1685),
.A2(n_1615),
.B(n_1585),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1695),
.B(n_1656),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1685),
.A2(n_1628),
.B1(n_1665),
.B2(n_1580),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1678),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1704),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1704),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1678),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1671),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1674),
.B(n_1691),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1680),
.B(n_1665),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1706),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1687),
.B(n_1682),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1687),
.B(n_1614),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1704),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1686),
.Y(n_1727)
);

INVxp67_ASAP7_75t_L g1728 ( 
.A(n_1689),
.Y(n_1728)
);

INVx5_ASAP7_75t_SL g1729 ( 
.A(n_1687),
.Y(n_1729)
);

BUFx3_ASAP7_75t_L g1730 ( 
.A(n_1682),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1680),
.B(n_1661),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1700),
.B(n_1656),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1683),
.B(n_1614),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1707),
.B(n_1659),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1686),
.Y(n_1735)
);

NOR2x1_ASAP7_75t_L g1736 ( 
.A(n_1670),
.B(n_1638),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1671),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1694),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1677),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1679),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1672),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1693),
.B(n_1659),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1694),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1701),
.A2(n_1628),
.B1(n_1579),
.B2(n_1570),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1672),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1690),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1675),
.B(n_1676),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1676),
.B(n_1613),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1728),
.B(n_1712),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1728),
.B(n_1705),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1716),
.B(n_1705),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_1724),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1739),
.B(n_1709),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_1730),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1723),
.Y(n_1755)
);

OAI221xp5_ASAP7_75t_L g1756 ( 
.A1(n_1736),
.A2(n_1681),
.B1(n_1711),
.B2(n_1690),
.C(n_1684),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1716),
.B(n_1710),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1719),
.B(n_1710),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1736),
.A2(n_1683),
.B1(n_1711),
.B2(n_1615),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1745),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1729),
.B(n_1707),
.Y(n_1761)
);

OA22x2_ASAP7_75t_L g1762 ( 
.A1(n_1713),
.A2(n_1683),
.B1(n_1699),
.B2(n_1673),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1719),
.B(n_1708),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1739),
.B(n_1703),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1713),
.A2(n_1721),
.B(n_1747),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1747),
.A2(n_1711),
.B(n_1699),
.Y(n_1766)
);

NOR2x1_ASAP7_75t_L g1767 ( 
.A(n_1730),
.B(n_1673),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1745),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1720),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1746),
.A2(n_1729),
.B1(n_1724),
.B2(n_1722),
.Y(n_1770)
);

CKINVDCx20_ASAP7_75t_R g1771 ( 
.A(n_1729),
.Y(n_1771)
);

NOR2x1_ASAP7_75t_L g1772 ( 
.A(n_1730),
.B(n_1688),
.Y(n_1772)
);

OAI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1715),
.A2(n_1696),
.B(n_1688),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1720),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1765),
.B(n_1746),
.Y(n_1775)
);

AND2x4_ASAP7_75t_L g1776 ( 
.A(n_1754),
.B(n_1724),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_SL g1777 ( 
.A(n_1771),
.B(n_1724),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1771),
.B(n_1729),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1755),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1752),
.B(n_1740),
.Y(n_1780)
);

NOR2x1_ASAP7_75t_L g1781 ( 
.A(n_1754),
.B(n_1740),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1755),
.B(n_1722),
.Y(n_1782)
);

AND2x4_ASAP7_75t_SL g1783 ( 
.A(n_1761),
.B(n_1725),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1749),
.B(n_1729),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1770),
.B(n_1731),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1760),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1762),
.B(n_1731),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1753),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1750),
.B(n_1714),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1751),
.B(n_1714),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1762),
.B(n_1734),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1768),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1769),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1773),
.B(n_1734),
.Y(n_1794)
);

NAND2x1_ASAP7_75t_L g1795 ( 
.A(n_1776),
.B(n_1767),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1775),
.A2(n_1756),
.B(n_1759),
.Y(n_1796)
);

AOI21xp5_ASAP7_75t_SL g1797 ( 
.A1(n_1778),
.A2(n_1327),
.B(n_1766),
.Y(n_1797)
);

AOI221x1_ASAP7_75t_L g1798 ( 
.A1(n_1779),
.A2(n_1774),
.B1(n_1757),
.B2(n_1758),
.C(n_1763),
.Y(n_1798)
);

O2A1O1Ixp5_ASAP7_75t_SL g1799 ( 
.A1(n_1786),
.A2(n_1737),
.B(n_1741),
.C(n_1764),
.Y(n_1799)
);

AOI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1794),
.A2(n_1787),
.B1(n_1791),
.B2(n_1788),
.C(n_1780),
.Y(n_1800)
);

O2A1O1Ixp33_ASAP7_75t_SL g1801 ( 
.A1(n_1782),
.A2(n_1732),
.B(n_1772),
.C(n_1737),
.Y(n_1801)
);

NAND4xp25_ASAP7_75t_L g1802 ( 
.A(n_1777),
.B(n_1744),
.C(n_1725),
.D(n_1732),
.Y(n_1802)
);

OAI221xp5_ASAP7_75t_L g1803 ( 
.A1(n_1778),
.A2(n_1744),
.B1(n_1742),
.B2(n_1741),
.C(n_1748),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1784),
.B(n_1438),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1781),
.A2(n_1725),
.B(n_1718),
.Y(n_1805)
);

XNOR2xp5_ASAP7_75t_L g1806 ( 
.A(n_1785),
.B(n_1327),
.Y(n_1806)
);

AOI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1796),
.A2(n_1794),
.B1(n_1785),
.B2(n_1791),
.Y(n_1807)
);

NAND5xp2_ASAP7_75t_L g1808 ( 
.A(n_1800),
.B(n_1787),
.C(n_1789),
.D(n_1790),
.E(n_1792),
.Y(n_1808)
);

NOR2x1_ASAP7_75t_L g1809 ( 
.A(n_1795),
.B(n_1776),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1798),
.B(n_1776),
.Y(n_1810)
);

NAND4xp75_ASAP7_75t_L g1811 ( 
.A(n_1805),
.B(n_1793),
.C(n_1727),
.D(n_1735),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1801),
.Y(n_1812)
);

OA22x2_ASAP7_75t_L g1813 ( 
.A1(n_1806),
.A2(n_1783),
.B1(n_1725),
.B2(n_1733),
.Y(n_1813)
);

NOR3xp33_ASAP7_75t_SL g1814 ( 
.A(n_1802),
.B(n_1783),
.C(n_1586),
.Y(n_1814)
);

NOR2x1_ASAP7_75t_L g1815 ( 
.A(n_1797),
.B(n_1381),
.Y(n_1815)
);

NOR2x1_ASAP7_75t_L g1816 ( 
.A(n_1804),
.B(n_1343),
.Y(n_1816)
);

NOR3xp33_ASAP7_75t_L g1817 ( 
.A(n_1803),
.B(n_1735),
.C(n_1727),
.Y(n_1817)
);

NAND3xp33_ASAP7_75t_SL g1818 ( 
.A(n_1807),
.B(n_1799),
.C(n_1810),
.Y(n_1818)
);

NAND3xp33_ASAP7_75t_SL g1819 ( 
.A(n_1812),
.B(n_1692),
.C(n_1742),
.Y(n_1819)
);

NOR3x1_ASAP7_75t_L g1820 ( 
.A(n_1811),
.B(n_1748),
.C(n_1702),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1808),
.B(n_1727),
.Y(n_1821)
);

NAND4xp25_ASAP7_75t_SL g1822 ( 
.A(n_1815),
.B(n_1717),
.C(n_1718),
.D(n_1726),
.Y(n_1822)
);

NOR2x1_ASAP7_75t_L g1823 ( 
.A(n_1809),
.B(n_1717),
.Y(n_1823)
);

NAND4xp25_ASAP7_75t_L g1824 ( 
.A(n_1816),
.B(n_1733),
.C(n_1738),
.D(n_1735),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1813),
.B(n_1438),
.Y(n_1825)
);

AOI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1818),
.A2(n_1814),
.B1(n_1817),
.B2(n_1733),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1823),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1821),
.Y(n_1828)
);

INVxp67_ASAP7_75t_L g1829 ( 
.A(n_1825),
.Y(n_1829)
);

AOI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1819),
.A2(n_1733),
.B1(n_1738),
.B2(n_1743),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1824),
.Y(n_1831)
);

AOI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1822),
.A2(n_1743),
.B1(n_1738),
.B2(n_1726),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1828),
.B(n_1743),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1827),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1826),
.A2(n_1726),
.B1(n_1718),
.B2(n_1717),
.Y(n_1835)
);

NAND3xp33_ASAP7_75t_L g1836 ( 
.A(n_1831),
.B(n_1820),
.C(n_1697),
.Y(n_1836)
);

OAI211xp5_ASAP7_75t_L g1837 ( 
.A1(n_1830),
.A2(n_1696),
.B(n_1697),
.C(n_1698),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1833),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1834),
.B(n_1829),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1836),
.B(n_1832),
.Y(n_1840)
);

OAI22x1_ASAP7_75t_L g1841 ( 
.A1(n_1839),
.A2(n_1838),
.B1(n_1840),
.B2(n_1835),
.Y(n_1841)
);

NAND4xp75_ASAP7_75t_L g1842 ( 
.A(n_1841),
.B(n_1837),
.C(n_1402),
.D(n_1403),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1842),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1842),
.A2(n_1698),
.B(n_1702),
.Y(n_1844)
);

OA21x2_ASAP7_75t_L g1845 ( 
.A1(n_1843),
.A2(n_1619),
.B(n_1620),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1844),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1846),
.B(n_1403),
.Y(n_1847)
);

AOI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1845),
.A2(n_1403),
.B(n_1652),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1847),
.B(n_1845),
.Y(n_1849)
);

OAI211xp5_ASAP7_75t_L g1850 ( 
.A1(n_1849),
.A2(n_1848),
.B(n_1845),
.C(n_1639),
.Y(n_1850)
);

AOI221xp5_ASAP7_75t_L g1851 ( 
.A1(n_1850),
.A2(n_1652),
.B1(n_1658),
.B2(n_1655),
.C(n_1668),
.Y(n_1851)
);

AOI211xp5_ASAP7_75t_L g1852 ( 
.A1(n_1851),
.A2(n_1669),
.B(n_1668),
.C(n_1605),
.Y(n_1852)
);


endmodule