module fake_ariane_3258_n_97 (n_8, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_10, n_97);

input n_8;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_10;

output n_97;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_74;
wire n_33;
wire n_40;
wire n_53;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_88;
wire n_68;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_35;
wire n_54;
wire n_25;

INVx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

OA21x2_ASAP7_75t_L g28 ( 
.A1(n_4),
.A2(n_19),
.B(n_6),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_11),
.A2(n_4),
.B1(n_16),
.B2(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

OA21x2_ASAP7_75t_L g35 ( 
.A1(n_0),
.A2(n_6),
.B(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

AND2x4_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_5),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_3),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_3),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_7),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_23),
.B(n_7),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_29),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_38),
.B(n_25),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_38),
.B(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

OAI21x1_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_50),
.B(n_44),
.Y(n_55)
);

AOI21x1_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_28),
.B(n_31),
.Y(n_56)
);

AO31x2_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_30),
.A3(n_35),
.B(n_28),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_54),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_41),
.C(n_42),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_35),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_57),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVxp33_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_58),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_63),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_64),
.B1(n_51),
.B2(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_59),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_75),
.A2(n_69),
.B(n_51),
.C(n_67),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_67),
.B(n_68),
.Y(n_78)
);

AOI322xp5_ASAP7_75t_L g79 ( 
.A1(n_74),
.A2(n_40),
.A3(n_36),
.B1(n_32),
.B2(n_23),
.C1(n_35),
.C2(n_34),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_28),
.C(n_32),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_65),
.Y(n_81)
);

AOI221xp5_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_36),
.B1(n_32),
.B2(n_76),
.C(n_34),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_40),
.Y(n_83)
);

NAND4xp75_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_29),
.C(n_23),
.D(n_32),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_36),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_36),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_84),
.Y(n_87)
);

XOR2x1_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_86),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_87),
.Y(n_90)
);

AO22x2_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_88),
.B1(n_61),
.B2(n_36),
.Y(n_91)
);

AOI221xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_24),
.B1(n_34),
.B2(n_23),
.C(n_61),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

AOI22x1_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_24),
.B1(n_34),
.B2(n_61),
.Y(n_94)
);

OA21x2_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_24),
.B(n_34),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_91),
.B1(n_92),
.B2(n_24),
.Y(n_96)
);

OR2x6_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_95),
.Y(n_97)
);


endmodule