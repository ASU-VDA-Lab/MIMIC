module fake_jpeg_3016_n_66 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_66);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_66;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_31;
wire n_25;
wire n_17;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_8),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx8_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_22),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_9),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_16),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_16),
.B1(n_23),
.B2(n_12),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_37),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_15),
.C(n_14),
.Y(n_35)
);

FAx1_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_22),
.CI(n_36),
.CON(n_43),
.SN(n_43)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_18),
.Y(n_36)
);

NOR2xp67_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_22),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_11),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_18),
.Y(n_39)
);

NOR3xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_43),
.C(n_19),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_17),
.B(n_11),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_32),
.B(n_34),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_36),
.B(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_48),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_45),
.B1(n_40),
.B2(n_31),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_33),
.B(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_16),
.B1(n_17),
.B2(n_13),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_51),
.C(n_25),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_55),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_53),
.C(n_54),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_6),
.Y(n_60)
);

AO221x1_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_51),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_SL g59 ( 
.A1(n_58),
.A2(n_43),
.B(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_59),
.B(n_60),
.Y(n_61)
);

AOI322xp5_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_56),
.A3(n_57),
.B1(n_13),
.B2(n_7),
.C1(n_6),
.C2(n_0),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_62),
.A2(n_13),
.B(n_0),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_63),
.A2(n_61),
.B1(n_13),
.B2(n_3),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_0),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_3),
.Y(n_66)
);


endmodule