module fake_jpeg_1015_n_444 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_444);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_444;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g127 ( 
.A(n_51),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_16),
.A2(n_8),
.B1(n_12),
.B2(n_11),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_36),
.B1(n_22),
.B2(n_42),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_8),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_75),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_30),
.B(n_8),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_62),
.B(n_67),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_63),
.A2(n_42),
.B1(n_37),
.B2(n_36),
.Y(n_108)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_17),
.B(n_6),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_17),
.B(n_6),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_69),
.B(n_76),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_21),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_70),
.B(n_81),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_71),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_73),
.B(n_74),
.Y(n_118)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_23),
.B(n_4),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_23),
.B(n_27),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_84),
.Y(n_97)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_80),
.B(n_86),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_21),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_25),
.B(n_13),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_25),
.Y(n_109)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

INVx2_ASAP7_75t_R g131 ( 
.A(n_83),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_21),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_27),
.B(n_4),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_25),
.Y(n_106)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g154 ( 
.A1(n_87),
.A2(n_117),
.B(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_20),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_88),
.B(n_114),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_40),
.C(n_39),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_102),
.B(n_31),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_106),
.B(n_115),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_108),
.A2(n_121),
.B1(n_29),
.B2(n_38),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_113),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_51),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_22),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_41),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_41),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_37),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_120),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_37),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_47),
.A2(n_31),
.B1(n_38),
.B2(n_40),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_46),
.B(n_34),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_55),
.B(n_34),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_86),
.A2(n_15),
.B1(n_32),
.B2(n_28),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_134),
.B1(n_43),
.B2(n_32),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_70),
.B(n_15),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_126),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_48),
.A2(n_15),
.B1(n_32),
.B2(n_28),
.Y(n_134)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_136),
.Y(n_193)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_81),
.B1(n_54),
.B2(n_28),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_127),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_141),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_43),
.B1(n_83),
.B2(n_40),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_143),
.A2(n_156),
.B1(n_166),
.B2(n_168),
.Y(n_181)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_147),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_88),
.A2(n_63),
.B(n_43),
.C(n_72),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_157),
.B(n_111),
.C(n_135),
.Y(n_187)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_150),
.Y(n_214)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_102),
.B1(n_129),
.B2(n_93),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_152),
.A2(n_160),
.B1(n_163),
.B2(n_169),
.Y(n_213)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_97),
.A2(n_61),
.B1(n_45),
.B2(n_50),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_91),
.B(n_89),
.C(n_93),
.D(n_100),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_133),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_172),
.Y(n_186)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_100),
.A2(n_52),
.B1(n_71),
.B2(n_68),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_161),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_164),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_109),
.A2(n_65),
.B1(n_59),
.B2(n_56),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_101),
.B(n_0),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_0),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_165),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_116),
.A2(n_128),
.B1(n_127),
.B2(n_104),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_99),
.Y(n_167)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_116),
.A2(n_79),
.B1(n_64),
.B2(n_21),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_95),
.A2(n_53),
.B1(n_38),
.B2(n_18),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_128),
.A2(n_18),
.B1(n_44),
.B2(n_29),
.Y(n_170)
);

INVx11_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_101),
.B(n_0),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_171),
.B(n_175),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_133),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_126),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_111),
.B(n_0),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_131),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_177),
.A2(n_103),
.B1(n_131),
.B2(n_105),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_127),
.A2(n_29),
.B1(n_9),
.B2(n_3),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_178),
.A2(n_103),
.B1(n_104),
.B2(n_131),
.Y(n_182)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_92),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_179),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_95),
.A2(n_29),
.B1(n_2),
.B2(n_1),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_130),
.B1(n_96),
.B2(n_1),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_182),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_185),
.A2(n_191),
.B1(n_202),
.B2(n_207),
.Y(n_228)
);

A2O1A1O1Ixp25_ASAP7_75t_L g254 ( 
.A1(n_187),
.A2(n_212),
.B(n_186),
.C(n_188),
.D(n_190),
.Y(n_254)
);

O2A1O1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_135),
.B(n_90),
.C(n_124),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_190),
.A2(n_206),
.B(n_184),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_137),
.A2(n_105),
.B1(n_107),
.B2(n_92),
.Y(n_191)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_145),
.B(n_135),
.CI(n_94),
.CON(n_196),
.SN(n_196)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_196),
.B(n_201),
.Y(n_238)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_145),
.A2(n_140),
.A3(n_146),
.B1(n_155),
.B2(n_162),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_157),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_142),
.B(n_110),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_177),
.A2(n_92),
.B1(n_107),
.B2(n_132),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_155),
.B(n_124),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_204),
.B(n_210),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_147),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_139),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_172),
.A2(n_135),
.B(n_90),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_142),
.A2(n_107),
.B1(n_132),
.B2(n_130),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_209),
.A2(n_141),
.B1(n_176),
.B2(n_180),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_173),
.B(n_12),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_140),
.B(n_96),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_212),
.C(n_158),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_152),
.B(n_112),
.C(n_4),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_162),
.B(n_112),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_218),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_149),
.B(n_112),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_222),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_214),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_234),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_224),
.B(n_227),
.Y(n_289)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_225),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_149),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_226),
.Y(n_290)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_229),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_163),
.B1(n_148),
.B2(n_154),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_230),
.A2(n_213),
.B1(n_208),
.B2(n_184),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_183),
.A2(n_192),
.B1(n_194),
.B2(n_201),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_258),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_186),
.A2(n_161),
.B(n_165),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_232),
.A2(n_254),
.B(n_259),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_144),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_233),
.B(n_237),
.Y(n_269)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_235),
.B(n_242),
.Y(n_277)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_236),
.B(n_239),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_144),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_164),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_240),
.B(n_248),
.C(n_252),
.Y(n_292)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_193),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_243),
.B(n_247),
.Y(n_278)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_244),
.B(n_246),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_171),
.C(n_175),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_193),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_250),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_183),
.B(n_150),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_188),
.B(n_165),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_192),
.B(n_160),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_217),
.Y(n_283)
);

BUFx12_ASAP7_75t_L g255 ( 
.A(n_205),
.Y(n_255)
);

INVx13_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_220),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_256),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_219),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_257),
.B(n_190),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_184),
.A2(n_179),
.B1(n_167),
.B2(n_159),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_221),
.A2(n_147),
.B(n_153),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_197),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_270),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_263),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_187),
.B(n_221),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_264),
.A2(n_266),
.B(n_136),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_189),
.B(n_181),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_232),
.B(n_203),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_268),
.B(n_251),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_197),
.Y(n_270)
);

INVx13_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_271),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_272),
.A2(n_202),
.B1(n_258),
.B2(n_207),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_196),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_273),
.B(n_276),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_230),
.A2(n_228),
.B1(n_227),
.B2(n_224),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_275),
.A2(n_292),
.B1(n_288),
.B2(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_241),
.B(n_196),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_224),
.B(n_216),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_288),
.C(n_268),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_283),
.B(n_191),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_241),
.B(n_216),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_286),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_222),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_285),
.B(n_243),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_238),
.B(n_210),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_238),
.B(n_200),
.Y(n_287)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_287),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_185),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_269),
.B(n_251),
.Y(n_295)
);

NAND3xp33_ASAP7_75t_L g346 ( 
.A(n_295),
.B(n_265),
.C(n_279),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_322),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_261),
.A2(n_245),
.B1(n_254),
.B2(n_208),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_300),
.B(n_313),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_260),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_324),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_228),
.B1(n_245),
.B2(n_208),
.Y(n_302)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_302),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_244),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_304),
.B(n_307),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_262),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_305),
.B(n_286),
.Y(n_332)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_294),
.Y(n_306)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_306),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_236),
.C(n_229),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_309),
.C(n_314),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_235),
.C(n_259),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_311),
.A2(n_316),
.B1(n_318),
.B2(n_263),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_198),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_294),
.Y(n_315)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_315),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_293),
.A2(n_209),
.B1(n_223),
.B2(n_200),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_293),
.A2(n_222),
.B1(n_249),
.B2(n_242),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_275),
.A2(n_293),
.B1(n_261),
.B2(n_274),
.Y(n_319)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_278),
.A2(n_234),
.B1(n_198),
.B2(n_255),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_280),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_274),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_321),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_323),
.A2(n_266),
.B(n_278),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_260),
.Y(n_324)
);

O2A1O1Ixp33_ASAP7_75t_L g326 ( 
.A1(n_298),
.A2(n_264),
.B(n_276),
.C(n_273),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_326),
.A2(n_335),
.B(n_336),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_331),
.A2(n_311),
.B1(n_310),
.B2(n_309),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_332),
.A2(n_346),
.B1(n_285),
.B2(n_267),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_333),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_323),
.A2(n_280),
.B(n_281),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_282),
.C(n_270),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_339),
.C(n_307),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_283),
.C(n_281),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_312),
.A2(n_287),
.B1(n_280),
.B2(n_284),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_341),
.A2(n_347),
.B1(n_277),
.B2(n_303),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_322),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_345),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_299),
.B(n_265),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_312),
.A2(n_298),
.B1(n_317),
.B2(n_316),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_320),
.Y(n_348)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_348),
.Y(n_369)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_306),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_350),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_299),
.B(n_279),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_351),
.B(n_317),
.Y(n_352)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_354),
.B(n_357),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_355),
.A2(n_342),
.B1(n_327),
.B2(n_325),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_340),
.B(n_314),
.C(n_313),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_368),
.C(n_373),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_328),
.B(n_300),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_310),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_358),
.B(n_360),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_303),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_359),
.B(n_333),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_328),
.B(n_318),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_277),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_361),
.B(n_365),
.Y(n_383)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_363),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_349),
.B(n_322),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_271),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_366),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_271),
.Y(n_368)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_370),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_326),
.B(n_267),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_371),
.B(n_372),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_327),
.A2(n_291),
.B1(n_267),
.B2(n_255),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_330),
.B(n_291),
.C(n_219),
.Y(n_373)
);

OAI21x1_ASAP7_75t_SL g381 ( 
.A1(n_364),
.A2(n_337),
.B(n_336),
.Y(n_381)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_381),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_360),
.B(n_330),
.C(n_342),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_387),
.C(n_390),
.Y(n_400)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_384),
.Y(n_404)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_362),
.Y(n_385)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_385),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_386),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_366),
.B(n_333),
.C(n_348),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_362),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_389),
.B(n_334),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_361),
.B(n_344),
.C(n_325),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g391 ( 
.A(n_353),
.B(n_341),
.CI(n_331),
.CON(n_391),
.SN(n_391)
);

BUFx24_ASAP7_75t_SL g392 ( 
.A(n_391),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_376),
.A2(n_353),
.B(n_367),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_395),
.A2(n_396),
.B(n_391),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_375),
.A2(n_371),
.B(n_367),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_388),
.B(n_358),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_379),
.Y(n_410)
);

AO221x1_ASAP7_75t_L g398 ( 
.A1(n_374),
.A2(n_347),
.B1(n_373),
.B2(n_357),
.C(n_369),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_398),
.B(n_405),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_382),
.A2(n_335),
.B1(n_329),
.B2(n_350),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_401),
.A2(n_403),
.B1(n_387),
.B2(n_379),
.Y(n_408)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_402),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_390),
.Y(n_403)
);

AOI322xp5_ASAP7_75t_SL g405 ( 
.A1(n_383),
.A2(n_354),
.A3(n_365),
.B1(n_334),
.B2(n_356),
.C1(n_368),
.C2(n_329),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_394),
.A2(n_380),
.B1(n_391),
.B2(n_378),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_406),
.B(n_409),
.Y(n_419)
);

AOI21xp33_ASAP7_75t_L g420 ( 
.A1(n_408),
.A2(n_412),
.B(n_393),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_400),
.B(n_377),
.C(n_388),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_410),
.B(n_411),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_SL g411 ( 
.A(n_400),
.B(n_377),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_SL g413 ( 
.A(n_392),
.B(n_383),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_414),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_397),
.B(n_219),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_395),
.B(n_151),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_415),
.B(n_416),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_404),
.B(n_179),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_153),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_399),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_420),
.A2(n_422),
.B(n_428),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_407),
.A2(n_393),
.B(n_399),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_417),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_418),
.B(n_4),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_427),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_10),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_415),
.A2(n_13),
.B(n_10),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_419),
.B(n_421),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_429),
.A2(n_432),
.B(n_426),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_430),
.B(n_431),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_425),
.B(n_410),
.C(n_414),
.Y(n_431)
);

AOI31xp67_ASAP7_75t_L g432 ( 
.A1(n_425),
.A2(n_12),
.A3(n_13),
.B(n_1),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_426),
.A2(n_2),
.B1(n_408),
.B2(n_407),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_434),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_437),
.B(n_438),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_429),
.B(n_428),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_439),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_440),
.B(n_433),
.C(n_436),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_442),
.B(n_441),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_443),
.B(n_435),
.Y(n_444)
);


endmodule