module fake_jpeg_29553_n_439 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_439);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_439;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_332;
wire n_92;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_54),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_23),
.B(n_9),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_21),
.Y(n_101)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_71),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_22),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_78),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_39),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g104 ( 
.A(n_75),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_25),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_79),
.B(n_86),
.Y(n_136)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_31),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_83),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_25),
.Y(n_82)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_85),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_23),
.B(n_9),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_28),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_51),
.B(n_36),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_93),
.B(n_101),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_28),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_105),
.B(n_129),
.Y(n_148)
);

FAx1_ASAP7_75t_SL g152 ( 
.A(n_107),
.B(n_124),
.CI(n_132),
.CON(n_152),
.SN(n_152)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_28),
.B(n_41),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_110),
.C(n_69),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_72),
.A2(n_25),
.B(n_1),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_61),
.B(n_38),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_135),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_82),
.A2(n_21),
.B1(n_44),
.B2(n_40),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_122),
.A2(n_123),
.B1(n_104),
.B2(n_68),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_86),
.A2(n_40),
.B1(n_39),
.B2(n_30),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_67),
.B(n_36),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_70),
.B(n_41),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_76),
.B(n_38),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_30),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_84),
.B1(n_59),
.B2(n_58),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_139),
.B(n_142),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_140),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_141),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_122),
.A2(n_47),
.B1(n_49),
.B2(n_55),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_39),
.B1(n_40),
.B2(n_71),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_145),
.Y(n_179)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

AO22x1_ASAP7_75t_SL g145 ( 
.A1(n_89),
.A2(n_64),
.B1(n_77),
.B2(n_56),
.Y(n_145)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_102),
.A2(n_48),
.B1(n_57),
.B2(n_65),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_157),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_155),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_29),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_154),
.B(n_156),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_97),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_29),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_107),
.A2(n_35),
.B1(n_12),
.B2(n_3),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_90),
.B(n_29),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_161),
.Y(n_186)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_100),
.B(n_94),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_104),
.A2(n_137),
.B1(n_115),
.B2(n_119),
.Y(n_163)
);

NAND2xp33_ASAP7_75t_SL g185 ( 
.A(n_163),
.B(n_166),
.Y(n_185)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

CKINVDCx9p33_ASAP7_75t_R g166 ( 
.A(n_108),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

BUFx16f_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_118),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_171),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_29),
.Y(n_171)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_173),
.Y(n_183)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_125),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_201),
.C(n_180),
.Y(n_210)
);

FAx1_ASAP7_75t_SL g180 ( 
.A(n_148),
.B(n_103),
.CI(n_117),
.CON(n_180),
.SN(n_180)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_180),
.B(n_145),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_98),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_188),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_98),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_117),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_157),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_152),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_202),
.B(n_169),
.Y(n_246)
);

INVx4_ASAP7_75t_SL g203 ( 
.A(n_187),
.Y(n_203)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_211),
.Y(n_238)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_143),
.B(n_150),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_185),
.B(n_177),
.Y(n_231)
);

AOI32xp33_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_151),
.A3(n_167),
.B1(n_155),
.B2(n_142),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_206),
.A2(n_208),
.B(n_190),
.Y(n_228)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_196),
.A2(n_188),
.B(n_184),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_215),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_165),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_192),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_214),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_213),
.B(n_177),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_158),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_139),
.B1(n_149),
.B2(n_145),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_216),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_176),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_220),
.Y(n_239)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_138),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_194),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_181),
.A2(n_144),
.B1(n_146),
.B2(n_173),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_223),
.A2(n_175),
.B1(n_198),
.B2(n_193),
.Y(n_227)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_174),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_224),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_227),
.A2(n_229),
.B1(n_232),
.B2(n_241),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_228),
.B(n_246),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_179),
.B1(n_182),
.B2(n_197),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_230),
.A2(n_202),
.B1(n_213),
.B2(n_215),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_SL g265 ( 
.A(n_231),
.B(n_236),
.C(n_218),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_212),
.A2(n_222),
.B1(n_214),
.B2(n_205),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_175),
.B(n_199),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_233),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_242),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_208),
.A2(n_106),
.B(n_164),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_205),
.A2(n_140),
.B1(n_141),
.B2(n_130),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_141),
.B1(n_140),
.B2(n_130),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_244),
.A2(n_203),
.B1(n_200),
.B2(n_207),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_210),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_271),
.C(n_246),
.Y(n_279)
);

INVx13_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_251),
.Y(n_297)
);

AND2x6_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_206),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_259),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

INVx5_ASAP7_75t_SL g258 ( 
.A(n_238),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_258),
.Y(n_290)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_238),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_261),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_263),
.A2(n_233),
.B1(n_246),
.B2(n_227),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_235),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_264),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_265),
.A2(n_269),
.B(n_246),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_266),
.A2(n_200),
.B1(n_189),
.B2(n_137),
.Y(n_300)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_267),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_209),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_268),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_229),
.A2(n_202),
.B1(n_224),
.B2(n_209),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_221),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_270),
.B(n_272),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_226),
.B(n_220),
.C(n_195),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_203),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_236),
.B(n_219),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_261),
.Y(n_283)
);

AO22x1_ASAP7_75t_L g275 ( 
.A1(n_265),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_275)
);

O2A1O1Ixp33_ASAP7_75t_L g325 ( 
.A1(n_275),
.A2(n_266),
.B(n_166),
.C(n_168),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_294),
.C(n_299),
.Y(n_303)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_258),
.A2(n_243),
.B1(n_247),
.B2(n_207),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_284),
.A2(n_272),
.B(n_255),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_292),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_260),
.A2(n_227),
.B1(n_241),
.B2(n_225),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_287),
.B(n_250),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_249),
.B(n_233),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_289),
.B(n_262),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_269),
.A2(n_225),
.B1(n_244),
.B2(n_247),
.Y(n_291)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_291),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_248),
.B(n_168),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_195),
.C(n_193),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_160),
.Y(n_298)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_248),
.B(n_99),
.C(n_106),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_300),
.A2(n_257),
.B1(n_256),
.B2(n_204),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_267),
.Y(n_304)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_304),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_306),
.B(n_304),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_264),
.Y(n_308)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_308),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_309),
.A2(n_319),
.B1(n_189),
.B2(n_134),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_275),
.A2(n_250),
.B1(n_256),
.B2(n_252),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_310),
.A2(n_302),
.B1(n_314),
.B2(n_325),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_279),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_311),
.B(n_287),
.Y(n_331)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_313),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_274),
.B(n_263),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_317),
.Y(n_327)
);

AOI21xp33_ASAP7_75t_L g316 ( 
.A1(n_281),
.A2(n_262),
.B(n_251),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_316),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_259),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_294),
.C(n_299),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_291),
.C(n_276),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_275),
.A2(n_285),
.B1(n_282),
.B2(n_290),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_297),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_320),
.Y(n_346)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_280),
.Y(n_321)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_321),
.Y(n_334)
);

XNOR2x1_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_297),
.Y(n_343)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_280),
.Y(n_323)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_324),
.B(n_147),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_326),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_290),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_342),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_320),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_333),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_335),
.B(n_337),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_276),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_336),
.B(n_343),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_303),
.B(n_278),
.C(n_293),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_306),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_338),
.B(n_340),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_303),
.B(n_278),
.C(n_293),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_307),
.B(n_300),
.Y(n_342)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_344),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_331),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_348),
.A2(n_312),
.B1(n_307),
.B2(n_204),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_349),
.A2(n_309),
.B1(n_305),
.B2(n_310),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_318),
.B(n_170),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_350),
.B(n_324),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_330),
.A2(n_314),
.B(n_319),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_352),
.B(n_362),
.Y(n_376)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_334),
.Y(n_353)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_353),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_354),
.B(n_127),
.Y(n_385)
);

A2O1A1Ixp33_ASAP7_75t_L g357 ( 
.A1(n_339),
.A2(n_308),
.B(n_301),
.C(n_321),
.Y(n_357)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_357),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_361),
.Y(n_375)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_332),
.Y(n_359)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_359),
.Y(n_386)
);

AOI322xp5_ASAP7_75t_L g362 ( 
.A1(n_341),
.A2(n_328),
.A3(n_329),
.B1(n_343),
.B2(n_327),
.C1(n_345),
.C2(n_338),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_346),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_365),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_364),
.B(n_346),
.Y(n_377)
);

BUFx24_ASAP7_75t_SL g365 ( 
.A(n_336),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_337),
.B(n_204),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_367),
.B(n_368),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_17),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_342),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_370),
.B(n_371),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_369),
.B(n_335),
.C(n_347),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_95),
.C(n_92),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_377),
.B(n_380),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_351),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_379),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_19),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_134),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_371),
.Y(n_384)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_384),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_385),
.A2(n_364),
.B1(n_357),
.B2(n_172),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_355),
.B(n_15),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_387),
.B(n_13),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_360),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_388),
.B(n_393),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_352),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_400),
.Y(n_409)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_391),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_383),
.B(n_366),
.C(n_358),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_354),
.C(n_360),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_397),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_396),
.A2(n_382),
.B1(n_372),
.B2(n_386),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_375),
.B(n_111),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_380),
.B(n_113),
.C(n_111),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_398),
.B(n_399),
.C(n_400),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_377),
.B(n_113),
.C(n_92),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_389),
.B(n_381),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_402),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_384),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_405),
.B(n_411),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_392),
.A2(n_385),
.B(n_96),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_406),
.B(n_29),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_409),
.B(n_410),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_394),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_394),
.B(n_12),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_389),
.A2(n_95),
.B(n_12),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_412),
.A2(n_10),
.B(n_16),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_408),
.B(n_96),
.C(n_11),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_418),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_404),
.Y(n_414)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_414),
.Y(n_425)
);

MAJx2_ASAP7_75t_L g416 ( 
.A(n_409),
.B(n_11),
.C(n_15),
.Y(n_416)
);

OAI21x1_ASAP7_75t_L g424 ( 
.A1(n_416),
.A2(n_417),
.B(n_406),
.Y(n_424)
);

AOI322xp5_ASAP7_75t_L g418 ( 
.A1(n_410),
.A2(n_69),
.A3(n_68),
.B1(n_61),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_8),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_419),
.B(n_421),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_424),
.B(n_426),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_422),
.A2(n_403),
.B(n_8),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_415),
.B(n_7),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_428),
.A2(n_10),
.B1(n_16),
.B2(n_4),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_422),
.B(n_6),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_429),
.A2(n_420),
.B1(n_35),
.B2(n_3),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_430),
.B(n_5),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_431),
.A2(n_432),
.B(n_13),
.Y(n_435)
);

AOI321xp33_ASAP7_75t_L g432 ( 
.A1(n_425),
.A2(n_423),
.A3(n_427),
.B1(n_5),
.B2(n_11),
.C(n_13),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_434),
.B(n_435),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_436),
.A2(n_433),
.B1(n_35),
.B2(n_1),
.Y(n_437)
);

FAx1_ASAP7_75t_SL g438 ( 
.A(n_437),
.B(n_0),
.CI(n_1),
.CON(n_438),
.SN(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_0),
.B(n_1),
.Y(n_439)
);


endmodule