module real_jpeg_15043_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_3),
.A2(n_66),
.B1(n_69),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_3),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_3),
.A2(n_52),
.B1(n_54),
.B2(n_81),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_81),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_3),
.A2(n_28),
.B1(n_32),
.B2(n_81),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_4),
.A2(n_28),
.B1(n_32),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_43),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_4),
.A2(n_43),
.B1(n_52),
.B2(n_54),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_4),
.A2(n_43),
.B1(n_66),
.B2(n_69),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_5),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_5),
.A2(n_32),
.B(n_35),
.C(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_5),
.B(n_41),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_5),
.A2(n_31),
.B1(n_52),
.B2(n_54),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_5),
.A2(n_90),
.B1(n_119),
.B2(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_5),
.B(n_56),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_10),
.A2(n_28),
.B1(n_32),
.B2(n_47),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_10),
.A2(n_47),
.B1(n_52),
.B2(n_54),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_10),
.A2(n_47),
.B1(n_66),
.B2(n_69),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_11),
.A2(n_66),
.B1(n_69),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_11),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_11),
.A2(n_52),
.B1(n_54),
.B2(n_83),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_83),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_11),
.A2(n_28),
.B1(n_32),
.B2(n_83),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_12),
.A2(n_52),
.B1(n_54),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_12),
.A2(n_66),
.B1(n_69),
.B2(n_74),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_74),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_12),
.A2(n_28),
.B1(n_32),
.B2(n_74),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_13),
.A2(n_52),
.B1(n_54),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_13),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_71),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_13),
.A2(n_66),
.B1(n_69),
.B2(n_71),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_13),
.A2(n_28),
.B1(n_32),
.B2(n_71),
.Y(n_249)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_15),
.A2(n_52),
.B1(n_54),
.B2(n_58),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_15),
.A2(n_58),
.B1(n_66),
.B2(n_69),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_15),
.A2(n_28),
.B1(n_32),
.B2(n_58),
.Y(n_224)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_320),
.C(n_324),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_318),
.B(n_322),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_310),
.B(n_317),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_276),
.B(n_307),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_254),
.B(n_275),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_227),
.B(n_253),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_128),
.B(n_206),
.C(n_226),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_101),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_24),
.B(n_101),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_75),
.C(n_88),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_25),
.B(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_44),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_26),
.B(n_45),
.C(n_59),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_26)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_31),
.A2(n_36),
.B(n_38),
.Y(n_85)
);

HAxp5_ASAP7_75t_SL g138 ( 
.A(n_31),
.B(n_39),
.CON(n_138),
.SN(n_138)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_31),
.B(n_63),
.C(n_69),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_31),
.B(n_90),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_31),
.B(n_65),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_33),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_33),
.A2(n_41),
.B1(n_110),
.B2(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_33),
.B(n_272),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_33),
.A2(n_41),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_33),
.A2(n_41),
.B(n_249),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_37),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_37),
.A2(n_289),
.B(n_290),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_39),
.B1(n_50),
.B2(n_51),
.Y(n_55)
);

NOR3xp33_ASAP7_75t_L g139 ( 
.A(n_38),
.B(n_51),
.C(n_52),
.Y(n_139)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_41),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_41),
.B(n_272),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_59),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B1(n_56),
.B2(n_57),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_46),
.Y(n_100)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_48),
.A2(n_56),
.B1(n_98),
.B2(n_138),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_48),
.A2(n_114),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_48),
.B(n_245),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_48),
.A2(n_56),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_48),
.A2(n_56),
.B(n_114),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_49),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_49),
.B(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_49),
.A2(n_243),
.B(n_244),
.Y(n_242)
);

OA22x2_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_SL g136 ( 
.A1(n_50),
.A2(n_54),
.B(n_137),
.C(n_139),
.Y(n_136)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_52),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_54),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_54),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_56),
.B(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_57),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_70),
.B(n_72),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_60),
.B(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_60),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_60),
.A2(n_145),
.B1(n_147),
.B2(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_60),
.A2(n_147),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_60),
.A2(n_147),
.B1(n_155),
.B2(n_165),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_60),
.A2(n_147),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_60),
.A2(n_72),
.B(n_215),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_60),
.A2(n_70),
.B(n_147),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_63),
.B1(n_66),
.B2(n_69),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_65),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

CKINVDCx6p67_ASAP7_75t_R g69 ( 
.A(n_66),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_69),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_70),
.B(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_75),
.B(n_88),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_82),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_77),
.A2(n_122),
.B(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_77),
.A2(n_78),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_78),
.B(n_141),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_82),
.Y(n_120)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_86),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.C(n_96),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_89),
.A2(n_94),
.B1(n_95),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_93),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_90),
.A2(n_119),
.B1(n_170),
.B2(n_178),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_90),
.A2(n_119),
.B(n_234),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_91),
.B(n_188),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_96),
.B(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g283 ( 
.A1(n_99),
.A2(n_284),
.B(n_285),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_116),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_102),
.B(n_117),
.C(n_127),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_115),
.Y(n_102)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_111),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_106),
.B(n_111),
.C(n_115),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_107),
.A2(n_247),
.B(n_248),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_107),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_107),
.A2(n_271),
.B(n_314),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_113),
.B(n_244),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_127),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_123),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_118),
.B(n_123),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B(n_121),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_119),
.A2(n_172),
.B(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_124),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_125),
.B(n_146),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_201),
.B(n_205),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_156),
.B(n_200),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_151),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_133),
.B(n_151),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_148),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_142),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_135),
.B(n_142),
.C(n_148),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_136),
.B(n_140),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_141),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B(n_146),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.C(n_154),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_154),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_195),
.B(n_199),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_184),
.B(n_194),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_173),
.B(n_183),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_168),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_168),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_163),
.B1(n_166),
.B2(n_167),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_161),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_166),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_179),
.B(n_182),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_181),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_186),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_190),
.C(n_193),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_192),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_198),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_204),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_225),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_225),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_210),
.C(n_217),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_217),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_216),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_216),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_213),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_220),
.C(n_223),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_221),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_224),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_229),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_252),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_237),
.B1(n_250),
.B2(n_251),
.Y(n_230)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_251),
.C(n_252),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_232),
.A2(n_233),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_235),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g292 ( 
.A1(n_233),
.A2(n_266),
.B(n_268),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_242),
.C(n_246),
.Y(n_257)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_243),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_248),
.B(n_290),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_249),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_274),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_274),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_273),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_256),
.B(n_259),
.C(n_265),
.Y(n_305)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_265),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_263),
.B(n_264),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_260),
.B(n_263),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_262),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_279),
.C(n_292),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g306 ( 
.A(n_264),
.B(n_279),
.CI(n_292),
.CON(n_306),
.SN(n_306)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_304),
.Y(n_276)
);

AOI21xp33_ASAP7_75t_L g307 ( 
.A1(n_277),
.A2(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_293),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_278),
.B(n_293),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_288),
.B2(n_291),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_286),
.B2(n_287),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_287),
.C(n_288),
.Y(n_294)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_287),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_297),
.C(n_302),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_288),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_291),
.B1(n_296),
.B2(n_303),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_294),
.C(n_303),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_289),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_296),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_299),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_301),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_306),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_306),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_316),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_316),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_311),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_320),
.Y(n_323)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_313),
.CI(n_315),
.CON(n_311),
.SN(n_311)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_321),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);


endmodule