module fake_jpeg_1705_n_619 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_619);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_619;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_539;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx2_ASAP7_75t_R g58 ( 
.A(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_58),
.B(n_60),
.Y(n_134)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_51),
.Y(n_59)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_21),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_61),
.B(n_62),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_54),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_63),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_64),
.Y(n_135)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_66),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_22),
.B(n_11),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_69),
.B(n_78),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_71),
.B(n_74),
.Y(n_184)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_43),
.B(n_11),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_22),
.B(n_11),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_79),
.B(n_83),
.Y(n_196)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_81),
.Y(n_155)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_40),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_84),
.Y(n_163)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_34),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_86),
.B(n_92),
.Y(n_214)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_87),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_88),
.Y(n_171)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_89),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_90),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_91),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_17),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_94),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_18),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_99),
.B(n_102),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_40),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_24),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_104),
.B(n_108),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_48),
.Y(n_105)
);

CKINVDCx6p67_ASAP7_75t_R g140 ( 
.A(n_105),
.Y(n_140)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_106),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_15),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_48),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_26),
.Y(n_113)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_34),
.Y(n_114)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_34),
.Y(n_115)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_115),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_37),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_34),
.Y(n_117)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_117),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_56),
.B(n_15),
.Y(n_118)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_23),
.Y(n_122)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_122),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_19),
.Y(n_123)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_123),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_27),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_124),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_23),
.Y(n_125)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_125),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_19),
.Y(n_126)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_126),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_19),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_127),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_58),
.B(n_28),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_129),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_28),
.C(n_30),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_131),
.B(n_205),
.Y(n_230)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_136),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_111),
.A2(n_27),
.B1(n_25),
.B2(n_29),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_152),
.A2(n_158),
.B1(n_194),
.B2(n_50),
.Y(n_248)
);

CKINVDCx10_ASAP7_75t_R g157 ( 
.A(n_68),
.Y(n_157)
);

INVx4_ASAP7_75t_SL g293 ( 
.A(n_157),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_67),
.A2(n_27),
.B1(n_25),
.B2(n_29),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_80),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_164),
.B(n_188),
.Y(n_289)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_77),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_174),
.Y(n_292)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_63),
.Y(n_177)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_65),
.Y(n_179)
);

INVx11_ASAP7_75t_L g288 ( 
.A(n_179),
.Y(n_288)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_93),
.Y(n_183)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_183),
.Y(n_286)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_187),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_81),
.Y(n_188)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_70),
.A2(n_25),
.B1(n_50),
.B2(n_36),
.Y(n_194)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_86),
.Y(n_199)
);

INVx3_ASAP7_75t_SL g252 ( 
.A(n_199),
.Y(n_252)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_120),
.Y(n_202)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_202),
.Y(n_260)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_203),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_87),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_73),
.Y(n_206)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_96),
.Y(n_207)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_59),
.Y(n_210)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_210),
.Y(n_255)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_94),
.Y(n_211)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_64),
.B(n_30),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_215),
.Y(n_222)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_66),
.Y(n_213)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_109),
.B(n_47),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_106),
.Y(n_217)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_217),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_114),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_127),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_134),
.A2(n_91),
.B1(n_95),
.B2(n_42),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_220),
.A2(n_234),
.B1(n_251),
.B2(n_207),
.Y(n_307)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_176),
.Y(n_224)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_224),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_216),
.A2(n_155),
.B1(n_151),
.B2(n_208),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_225),
.A2(n_246),
.B1(n_264),
.B2(n_181),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_143),
.B(n_42),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_226),
.B(n_227),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_132),
.B(n_38),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_196),
.Y(n_228)
);

NAND3xp33_ASAP7_75t_L g325 ( 
.A(n_228),
.B(n_229),
.C(n_233),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_134),
.B(n_47),
.Y(n_229)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_147),
.Y(n_231)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_231),
.Y(n_308)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_204),
.Y(n_232)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_232),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_196),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_165),
.A2(n_45),
.B1(n_39),
.B2(n_38),
.Y(n_234)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_138),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_236),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_138),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_237),
.Y(n_341)
);

BUFx4f_ASAP7_75t_L g238 ( 
.A(n_150),
.Y(n_238)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_238),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_135),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_240),
.B(n_249),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_160),
.A2(n_75),
.B1(n_107),
.B2(n_88),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_241),
.A2(n_253),
.B1(n_275),
.B2(n_169),
.Y(n_297)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_146),
.Y(n_242)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_242),
.Y(n_335)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_179),
.Y(n_245)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_245),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_L g246 ( 
.A1(n_152),
.A2(n_84),
.B1(n_90),
.B2(n_100),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_248),
.B(n_195),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_135),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_128),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_250),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_140),
.A2(n_33),
.B1(n_39),
.B2(n_45),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_158),
.A2(n_110),
.B1(n_119),
.B2(n_115),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_184),
.B(n_33),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_254),
.B(n_257),
.Y(n_315)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_200),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_256),
.Y(n_332)
);

NAND3xp33_ASAP7_75t_L g257 ( 
.A(n_212),
.B(n_41),
.C(n_36),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_184),
.B(n_41),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_258),
.B(n_265),
.Y(n_317)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_159),
.Y(n_262)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_262),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_263),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_151),
.A2(n_126),
.B1(n_52),
.B2(n_49),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_182),
.B(n_153),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_175),
.Y(n_266)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_167),
.B(n_12),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_267),
.B(n_271),
.Y(n_319)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_170),
.Y(n_268)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_268),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_214),
.B(n_16),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_269),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_153),
.B(n_16),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_137),
.Y(n_272)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_272),
.Y(n_322)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_178),
.Y(n_273)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_273),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_214),
.B(n_154),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_274),
.B(n_276),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_194),
.A2(n_52),
.B1(n_49),
.B2(n_46),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_140),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_149),
.B(n_14),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_277),
.B(n_281),
.Y(n_353)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_150),
.Y(n_278)
);

BUFx4f_ASAP7_75t_L g344 ( 
.A(n_278),
.Y(n_344)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_129),
.A2(n_14),
.B(n_13),
.C(n_52),
.Y(n_279)
);

O2A1O1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_279),
.A2(n_284),
.B(n_1),
.C(n_2),
.Y(n_316)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_162),
.Y(n_280)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_280),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_133),
.B(n_0),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_215),
.B(n_0),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_285),
.Y(n_305)
);

CKINVDCx12_ASAP7_75t_R g283 ( 
.A(n_201),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_283),
.Y(n_306)
);

OA22x2_ASAP7_75t_L g284 ( 
.A1(n_198),
.A2(n_49),
.B1(n_19),
.B2(n_2),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_139),
.B(n_0),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_142),
.B(n_0),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_287),
.B(n_290),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_161),
.B(n_1),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_145),
.Y(n_291)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_291),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_192),
.Y(n_295)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_295),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_296),
.B(n_297),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_246),
.A2(n_166),
.B1(n_208),
.B2(n_155),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_298),
.A2(n_313),
.B1(n_323),
.B2(n_334),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_289),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_299),
.B(n_348),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_220),
.A2(n_186),
.B(n_173),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_300),
.A2(n_260),
.B(n_280),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_222),
.A2(n_180),
.B1(n_166),
.B2(n_148),
.Y(n_304)
);

AO21x2_ASAP7_75t_L g390 ( 
.A1(n_304),
.A2(n_326),
.B(n_336),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_307),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_247),
.A2(n_189),
.B1(n_168),
.B2(n_191),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_309),
.Y(n_378)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_237),
.Y(n_310)
);

INVx3_ASAP7_75t_SL g373 ( 
.A(n_310),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_230),
.B(n_172),
.C(n_156),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_312),
.B(n_349),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_264),
.A2(n_225),
.B1(n_247),
.B2(n_257),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_316),
.A2(n_338),
.B1(n_284),
.B2(n_259),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_275),
.A2(n_235),
.B1(n_270),
.B2(n_190),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_269),
.A2(n_209),
.B1(n_130),
.B2(n_190),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_279),
.B(n_171),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_328),
.B(n_330),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_229),
.B(n_171),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_262),
.A2(n_195),
.B1(n_163),
.B2(n_141),
.Y(n_333)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_333),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_234),
.A2(n_163),
.B1(n_141),
.B2(n_144),
.Y(n_336)
);

OAI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_251),
.A2(n_144),
.B1(n_172),
.B2(n_156),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_197),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_293),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_238),
.A2(n_19),
.B1(n_3),
.B2(n_4),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_345),
.A2(n_259),
.B1(n_250),
.B2(n_252),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_294),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_294),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_244),
.B(n_201),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_350),
.B(n_243),
.Y(n_397)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_238),
.Y(n_351)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_351),
.Y(n_356)
);

INVx13_ASAP7_75t_L g354 ( 
.A(n_306),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_354),
.Y(n_410)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_357),
.Y(n_400)
);

INVx13_ASAP7_75t_L g358 ( 
.A(n_347),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g432 ( 
.A1(n_358),
.A2(n_361),
.B1(n_376),
.B2(n_383),
.Y(n_432)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_327),
.Y(n_359)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_359),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_360),
.A2(n_389),
.B(n_221),
.Y(n_404)
);

BUFx24_ASAP7_75t_L g361 ( 
.A(n_344),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_317),
.B(n_255),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_362),
.B(n_384),
.Y(n_406)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_327),
.Y(n_363)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_363),
.Y(n_414)
);

AND2x6_ASAP7_75t_L g366 ( 
.A(n_325),
.B(n_302),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_366),
.B(n_385),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_367),
.B(n_371),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_300),
.A2(n_278),
.B(n_291),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_369),
.A2(n_395),
.B(n_337),
.Y(n_405)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_322),
.Y(n_370)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_370),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_305),
.B(n_223),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_334),
.A2(n_236),
.B1(n_295),
.B2(n_284),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_374),
.A2(n_386),
.B1(n_387),
.B2(n_326),
.Y(n_411)
);

INVx13_ASAP7_75t_L g376 ( 
.A(n_347),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_305),
.B(n_260),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_377),
.B(n_379),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_328),
.B(n_219),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_308),
.Y(n_380)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_380),
.Y(n_419)
);

OAI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_381),
.A2(n_355),
.B1(n_378),
.B2(n_390),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_329),
.Y(n_382)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_382),
.Y(n_423)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_352),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_331),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_334),
.A2(n_286),
.B1(n_231),
.B2(n_239),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_313),
.A2(n_256),
.B1(n_273),
.B2(n_266),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_320),
.B(n_292),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_388),
.B(n_396),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_316),
.A2(n_252),
.B(n_261),
.Y(n_389)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_308),
.Y(n_391)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_391),
.Y(n_429)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_321),
.Y(n_392)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_392),
.Y(n_433)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_340),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_393),
.B(n_397),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_312),
.A2(n_261),
.B(n_243),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_321),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_398),
.B(n_329),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_390),
.A2(n_296),
.B1(n_298),
.B2(n_330),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_399),
.A2(n_407),
.B1(n_411),
.B2(n_368),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_372),
.B(n_350),
.C(n_314),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_401),
.B(n_403),
.C(n_415),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_395),
.B(n_320),
.C(n_332),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_404),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_405),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_390),
.A2(n_301),
.B1(n_336),
.B2(n_315),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_360),
.A2(n_337),
.B(n_303),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_409),
.B(n_420),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_319),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_412),
.B(n_344),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_390),
.A2(n_353),
.B1(n_304),
.B2(n_343),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_413),
.A2(n_417),
.B1(n_386),
.B2(n_396),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_393),
.B(n_364),
.C(n_377),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_416),
.B(n_356),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_390),
.A2(n_343),
.B1(n_341),
.B2(n_346),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_369),
.A2(n_303),
.B(n_339),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_371),
.B(n_324),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_422),
.B(n_435),
.C(n_356),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_364),
.A2(n_324),
.B(n_342),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_424),
.B(n_430),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_379),
.B(n_342),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g445 ( 
.A(n_427),
.B(n_422),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_355),
.A2(n_367),
.B(n_389),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_394),
.Y(n_431)
);

INVx13_ASAP7_75t_L g459 ( 
.A(n_431),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g440 ( 
.A1(n_434),
.A2(n_407),
.B1(n_399),
.B2(n_405),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_370),
.B(n_311),
.C(n_318),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_411),
.A2(n_368),
.B1(n_381),
.B2(n_365),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_436),
.B(n_442),
.Y(n_478)
);

BUFx24_ASAP7_75t_SL g437 ( 
.A(n_408),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_437),
.B(n_454),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_431),
.B(n_406),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_438),
.B(n_452),
.Y(n_482)
);

MAJx2_ASAP7_75t_L g439 ( 
.A(n_401),
.B(n_366),
.C(n_398),
.Y(n_439)
);

FAx1_ASAP7_75t_SL g500 ( 
.A(n_439),
.B(n_376),
.CI(n_358),
.CON(n_500),
.SN(n_500)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_440),
.A2(n_446),
.B1(n_448),
.B2(n_456),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_374),
.Y(n_444)
);

AO21x1_ASAP7_75t_L g481 ( 
.A1(n_444),
.A2(n_458),
.B(n_404),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_445),
.B(n_469),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_415),
.B(n_368),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_460),
.C(n_423),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_425),
.A2(n_378),
.B1(n_375),
.B2(n_373),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_418),
.Y(n_450)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_450),
.Y(n_474)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_418),
.Y(n_451)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_451),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_416),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_406),
.B(n_335),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_402),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_457),
.B(n_419),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_409),
.B(n_391),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_402),
.B(n_311),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_413),
.A2(n_375),
.B1(n_373),
.B2(n_380),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_461),
.A2(n_432),
.B1(n_410),
.B2(n_423),
.Y(n_471)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_400),
.Y(n_462)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_462),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_425),
.A2(n_375),
.B1(n_341),
.B2(n_310),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_463),
.B(n_428),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_403),
.B(n_335),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_464),
.B(n_465),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_426),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_421),
.B(n_363),
.Y(n_467)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_467),
.Y(n_475)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_400),
.Y(n_468)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_468),
.Y(n_488)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_354),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_471),
.B(n_473),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_472),
.B(n_439),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_442),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_476),
.B(n_477),
.C(n_496),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_421),
.C(n_424),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_459),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_479),
.B(n_487),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_481),
.A2(n_490),
.B(n_428),
.Y(n_526)
);

OA22x2_ASAP7_75t_L g483 ( 
.A1(n_466),
.A2(n_417),
.B1(n_375),
.B2(n_410),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_483),
.Y(n_510)
);

XNOR2x1_ASAP7_75t_L g484 ( 
.A(n_447),
.B(n_426),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_484),
.B(n_489),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_456),
.A2(n_427),
.B1(n_433),
.B2(n_429),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_486),
.A2(n_499),
.B1(n_501),
.B2(n_462),
.Y(n_522)
);

NOR2x1_ASAP7_75t_L g487 ( 
.A(n_467),
.B(n_433),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_453),
.B(n_435),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_443),
.A2(n_410),
.B(n_414),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_450),
.Y(n_491)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_491),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_414),
.Y(n_492)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_492),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_449),
.Y(n_494)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_494),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_455),
.B(n_429),
.C(n_419),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_451),
.Y(n_497)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_497),
.Y(n_517)
);

AOI21xp33_ASAP7_75t_L g523 ( 
.A1(n_500),
.A2(n_346),
.B(n_339),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_496),
.C(n_477),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_505),
.B(n_511),
.C(n_513),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_478),
.A2(n_466),
.B1(n_443),
.B2(n_444),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_506),
.A2(n_521),
.B1(n_490),
.B2(n_495),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_507),
.B(n_512),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_472),
.B(n_445),
.C(n_436),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_476),
.B(n_444),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_484),
.B(n_441),
.C(n_458),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_482),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_514),
.B(n_515),
.Y(n_549)
);

NOR3xp33_ASAP7_75t_SL g515 ( 
.A(n_485),
.B(n_459),
.C(n_469),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_498),
.B(n_441),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_518),
.B(n_475),
.Y(n_544)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_487),
.Y(n_519)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_519),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_492),
.B(n_441),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_520),
.B(n_486),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_478),
.A2(n_461),
.B1(n_458),
.B2(n_468),
.Y(n_521)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_522),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_523),
.A2(n_499),
.B(n_500),
.Y(n_536)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_491),
.Y(n_524)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_524),
.Y(n_545)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_470),
.Y(n_525)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_525),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_526),
.A2(n_481),
.B(n_501),
.Y(n_542)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_497),
.Y(n_528)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_528),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_516),
.A2(n_485),
.B1(n_510),
.B2(n_527),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_529),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_530),
.B(n_542),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_518),
.B(n_493),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_535),
.B(n_541),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_536),
.B(n_544),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_508),
.B(n_475),
.Y(n_537)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_537),
.Y(n_552)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_525),
.Y(n_539)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_539),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_540),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_502),
.B(n_474),
.Y(n_541)
);

CKINVDCx14_ASAP7_75t_R g543 ( 
.A(n_509),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_543),
.B(n_546),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_505),
.B(n_483),
.C(n_471),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_502),
.B(n_483),
.C(n_480),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_547),
.B(n_506),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_510),
.A2(n_500),
.B1(n_488),
.B2(n_470),
.Y(n_550)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_550),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_547),
.B(n_511),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_551),
.B(n_553),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_534),
.B(n_512),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_532),
.B(n_503),
.C(n_507),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_556),
.B(n_562),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_538),
.B(n_503),
.Y(n_561)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_561),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_532),
.B(n_513),
.C(n_526),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_549),
.B(n_504),
.Y(n_563)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_563),
.Y(n_578)
);

OAI21x1_ASAP7_75t_L g577 ( 
.A1(n_565),
.A2(n_550),
.B(n_533),
.Y(n_577)
);

BUFx12_ASAP7_75t_L g567 ( 
.A(n_530),
.Y(n_567)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_567),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_562),
.B(n_546),
.C(n_531),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_568),
.B(n_570),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_556),
.B(n_531),
.C(n_540),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_558),
.B(n_542),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_571),
.B(n_573),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_559),
.B(n_544),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_552),
.B(n_536),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_574),
.A2(n_581),
.B1(n_545),
.B2(n_517),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_557),
.B(n_548),
.Y(n_575)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_575),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_554),
.B(n_564),
.C(n_558),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_576),
.B(n_555),
.C(n_566),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_577),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_SL g579 ( 
.A(n_559),
.B(n_520),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_579),
.B(n_567),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_555),
.A2(n_515),
.B1(n_537),
.B2(n_539),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_SL g583 ( 
.A1(n_582),
.A2(n_566),
.B(n_560),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_583),
.B(n_584),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_569),
.B(n_533),
.C(n_521),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_585),
.B(n_594),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_587),
.B(n_288),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_570),
.B(n_567),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_589),
.B(n_593),
.C(n_361),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_590),
.A2(n_576),
.B1(n_568),
.B2(n_579),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_571),
.B(n_483),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_SL g594 ( 
.A1(n_574),
.A2(n_488),
.B(n_359),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_586),
.A2(n_578),
.B1(n_572),
.B2(n_580),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_595),
.B(n_599),
.Y(n_606)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_596),
.Y(n_608)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_586),
.A2(n_318),
.B(n_361),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_597),
.A2(n_602),
.B(n_344),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_588),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_600),
.B(n_601),
.Y(n_607)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_592),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_604),
.A2(n_609),
.B(n_245),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_SL g605 ( 
.A(n_603),
.B(n_591),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_605),
.A2(n_587),
.B1(n_602),
.B2(n_593),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_596),
.A2(n_589),
.B(n_585),
.Y(n_609)
);

A2O1A1Ixp33_ASAP7_75t_SL g610 ( 
.A1(n_607),
.A2(n_608),
.B(n_606),
.C(n_598),
.Y(n_610)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_610),
.A2(n_611),
.B(n_612),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_612),
.B(n_221),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_614),
.A2(n_288),
.B(n_3),
.Y(n_615)
);

AO21x1_ASAP7_75t_L g616 ( 
.A1(n_615),
.A2(n_613),
.B(n_4),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_616),
.B(n_2),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_617),
.B(n_9),
.C(n_6),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_618),
.Y(n_619)
);


endmodule