module real_aes_2570_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_594;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_231;
wire n_547;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_246;
wire n_412;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_613;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_498;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_294;
wire n_393;
wire n_258;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_0), .A2(n_194), .B1(n_372), .B2(n_396), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_1), .A2(n_87), .B1(n_334), .B2(n_337), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_2), .A2(n_117), .B1(n_371), .B2(n_372), .Y(n_492) );
AO22x2_ASAP7_75t_L g247 ( .A1(n_3), .A2(n_161), .B1(n_248), .B2(n_249), .Y(n_247) );
INVx1_ASAP7_75t_L g584 ( .A(n_3), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_4), .A2(n_164), .B1(n_312), .B2(n_316), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_5), .A2(n_133), .B1(n_420), .B2(n_422), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_6), .A2(n_111), .B1(n_368), .B2(n_369), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_7), .A2(n_193), .B1(n_307), .B2(n_436), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_8), .A2(n_56), .B1(n_542), .B2(n_543), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_9), .A2(n_110), .B1(n_268), .B2(n_274), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_10), .A2(n_106), .B1(n_385), .B2(n_388), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_11), .A2(n_85), .B1(n_276), .B2(n_331), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_12), .A2(n_55), .B1(n_387), .B2(n_388), .Y(n_386) );
OA22x2_ASAP7_75t_L g389 ( .A1(n_13), .A2(n_390), .B1(n_391), .B2(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_13), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_14), .A2(n_47), .B1(n_303), .B2(n_307), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_15), .A2(n_26), .B1(n_384), .B2(n_387), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_16), .A2(n_79), .B1(n_385), .B2(n_388), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_17), .A2(n_163), .B1(n_378), .B2(n_379), .Y(n_498) );
AO22x2_ASAP7_75t_L g251 ( .A1(n_18), .A2(n_53), .B1(n_248), .B2(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_18), .B(n_583), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_19), .A2(n_41), .B1(n_384), .B2(n_385), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_20), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_21), .A2(n_131), .B1(n_387), .B2(n_388), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_22), .A2(n_118), .B1(n_320), .B2(n_427), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_23), .A2(n_48), .B1(n_340), .B2(n_344), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_24), .A2(n_82), .B1(n_348), .B2(n_439), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_25), .A2(n_206), .B1(n_384), .B2(n_387), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_27), .A2(n_50), .B1(n_520), .B2(n_604), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_28), .A2(n_67), .B1(n_439), .B2(n_478), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_29), .A2(n_49), .B1(n_381), .B2(n_382), .Y(n_402) );
AOI222xp33_ASAP7_75t_L g394 ( .A1(n_30), .A2(n_195), .B1(n_217), .B2(n_366), .C1(n_395), .C2(n_396), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_31), .A2(n_176), .B1(n_378), .B2(n_379), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_32), .A2(n_221), .B1(n_385), .B2(n_388), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_33), .A2(n_198), .B1(n_384), .B2(n_385), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_34), .A2(n_103), .B1(n_385), .B2(n_388), .Y(n_403) );
AO22x1_ASAP7_75t_L g518 ( .A1(n_35), .A2(n_166), .B1(n_519), .B2(n_520), .Y(n_518) );
OA22x2_ASAP7_75t_L g508 ( .A1(n_36), .A2(n_509), .B1(n_510), .B2(n_533), .Y(n_508) );
INVx1_ASAP7_75t_L g533 ( .A(n_36), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_37), .A2(n_138), .B1(n_595), .B2(n_596), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_38), .A2(n_93), .B1(n_382), .B2(n_454), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_39), .A2(n_100), .B1(n_372), .B2(n_396), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_40), .A2(n_148), .B1(n_371), .B2(n_372), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_42), .A2(n_92), .B1(n_433), .B2(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_43), .B(n_366), .Y(n_490) );
AOI22xp33_ASAP7_75t_SL g399 ( .A1(n_44), .A2(n_219), .B1(n_374), .B2(n_400), .Y(n_399) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_45), .A2(n_178), .B1(n_382), .B2(n_387), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_46), .A2(n_109), .B1(n_430), .B2(n_433), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_51), .A2(n_66), .B1(n_374), .B2(n_375), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_52), .A2(n_81), .B1(n_352), .B2(n_513), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_54), .A2(n_99), .B1(n_371), .B2(n_372), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_57), .A2(n_155), .B1(n_244), .B2(n_261), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_58), .A2(n_209), .B1(n_374), .B2(n_375), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_59), .A2(n_218), .B1(n_378), .B2(n_379), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_60), .A2(n_123), .B1(n_420), .B2(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_61), .A2(n_102), .B1(n_368), .B2(n_398), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_62), .A2(n_91), .B1(n_598), .B2(n_599), .Y(n_597) );
INVx3_ASAP7_75t_L g248 ( .A(n_63), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_64), .A2(n_77), .B1(n_331), .B2(n_332), .Y(n_330) );
XOR2x1_ASAP7_75t_L g410 ( .A(n_65), .B(n_411), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_68), .A2(n_145), .B1(n_414), .B2(n_417), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_69), .A2(n_121), .B1(n_322), .B2(n_348), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_70), .A2(n_136), .B1(n_319), .B2(n_354), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_71), .A2(n_216), .B1(n_307), .B2(n_436), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_72), .A2(n_147), .B1(n_381), .B2(n_382), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_73), .B(n_424), .Y(n_423) );
XOR2x2_ASAP7_75t_L g487 ( .A(n_74), .B(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_75), .B(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_76), .A2(n_177), .B1(n_374), .B2(n_375), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_78), .A2(n_144), .B1(n_378), .B2(n_379), .Y(n_622) );
INVx1_ASAP7_75t_SL g256 ( .A(n_80), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_80), .B(n_108), .Y(n_585) );
INVx2_ASAP7_75t_L g232 ( .A(n_83), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_84), .A2(n_120), .B1(n_427), .B2(n_428), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_86), .A2(n_220), .B1(n_382), .B2(n_454), .Y(n_453) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_88), .A2(n_223), .B(n_233), .C(n_586), .Y(n_222) );
XOR2x2_ASAP7_75t_L g559 ( .A(n_89), .B(n_560), .Y(n_559) );
XOR2x2_ASAP7_75t_L g240 ( .A(n_90), .B(n_241), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_94), .A2(n_105), .B1(n_384), .B2(n_454), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_95), .A2(n_114), .B1(n_414), .B2(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_96), .B(n_424), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_97), .A2(n_129), .B1(n_319), .B2(n_322), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_98), .A2(n_115), .B1(n_354), .B2(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_101), .A2(n_202), .B1(n_368), .B2(n_369), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_104), .A2(n_192), .B1(n_381), .B2(n_382), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_107), .B(n_366), .Y(n_365) );
AO22x2_ASAP7_75t_L g259 ( .A1(n_108), .A2(n_167), .B1(n_248), .B2(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_112), .B(n_366), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_113), .A2(n_186), .B1(n_342), .B2(n_414), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_116), .A2(n_185), .B1(n_374), .B2(n_375), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_119), .A2(n_182), .B1(n_417), .B2(n_418), .Y(n_416) );
AO22x1_ASAP7_75t_L g515 ( .A1(n_122), .A2(n_154), .B1(n_516), .B2(n_517), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_124), .Y(n_466) );
AO22x1_ASAP7_75t_L g521 ( .A1(n_125), .A2(n_158), .B1(n_313), .B2(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g257 ( .A(n_126), .Y(n_257) );
AOI22xp33_ASAP7_75t_SL g473 ( .A1(n_127), .A2(n_174), .B1(n_379), .B2(n_474), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_128), .A2(n_190), .B1(n_374), .B2(n_400), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_130), .A2(n_152), .B1(n_378), .B2(n_379), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_132), .A2(n_197), .B1(n_342), .B2(n_369), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_134), .A2(n_188), .B1(n_321), .B2(n_566), .Y(n_565) );
AOI22xp33_ASAP7_75t_SL g469 ( .A1(n_135), .A2(n_215), .B1(n_368), .B2(n_369), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_137), .A2(n_159), .B1(n_378), .B2(n_379), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_139), .A2(n_169), .B1(n_378), .B2(n_379), .Y(n_452) );
INVx1_ASAP7_75t_L g326 ( .A(n_140), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_141), .A2(n_210), .B1(n_279), .B2(n_282), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_142), .A2(n_187), .B1(n_358), .B2(n_430), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_143), .A2(n_151), .B1(n_295), .B2(n_298), .Y(n_294) );
XNOR2x1_ASAP7_75t_L g362 ( .A(n_146), .B(n_363), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_149), .A2(n_170), .B1(n_517), .B2(n_566), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_150), .A2(n_179), .B1(n_368), .B2(n_398), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_153), .A2(n_211), .B1(n_368), .B2(n_398), .Y(n_397) );
AOI21xp5_ASAP7_75t_SL g524 ( .A1(n_156), .A2(n_525), .B(n_526), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_157), .A2(n_212), .B1(n_357), .B2(n_358), .Y(n_356) );
CKINVDCx16_ASAP7_75t_R g627 ( .A(n_160), .Y(n_627) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_162), .A2(n_203), .B1(n_279), .B2(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g458 ( .A(n_165), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_168), .A2(n_175), .B1(n_348), .B2(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_171), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_172), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_173), .B(n_287), .Y(n_286) );
XOR2x2_ASAP7_75t_L g534 ( .A(n_180), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_181), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g580 ( .A(n_181), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_183), .A2(n_204), .B1(n_395), .B2(n_396), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_184), .A2(n_213), .B1(n_337), .B2(n_421), .Y(n_593) );
INVx1_ASAP7_75t_L g229 ( .A(n_189), .Y(n_229) );
AND2x2_ASAP7_75t_R g610 ( .A(n_189), .B(n_580), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_191), .A2(n_588), .B1(n_589), .B2(n_608), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_191), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_196), .A2(n_207), .B1(n_350), .B2(n_352), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_199), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_200), .B(n_287), .Y(n_329) );
INVx1_ASAP7_75t_L g480 ( .A(n_201), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_205), .B(n_366), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_208), .A2(n_214), .B1(n_385), .B2(n_388), .Y(n_562) );
CKINVDCx6p67_ASAP7_75t_R g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
BUFx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_SL g226 ( .A(n_227), .B(n_230), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
OR2x2_ASAP7_75t_L g631 ( .A(n_228), .B(n_230), .Y(n_631) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_229), .B(n_580), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_501), .B1(n_575), .B2(n_576), .C(n_577), .Y(n_233) );
INVxp67_ASAP7_75t_SL g575 ( .A(n_234), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_486), .B1(n_499), .B2(n_500), .Y(n_234) );
INVx1_ASAP7_75t_L g500 ( .A(n_235), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_409), .B1(n_484), .B2(n_485), .Y(n_235) );
INVx1_ASAP7_75t_L g484 ( .A(n_236), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_360), .B1(n_361), .B2(n_408), .Y(n_236) );
INVx1_ASAP7_75t_L g408 ( .A(n_237), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B1(n_325), .B2(n_359), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
BUFx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp67_ASAP7_75t_L g241 ( .A(n_242), .B(n_293), .Y(n_241) );
NAND4xp25_ASAP7_75t_L g242 ( .A(n_243), .B(n_267), .C(n_278), .D(n_286), .Y(n_242) );
BUFx6f_ASAP7_75t_SL g525 ( .A(n_244), .Y(n_525) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx3_ASAP7_75t_L g343 ( .A(n_245), .Y(n_343) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_245), .Y(n_598) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_253), .Y(n_245) );
AND2x4_ASAP7_75t_L g300 ( .A(n_246), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g306 ( .A(n_246), .B(n_272), .Y(n_306) );
AND2x4_ASAP7_75t_L g368 ( .A(n_246), .B(n_253), .Y(n_368) );
AND2x2_ASAP7_75t_L g378 ( .A(n_246), .B(n_272), .Y(n_378) );
AND2x6_ASAP7_75t_L g388 ( .A(n_246), .B(n_301), .Y(n_388) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_250), .Y(n_246) );
INVx2_ASAP7_75t_L g271 ( .A(n_247), .Y(n_271) );
AND2x2_ASAP7_75t_L g284 ( .A(n_247), .B(n_251), .Y(n_284) );
INVx1_ASAP7_75t_L g249 ( .A(n_248), .Y(n_249) );
INVx2_ASAP7_75t_L g252 ( .A(n_248), .Y(n_252) );
OAI22x1_ASAP7_75t_L g254 ( .A1(n_248), .A2(n_255), .B1(n_256), .B2(n_257), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_248), .Y(n_255) );
INVx1_ASAP7_75t_L g260 ( .A(n_248), .Y(n_260) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_250), .Y(n_266) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x4_ASAP7_75t_L g270 ( .A(n_251), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g292 ( .A(n_251), .Y(n_292) );
AND2x2_ASAP7_75t_L g281 ( .A(n_253), .B(n_270), .Y(n_281) );
AND2x4_ASAP7_75t_L g324 ( .A(n_253), .B(n_291), .Y(n_324) );
AND2x4_ASAP7_75t_L g374 ( .A(n_253), .B(n_270), .Y(n_374) );
AND2x2_ASAP7_75t_L g381 ( .A(n_253), .B(n_291), .Y(n_381) );
AND2x2_ASAP7_75t_L g454 ( .A(n_253), .B(n_291), .Y(n_454) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_258), .Y(n_253) );
AND2x2_ASAP7_75t_L g264 ( .A(n_254), .B(n_259), .Y(n_264) );
INVx2_ASAP7_75t_L g273 ( .A(n_254), .Y(n_273) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_254), .Y(n_285) );
AND2x4_ASAP7_75t_L g301 ( .A(n_258), .B(n_273), .Y(n_301) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g272 ( .A(n_259), .B(n_273), .Y(n_272) );
BUFx2_ASAP7_75t_L g310 ( .A(n_259), .Y(n_310) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
BUFx2_ASAP7_75t_L g345 ( .A(n_262), .Y(n_345) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx3_ASAP7_75t_L g415 ( .A(n_263), .Y(n_415) );
INVx1_ASAP7_75t_L g600 ( .A(n_263), .Y(n_600) );
AND2x4_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
AND2x4_ASAP7_75t_L g276 ( .A(n_264), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g290 ( .A(n_264), .B(n_291), .Y(n_290) );
AND2x4_ASAP7_75t_L g366 ( .A(n_264), .B(n_291), .Y(n_366) );
AND2x2_ASAP7_75t_L g369 ( .A(n_264), .B(n_265), .Y(n_369) );
AND2x2_ASAP7_75t_L g372 ( .A(n_264), .B(n_277), .Y(n_372) );
AND2x2_ASAP7_75t_L g395 ( .A(n_264), .B(n_277), .Y(n_395) );
AND2x2_ASAP7_75t_L g398 ( .A(n_264), .B(n_265), .Y(n_398) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
BUFx2_ASAP7_75t_L g331 ( .A(n_268), .Y(n_331) );
BUFx2_ASAP7_75t_L g417 ( .A(n_268), .Y(n_417) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx2_ASAP7_75t_L g595 ( .A(n_269), .Y(n_595) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
AND2x4_ASAP7_75t_L g321 ( .A(n_270), .B(n_301), .Y(n_321) );
AND2x2_ASAP7_75t_L g371 ( .A(n_270), .B(n_272), .Y(n_371) );
AND2x2_ASAP7_75t_L g384 ( .A(n_270), .B(n_301), .Y(n_384) );
AND2x2_ASAP7_75t_L g396 ( .A(n_270), .B(n_272), .Y(n_396) );
INVxp67_ASAP7_75t_L g277 ( .A(n_271), .Y(n_277) );
AND2x4_ASAP7_75t_L g291 ( .A(n_271), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g297 ( .A(n_272), .B(n_291), .Y(n_297) );
AND2x6_ASAP7_75t_L g385 ( .A(n_272), .B(n_291), .Y(n_385) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g332 ( .A(n_275), .Y(n_332) );
INVx2_ASAP7_75t_L g418 ( .A(n_275), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_275), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_SL g596 ( .A(n_275), .Y(n_596) );
INVx6_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx3_ASAP7_75t_L g336 ( .A(n_281), .Y(n_336) );
BUFx3_ASAP7_75t_L g421 ( .A(n_281), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_282), .Y(n_422) );
INVx2_ASAP7_75t_L g532 ( .A(n_282), .Y(n_532) );
BUFx12f_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx3_ASAP7_75t_L g338 ( .A(n_283), .Y(n_338) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x4_ASAP7_75t_L g309 ( .A(n_284), .B(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g317 ( .A(n_284), .B(n_301), .Y(n_317) );
AND2x2_ASAP7_75t_SL g375 ( .A(n_284), .B(n_285), .Y(n_375) );
AND2x4_ASAP7_75t_L g379 ( .A(n_284), .B(n_310), .Y(n_379) );
AND2x4_ASAP7_75t_L g382 ( .A(n_284), .B(n_301), .Y(n_382) );
AND2x2_ASAP7_75t_SL g400 ( .A(n_284), .B(n_285), .Y(n_400) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g546 ( .A(n_288), .Y(n_546) );
INVx3_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
INVx3_ASAP7_75t_L g424 ( .A(n_289), .Y(n_424) );
INVx4_ASAP7_75t_SL g574 ( .A(n_289), .Y(n_574) );
INVx4_ASAP7_75t_SL g592 ( .A(n_289), .Y(n_592) );
INVx6_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g315 ( .A(n_291), .B(n_301), .Y(n_315) );
AND2x2_ASAP7_75t_L g387 ( .A(n_291), .B(n_301), .Y(n_387) );
NAND4xp25_ASAP7_75t_L g293 ( .A(n_294), .B(n_302), .C(n_311), .D(n_318), .Y(n_293) );
INVx2_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_SL g357 ( .A(n_296), .Y(n_357) );
INVx3_ASAP7_75t_L g606 ( .A(n_296), .Y(n_606) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
BUFx2_ASAP7_75t_L g432 ( .A(n_297), .Y(n_432) );
BUFx2_ASAP7_75t_L g516 ( .A(n_297), .Y(n_516) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g358 ( .A(n_299), .Y(n_358) );
INVx2_ASAP7_75t_SL g428 ( .A(n_299), .Y(n_428) );
INVx2_ASAP7_75t_L g517 ( .A(n_299), .Y(n_517) );
INVx8_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g351 ( .A(n_304), .Y(n_351) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_304), .Y(n_513) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g437 ( .A(n_305), .Y(n_437) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx3_ASAP7_75t_L g474 ( .A(n_306), .Y(n_474) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx5_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
BUFx2_ASAP7_75t_L g352 ( .A(n_309), .Y(n_352) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g355 ( .A(n_313), .Y(n_355) );
INVx4_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx3_ASAP7_75t_SL g427 ( .A(n_314), .Y(n_427) );
INVx3_ASAP7_75t_L g566 ( .A(n_314), .Y(n_566) );
INVx8_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx2_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
BUFx2_ASAP7_75t_SL g348 ( .A(n_317), .Y(n_348) );
BUFx3_ASAP7_75t_L g478 ( .A(n_317), .Y(n_478) );
BUFx3_ASAP7_75t_L g520 ( .A(n_317), .Y(n_520) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g552 ( .A(n_320), .Y(n_552) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g434 ( .A(n_321), .Y(n_434) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g519 ( .A(n_323), .Y(n_519) );
INVx1_ASAP7_75t_SL g554 ( .A(n_323), .Y(n_554) );
INVx6_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx3_ASAP7_75t_L g439 ( .A(n_324), .Y(n_439) );
BUFx3_ASAP7_75t_L g604 ( .A(n_324), .Y(n_604) );
INVx2_ASAP7_75t_L g359 ( .A(n_325), .Y(n_359) );
XNOR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
NOR2x1_ASAP7_75t_L g327 ( .A(n_328), .B(n_346), .Y(n_327) );
NAND4xp25_ASAP7_75t_SL g328 ( .A(n_329), .B(n_330), .C(n_333), .D(n_339), .Y(n_328) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx6f_ASAP7_75t_SL g542 ( .A(n_336), .Y(n_542) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_337), .Y(n_543) );
INVx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g569 ( .A(n_338), .Y(n_569) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVx4_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g539 ( .A(n_343), .Y(n_539) );
INVx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND4xp25_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .C(n_353), .D(n_356), .Y(n_346) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AO22x2_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_389), .B1(n_406), .B2(n_407), .Y(n_361) );
INVx1_ASAP7_75t_L g406 ( .A(n_362), .Y(n_406) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_376), .Y(n_363) );
NAND4xp25_ASAP7_75t_SL g364 ( .A(n_365), .B(n_367), .C(n_370), .D(n_373), .Y(n_364) );
INVx2_ASAP7_75t_SL g465 ( .A(n_366), .Y(n_465) );
NAND4xp25_ASAP7_75t_SL g376 ( .A(n_377), .B(n_380), .C(n_383), .D(n_386), .Y(n_376) );
INVx1_ASAP7_75t_L g407 ( .A(n_389), .Y(n_407) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_393), .B(n_401), .Y(n_392) );
NAND3xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_397), .C(n_399), .Y(n_393) );
NAND4xp25_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .C(n_404), .D(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g485 ( .A(n_409), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_440), .B1(n_482), .B2(n_483), .Y(n_409) );
INVx1_ASAP7_75t_SL g482 ( .A(n_410), .Y(n_482) );
OR2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_425), .Y(n_411) );
NAND4xp25_ASAP7_75t_L g412 ( .A(n_413), .B(n_416), .C(n_419), .D(n_423), .Y(n_412) );
BUFx6f_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND4xp25_ASAP7_75t_L g425 ( .A(n_426), .B(n_429), .C(n_435), .D(n_438), .Y(n_425) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g522 ( .A(n_434), .Y(n_522) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g483 ( .A(n_440), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_459), .B1(n_460), .B2(n_481), .Y(n_440) );
INVx3_ASAP7_75t_SL g481 ( .A(n_441), .Y(n_481) );
XOR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_458), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_450), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_447), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_445), .B(n_446), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_455), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
XOR2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_480), .Y(n_461) );
NAND2x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_471), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_468), .Y(n_463) );
OAI21xp5_ASAP7_75t_SL g464 ( .A1(n_465), .A2(n_466), .B(n_467), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_472), .B(n_476), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_475), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_479), .Y(n_476) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_487), .Y(n_499) );
NOR2x1_ASAP7_75t_L g488 ( .A(n_489), .B(n_494), .Y(n_488) );
NAND4xp25_ASAP7_75t_SL g489 ( .A(n_490), .B(n_491), .C(n_492), .D(n_493), .Y(n_489) );
NAND4xp25_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .C(n_497), .D(n_498), .Y(n_494) );
INVx1_ASAP7_75t_L g576 ( .A(n_501), .Y(n_576) );
AOI22xp5_ASAP7_75t_SL g501 ( .A1(n_502), .A2(n_503), .B1(n_556), .B2(n_557), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B1(n_534), .B2(n_555), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NOR2xp67_ASAP7_75t_L g510 ( .A(n_511), .B(n_523), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_514), .Y(n_511) );
NOR3xp33_ASAP7_75t_L g514 ( .A(n_515), .B(n_518), .C(n_521), .Y(n_514) );
NAND4xp25_ASAP7_75t_L g523 ( .A(n_524), .B(n_528), .C(n_529), .D(n_530), .Y(n_523) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx4_ASAP7_75t_L g555 ( .A(n_534), .Y(n_555) );
NOR2x1_ASAP7_75t_L g535 ( .A(n_536), .B(n_547), .Y(n_535) );
NAND4xp25_ASAP7_75t_L g536 ( .A(n_537), .B(n_540), .C(n_541), .D(n_544), .Y(n_536) );
BUFx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND4xp25_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .C(n_550), .D(n_553), .Y(n_547) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NOR3xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_567), .C(n_571), .Y(n_560) );
NAND4xp25_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .C(n_564), .D(n_565), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
INVx3_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_579), .B(n_582), .Y(n_630) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
OAI222xp33_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_609), .B1(n_611), .B2(n_627), .C1(n_628), .C2(n_631), .Y(n_586) );
INVxp67_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_601), .Y(n_589) );
NAND4xp25_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .C(n_594), .D(n_597), .Y(n_590) );
INVx2_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
NAND4xp25_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .C(n_605), .D(n_607), .Y(n_601) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
XOR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_627), .Y(n_611) );
NAND2x1p5_ASAP7_75t_L g612 ( .A(n_613), .B(n_620), .Y(n_612) );
NOR2x1_ASAP7_75t_L g613 ( .A(n_614), .B(n_617), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
NOR2x1_ASAP7_75t_L g620 ( .A(n_621), .B(n_624), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_629), .Y(n_628) );
CKINVDCx6p67_ASAP7_75t_R g629 ( .A(n_630), .Y(n_629) );
endmodule