module real_jpeg_27840_n_12 (n_5, n_4, n_8, n_0, n_315, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_315;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_0),
.A2(n_6),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_0),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_0),
.A2(n_21),
.B1(n_46),
.B2(n_48),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_0),
.A2(n_21),
.B1(n_40),
.B2(n_44),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_1),
.B(n_48),
.Y(n_109)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_1),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_1),
.B(n_208),
.Y(n_213)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_1),
.Y(n_224)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_4),
.A2(n_6),
.B1(n_20),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_4),
.A2(n_31),
.B1(n_46),
.B2(n_48),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_4),
.A2(n_31),
.B1(n_40),
.B2(n_44),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_5),
.A2(n_40),
.B1(n_44),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_52),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_5),
.A2(n_20),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_5),
.B(n_20),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_5),
.B(n_71),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_5),
.A2(n_46),
.B1(n_48),
.B2(n_52),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_SL g168 ( 
.A1(n_5),
.A2(n_10),
.B(n_40),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_L g198 ( 
.A1(n_5),
.A2(n_7),
.B(n_46),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_5),
.B(n_56),
.Y(n_202)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_6),
.A2(n_8),
.B1(n_20),
.B2(n_123),
.Y(n_122)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_8),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_123),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_8),
.A2(n_40),
.B1(n_44),
.B2(n_123),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_8),
.A2(n_46),
.B1(n_48),
.B2(n_123),
.Y(n_208)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_11),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_99),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_97),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_84),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_15),
.B(n_84),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_69),
.C(n_77),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_16),
.A2(n_17),
.B1(n_69),
.B2(n_302),
.Y(n_307)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_34),
.B1(n_35),
.B2(n_68),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_18),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_22),
.B(n_28),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_19),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_20),
.A2(n_22),
.B(n_23),
.C(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_22),
.B(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_22),
.A2(n_32),
.B(n_75),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_22)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_24),
.B(n_27),
.Y(n_140)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_25),
.A2(n_56),
.B(n_64),
.C(n_65),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_25),
.B(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_25),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_25),
.A2(n_52),
.B(n_66),
.C(n_168),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_29),
.B(n_121),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_30),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_32),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_33),
.Y(n_142)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_53),
.Y(n_35)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_36),
.B(n_53),
.C(n_68),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_36),
.A2(n_78),
.B1(n_124),
.B2(n_125),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_36),
.B(n_79),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_49),
.B(n_50),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_37),
.A2(n_116),
.B(n_250),
.Y(n_276)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_38),
.B(n_51),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_38),
.B(n_117),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_38),
.B(n_178),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_45),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_40),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_44),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_40),
.A2(n_42),
.B(n_52),
.C(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_45),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_45),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_45),
.B(n_51),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_46),
.Y(n_48)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_48),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_49),
.B(n_52),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_49),
.A2(n_179),
.B(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_52),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_61),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_54),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_59),
.B(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_55),
.A2(n_62),
.B(n_81),
.Y(n_287)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_56),
.B(n_127),
.Y(n_126)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_60),
.B(n_63),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_62),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_80),
.B(n_82),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_63),
.B(n_127),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_78),
.C(n_79),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_69),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_69),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_70),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_71),
.B(n_270),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_75),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_77),
.B(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_120),
.C(n_124),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_82),
.B(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_83),
.B(n_137),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_91),
.B2(n_93),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B(n_90),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_88),
.B(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_91),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_91),
.A2(n_93),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_93),
.B(n_252),
.C(n_255),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI321xp33_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_299),
.A3(n_308),
.B1(n_311),
.B2(n_312),
.C(n_315),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_280),
.B(n_298),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_259),
.B(n_279),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_161),
.B(n_242),
.C(n_258),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_148),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_104),
.B(n_148),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_128),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_119),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_106),
.B(n_119),
.C(n_128),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_115),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_107),
.B(n_115),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_110),
.B(n_111),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_108),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_109),
.A2(n_113),
.B(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_109),
.B(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_111),
.B(n_207),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_113),
.B(n_160),
.Y(n_206)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_116),
.B(n_189),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_118),
.B(n_177),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_138),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_134),
.B2(n_135),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_130),
.B(n_135),
.C(n_138),
.Y(n_256)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_132),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_143),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_145),
.B(n_206),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_146),
.B(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_154),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_149),
.A2(n_150),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_154),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.C(n_158),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_158),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_159),
.B(n_213),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_241),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_234),
.B(n_240),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_191),
.B(n_233),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_180),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_165),
.B(n_180),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_172),
.C(n_175),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_166),
.B(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_167),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_170),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_169),
.A2(n_170),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_169),
.B(n_276),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_169),
.A2(n_170),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_170),
.A2(n_290),
.B(n_295),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_231)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_174),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_179),
.B(n_188),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_181),
.B(n_187),
.C(n_190),
.Y(n_235)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_228),
.B(n_232),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_209),
.B(n_227),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_194),
.B(n_199),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_197),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_204),
.C(n_205),
.Y(n_229)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_216),
.B(n_226),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_211),
.B(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_220),
.B(n_225),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_218),
.B(n_219),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_229),
.B(n_230),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_235),
.B(n_236),
.Y(n_240)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_243),
.B(n_244),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_256),
.B2(n_257),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_251),
.C(n_257),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_249),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_256),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_260),
.B(n_261),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_278),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_274),
.B2(n_275),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_275),
.C(n_278),
.Y(n_281)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_267),
.C(n_272),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_271),
.B2(n_272),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_276),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_281),
.B(n_282),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_296),
.B2(n_297),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_289),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_289),
.C(n_297),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B(n_288),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_287),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_301),
.C(n_305),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_288),
.B(n_301),
.CI(n_305),
.CON(n_310),
.SN(n_310)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_296),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_306),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_306),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_309),
.B(n_310),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_310),
.Y(n_313)
);


endmodule