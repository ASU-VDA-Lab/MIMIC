module fake_jpeg_21362_n_95 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_95);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_95;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_8),
.Y(n_27)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_20),
.B(n_8),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_27),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_20),
.B(n_22),
.C(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_35),
.Y(n_41)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_19),
.B1(n_21),
.B2(n_17),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_24),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_12),
.B(n_13),
.C(n_21),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_23),
.A2(n_19),
.B1(n_21),
.B2(n_15),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_23),
.B1(n_28),
.B2(n_26),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_19),
.B(n_17),
.Y(n_38)
);

AO21x1_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_40),
.B(n_44),
.Y(n_45)
);

AOI31xp33_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_12),
.A3(n_17),
.B(n_10),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_32),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_28),
.B1(n_36),
.B2(n_33),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_46),
.B(n_50),
.Y(n_60)
);

AO21x1_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_30),
.B(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_49),
.B(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_9),
.Y(n_63)
);

NAND4xp25_ASAP7_75t_SL g57 ( 
.A(n_45),
.B(n_25),
.C(n_42),
.D(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_40),
.C(n_16),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_16),
.C(n_34),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_49),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_66),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_14),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_42),
.B1(n_14),
.B2(n_15),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_25),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_16),
.C(n_18),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2x1_ASAP7_75t_SL g72 ( 
.A(n_61),
.B(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_72),
.B(n_75),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_64),
.A2(n_57),
.B(n_58),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_73),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_67),
.B(n_68),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_0),
.B(n_3),
.Y(n_86)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_81),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_71),
.C(n_16),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_83),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_71),
.C(n_25),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_18),
.C(n_2),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_86),
.B1(n_78),
.B2(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_87),
.B(n_88),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_4),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_90),
.A2(n_91),
.B(n_5),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_92),
.A2(n_93),
.B(n_5),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_6),
.Y(n_95)
);


endmodule