module fake_jpeg_22199_n_220 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_220);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_19),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_59),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_29),
.B1(n_17),
.B2(n_34),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_57),
.B1(n_21),
.B2(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_61),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_29),
.B1(n_24),
.B2(n_15),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_16),
.B1(n_20),
.B2(n_27),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_32),
.A2(n_29),
.B1(n_17),
.B2(n_26),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_26),
.B1(n_27),
.B2(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_23),
.B1(n_28),
.B2(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_18),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_25),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_67),
.B1(n_71),
.B2(n_80),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_69),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_25),
.B1(n_21),
.B2(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_61),
.B(n_56),
.C(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_77),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_54),
.B1(n_44),
.B2(n_51),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_63),
.B(n_48),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_54),
.B1(n_45),
.B2(n_50),
.Y(n_84)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_79),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_21),
.B(n_25),
.C(n_39),
.Y(n_77)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_44),
.B1(n_49),
.B2(n_45),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_0),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_58),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_87),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_86),
.B1(n_94),
.B2(n_101),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_38),
.B1(n_47),
.B2(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_46),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_50),
.B1(n_60),
.B2(n_21),
.Y(n_94)
);

AND2x4_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_77),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_74),
.C(n_82),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_47),
.Y(n_99)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

OAI32xp33_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_47),
.A3(n_8),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_122)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_103),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_87),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_98),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_118),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_77),
.B(n_67),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_97),
.B(n_85),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_65),
.B1(n_69),
.B2(n_73),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_115),
.B1(n_120),
.B2(n_93),
.Y(n_129)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_103),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_73),
.B1(n_78),
.B2(n_64),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_83),
.B(n_70),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_89),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_95),
.A2(n_70),
.B1(n_78),
.B2(n_75),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_121),
.B1(n_94),
.B2(n_84),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_81),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_124),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_79),
.B1(n_47),
.B2(n_66),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_79),
.B1(n_66),
.B2(n_0),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_102),
.B1(n_101),
.B2(n_100),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_1),
.Y(n_124)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_128),
.Y(n_157)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_129),
.B(n_117),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_106),
.Y(n_150)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_99),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_139),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_138),
.B(n_140),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_104),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_135),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_85),
.C(n_92),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_143),
.C(n_113),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_144),
.B(n_116),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_90),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_142),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_88),
.C(n_86),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_86),
.B(n_1),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_150),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_109),
.B(n_108),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_161),
.B(n_127),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_158),
.Y(n_174)
);

AOI221xp5_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_123),
.B1(n_124),
.B2(n_86),
.C(n_6),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_110),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_90),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_110),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_129),
.C(n_143),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_105),
.B(n_109),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_155),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_162),
.B(n_163),
.Y(n_185)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

OAI22x1_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_141),
.B1(n_109),
.B2(n_144),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_165),
.B1(n_173),
.B2(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

AOI321xp33_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_176),
.A3(n_161),
.B1(n_160),
.B2(n_158),
.C(n_152),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_133),
.A3(n_138),
.B1(n_107),
.B2(n_112),
.C1(n_127),
.C2(n_125),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_170),
.Y(n_177)
);

AOI322xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_107),
.A3(n_105),
.B1(n_123),
.B2(n_119),
.C1(n_140),
.C2(n_135),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_175),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_153),
.A2(n_128),
.B1(n_86),
.B2(n_124),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_90),
.C(n_3),
.Y(n_176)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_154),
.B1(n_153),
.B2(n_147),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_165),
.B1(n_173),
.B2(n_176),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_14),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_159),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_187),
.C(n_188),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_151),
.B1(n_147),
.B2(n_145),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_186),
.A2(n_172),
.B1(n_1),
.B2(n_6),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_175),
.B(n_9),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_192),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_197),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_179),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_194),
.A2(n_195),
.B(n_188),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_181),
.B(n_7),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_185),
.B(n_9),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_203),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_182),
.B(n_177),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_196),
.B(n_189),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_181),
.Y(n_203)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_204),
.B(n_194),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_177),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_12),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_209),
.Y(n_210)
);

OAI321xp33_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_10),
.A3(n_12),
.B1(n_13),
.B2(n_184),
.C(n_202),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_203),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_13),
.Y(n_216)
);

AO21x1_ASAP7_75t_SL g215 ( 
.A1(n_212),
.A2(n_13),
.B(n_213),
.Y(n_215)
);

INVx11_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g218 ( 
.A(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_215),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_218),
.A2(n_216),
.B(n_217),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_216),
.Y(n_220)
);


endmodule