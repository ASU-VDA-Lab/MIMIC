module fake_netlist_1_11066_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
AND2x4_ASAP7_75t_L g3 ( .A(n_0), .B(n_1), .Y(n_3) );
NAND2xp5_ASAP7_75t_SL g4 ( .A(n_2), .B(n_1), .Y(n_4) );
INVx4_ASAP7_75t_L g5 ( .A(n_3), .Y(n_5) );
CKINVDCx5p33_ASAP7_75t_R g6 ( .A(n_3), .Y(n_6) );
OR2x2_ASAP7_75t_L g7 ( .A(n_6), .B(n_0), .Y(n_7) );
NAND3x2_ASAP7_75t_L g8 ( .A(n_7), .B(n_5), .C(n_4), .Y(n_8) );
OAI21xp5_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_5), .B(n_0), .Y(n_9) );
OAI21x1_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_5), .B(n_2), .Y(n_10) );
INVx1_ASAP7_75t_SL g11 ( .A(n_10), .Y(n_11) );
endmodule