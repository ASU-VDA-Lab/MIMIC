module fake_ariane_808_n_769 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_769);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_769;

wire n_295;
wire n_556;
wire n_356;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_187;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_515;
wire n_445;
wire n_379;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_352;
wire n_538;
wire n_206;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_455;
wire n_429;
wire n_365;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_458;
wire n_361;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_203;
wire n_436;
wire n_150;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_147;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_484;
wire n_411;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_79),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_8),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_28),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_18),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVxp67_ASAP7_75t_SL g153 ( 
.A(n_136),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_36),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_102),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_47),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_41),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_98),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_24),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_51),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_74),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_61),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_24),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_56),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_13),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_109),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_52),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_37),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_67),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_23),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_46),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_48),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_70),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_122),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_45),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_12),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_8),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_65),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_141),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_100),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_35),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_53),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_30),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_96),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_76),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_38),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_77),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_6),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_34),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_40),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_105),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_142),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_19),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_0),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_149),
.B(n_0),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_149),
.B(n_1),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_1),
.Y(n_208)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_170),
.Y(n_209)
);

AND2x4_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_146),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_152),
.B(n_2),
.Y(n_211)
);

AND2x4_ASAP7_75t_L g212 ( 
.A(n_156),
.B(n_2),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_147),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_3),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_157),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_153),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_158),
.B(n_3),
.Y(n_219)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_159),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_165),
.B(n_4),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g226 ( 
.A(n_164),
.B(n_4),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_166),
.B(n_5),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_161),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

BUFx8_ASAP7_75t_SL g231 ( 
.A(n_169),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_176),
.B(n_5),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_6),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_210),
.A2(n_177),
.B1(n_197),
.B2(n_179),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_173),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_227),
.A2(n_151),
.B1(n_194),
.B2(n_193),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_210),
.A2(n_196),
.B1(n_194),
.B2(n_193),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_144),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_198),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_199),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_144),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_216),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_210),
.A2(n_196),
.B1(n_189),
.B2(n_186),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_L g250 ( 
.A1(n_228),
.A2(n_189),
.B1(n_186),
.B2(n_185),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_199),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_210),
.A2(n_185),
.B1(n_184),
.B2(n_182),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_210),
.A2(n_184),
.B1(n_182),
.B2(n_181),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

AO22x2_ASAP7_75t_L g255 ( 
.A1(n_208),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_198),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_214),
.B(n_148),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_148),
.Y(n_259)
);

AND2x4_ASAP7_75t_L g260 ( 
.A(n_214),
.B(n_150),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_181),
.B1(n_155),
.B2(n_150),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_198),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_222),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_219),
.A2(n_155),
.B1(n_178),
.B2(n_175),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_208),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_208),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_214),
.B(n_11),
.Y(n_267)
);

OA22x2_ASAP7_75t_L g268 ( 
.A1(n_213),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_198),
.Y(n_269)
);

AND2x6_ASAP7_75t_L g270 ( 
.A(n_212),
.B(n_26),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_L g271 ( 
.A1(n_215),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_205),
.B(n_17),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_205),
.B(n_17),
.Y(n_273)
);

AO22x2_ASAP7_75t_L g274 ( 
.A1(n_215),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_L g275 ( 
.A1(n_215),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_211),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_216),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_L g278 ( 
.A1(n_219),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_278)
);

BUFx6f_ASAP7_75t_SL g279 ( 
.A(n_235),
.Y(n_279)
);

AO22x2_ASAP7_75t_L g280 ( 
.A1(n_212),
.A2(n_25),
.B1(n_31),
.B2(n_32),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_L g281 ( 
.A1(n_201),
.A2(n_209),
.B1(n_229),
.B2(n_233),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_198),
.Y(n_282)
);

AO22x2_ASAP7_75t_L g283 ( 
.A1(n_212),
.A2(n_33),
.B1(n_39),
.B2(n_42),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_230),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_254),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_263),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_229),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_248),
.B(n_216),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_248),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_245),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_239),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_249),
.B(n_209),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_253),
.B(n_209),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_242),
.B(n_233),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_201),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_246),
.B(n_235),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_251),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_269),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_272),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_257),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_238),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_260),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_282),
.Y(n_306)
);

INVx4_ASAP7_75t_SL g307 ( 
.A(n_270),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_269),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_267),
.Y(n_309)
);

NAND2x1p5_ASAP7_75t_L g310 ( 
.A(n_265),
.B(n_212),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_244),
.A2(n_212),
.B(n_232),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_243),
.B(n_209),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_281),
.B(n_217),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_279),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_279),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_255),
.B(n_274),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g317 ( 
.A(n_270),
.B(n_201),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_240),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_281),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_277),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_270),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_270),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_283),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_247),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_258),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_259),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_252),
.B(n_209),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_283),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_241),
.B(n_209),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_283),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_280),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_280),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_264),
.B(n_209),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_280),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_268),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_268),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_255),
.B(n_226),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_266),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_255),
.B(n_235),
.Y(n_339)
);

NAND2x1p5_ASAP7_75t_L g340 ( 
.A(n_274),
.B(n_226),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_250),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_274),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_276),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_250),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_278),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_261),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_261),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_271),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_296),
.B(n_271),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_223),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_345),
.A2(n_226),
.B1(n_232),
.B2(n_275),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_318),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_298),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_223),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_321),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_291),
.Y(n_357)
);

OR2x6_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_226),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_336),
.B(n_223),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_291),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_321),
.Y(n_361)
);

NAND2x1p5_ASAP7_75t_L g362 ( 
.A(n_322),
.B(n_226),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_300),
.B(n_232),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_319),
.B(n_204),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_324),
.B(n_209),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_285),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_340),
.B(n_275),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_286),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_320),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_204),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_301),
.B(n_232),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_322),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_287),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_345),
.B(n_232),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_295),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_311),
.A2(n_326),
.B(n_325),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_302),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_290),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_309),
.B(n_204),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_296),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_303),
.B(n_218),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_297),
.B(n_211),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_308),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_290),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_296),
.B(n_218),
.Y(n_385)
);

NAND2x1p5_ASAP7_75t_L g386 ( 
.A(n_317),
.B(n_236),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_317),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_292),
.A2(n_202),
.B(n_278),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_304),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_317),
.B(n_236),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_339),
.B(n_230),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_340),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_295),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_306),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_288),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_308),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_288),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_337),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_313),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_297),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_346),
.B(n_230),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_346),
.B(n_234),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_337),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_347),
.B(n_234),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_305),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_307),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_341),
.B(n_348),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_344),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_303),
.B(n_338),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_293),
.B(n_236),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_342),
.B(n_234),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_305),
.B(n_213),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_307),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_344),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_294),
.B(n_236),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_307),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_409),
.B(n_343),
.Y(n_417)
);

OR2x6_ASAP7_75t_L g418 ( 
.A(n_392),
.B(n_310),
.Y(n_418)
);

NAND2x1_ASAP7_75t_SL g419 ( 
.A(n_378),
.B(n_331),
.Y(n_419)
);

CKINVDCx6p67_ASAP7_75t_R g420 ( 
.A(n_369),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_387),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_409),
.Y(n_422)
);

NOR2x1_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_332),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_380),
.B(n_314),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_343),
.Y(n_425)
);

AND2x2_ASAP7_75t_SL g426 ( 
.A(n_367),
.B(n_328),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_380),
.B(n_315),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_384),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_352),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_407),
.B(n_307),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_377),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_401),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_381),
.B(n_367),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_401),
.B(n_310),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_402),
.Y(n_435)
);

NAND2x1_ASAP7_75t_L g436 ( 
.A(n_358),
.B(n_334),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_355),
.B(n_316),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_349),
.B(n_316),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_413),
.Y(n_439)
);

BUFx5_ASAP7_75t_L g440 ( 
.A(n_406),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_387),
.B(n_334),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_395),
.B(n_310),
.Y(n_442)
);

BUFx6f_ASAP7_75t_SL g443 ( 
.A(n_358),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_391),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_402),
.B(n_224),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_386),
.Y(n_446)
);

INVx6_ASAP7_75t_L g447 ( 
.A(n_404),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_391),
.B(n_328),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_405),
.B(n_323),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_408),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_377),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_414),
.B(n_329),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_412),
.B(n_323),
.Y(n_453)
);

AND2x2_ASAP7_75t_SL g454 ( 
.A(n_351),
.B(n_312),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_412),
.B(n_224),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_377),
.Y(n_456)
);

NOR2x1_ASAP7_75t_L g457 ( 
.A(n_416),
.B(n_313),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_398),
.B(n_327),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_405),
.B(n_330),
.Y(n_459)
);

OR2x6_ASAP7_75t_L g460 ( 
.A(n_358),
.B(n_330),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_375),
.B(n_333),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_386),
.Y(n_463)
);

CKINVDCx8_ASAP7_75t_R g464 ( 
.A(n_358),
.Y(n_464)
);

CKINVDCx6p67_ASAP7_75t_R g465 ( 
.A(n_358),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_404),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_370),
.B(n_299),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_403),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_375),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_357),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_393),
.B(n_205),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_386),
.Y(n_472)
);

CKINVDCx8_ASAP7_75t_R g473 ( 
.A(n_351),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_429),
.Y(n_474)
);

BUFx4f_ASAP7_75t_L g475 ( 
.A(n_420),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_425),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_464),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_433),
.A2(n_385),
.B1(n_370),
.B2(n_399),
.Y(n_478)
);

BUFx12f_ASAP7_75t_L g479 ( 
.A(n_428),
.Y(n_479)
);

NAND2x1p5_ASAP7_75t_L g480 ( 
.A(n_430),
.B(n_399),
.Y(n_480)
);

BUFx4_ASAP7_75t_SL g481 ( 
.A(n_450),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_448),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_470),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_447),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_446),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_446),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_422),
.Y(n_487)
);

BUFx2_ASAP7_75t_SL g488 ( 
.A(n_443),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_417),
.B(n_422),
.Y(n_489)
);

INVx5_ASAP7_75t_L g490 ( 
.A(n_460),
.Y(n_490)
);

BUFx2_ASAP7_75t_SL g491 ( 
.A(n_443),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_468),
.Y(n_492)
);

INVx5_ASAP7_75t_L g493 ( 
.A(n_460),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_446),
.Y(n_494)
);

INVx3_ASAP7_75t_SL g495 ( 
.A(n_465),
.Y(n_495)
);

INVx5_ASAP7_75t_SL g496 ( 
.A(n_460),
.Y(n_496)
);

NAND2x1p5_ASAP7_75t_L g497 ( 
.A(n_430),
.B(n_416),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_447),
.Y(n_498)
);

OR2x6_ASAP7_75t_L g499 ( 
.A(n_418),
.B(n_393),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_458),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_469),
.Y(n_501)
);

BUFx4_ASAP7_75t_SL g502 ( 
.A(n_418),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_461),
.Y(n_503)
);

OAI22xp33_ASAP7_75t_L g504 ( 
.A1(n_473),
.A2(n_397),
.B1(n_388),
.B2(n_400),
.Y(n_504)
);

BUFx2_ASAP7_75t_SL g505 ( 
.A(n_424),
.Y(n_505)
);

INVx5_ASAP7_75t_L g506 ( 
.A(n_418),
.Y(n_506)
);

CKINVDCx8_ASAP7_75t_R g507 ( 
.A(n_461),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_419),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_463),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_449),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_466),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_452),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_424),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_421),
.Y(n_514)
);

NOR2xp67_ASAP7_75t_L g515 ( 
.A(n_438),
.B(n_382),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_427),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_427),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_454),
.A2(n_397),
.B1(n_218),
.B2(n_221),
.Y(n_518)
);

OAI22x1_ASAP7_75t_L g519 ( 
.A1(n_518),
.A2(n_437),
.B1(n_442),
.B2(n_435),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_504),
.A2(n_388),
.B1(n_426),
.B2(n_455),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_515),
.A2(n_432),
.B1(n_434),
.B2(n_421),
.Y(n_521)
);

NAND2x1p5_ASAP7_75t_L g522 ( 
.A(n_506),
.B(n_472),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_512),
.A2(n_445),
.B1(n_472),
.B2(n_444),
.Y(n_523)
);

BUFx12f_ASAP7_75t_L g524 ( 
.A(n_479),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_474),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_492),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_504),
.A2(n_441),
.B1(n_353),
.B2(n_366),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_476),
.A2(n_441),
.B1(n_353),
.B2(n_366),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_483),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_481),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_483),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_499),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_479),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_478),
.A2(n_237),
.B(n_202),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_476),
.A2(n_512),
.B1(n_489),
.B2(n_500),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_511),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_487),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_482),
.A2(n_368),
.B1(n_373),
.B2(n_400),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_475),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_503),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_490),
.Y(n_541)
);

INVx6_ASAP7_75t_L g542 ( 
.A(n_501),
.Y(n_542)
);

BUFx10_ASAP7_75t_L g543 ( 
.A(n_484),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_513),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_510),
.Y(n_545)
);

OAI22xp33_ASAP7_75t_L g546 ( 
.A1(n_507),
.A2(n_467),
.B1(n_453),
.B2(n_374),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_510),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_482),
.A2(n_376),
.B(n_390),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_501),
.Y(n_549)
);

INVx5_ASAP7_75t_L g550 ( 
.A(n_499),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_490),
.B(n_431),
.Y(n_551)
);

INVx6_ASAP7_75t_L g552 ( 
.A(n_490),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_505),
.A2(n_368),
.B1(n_373),
.B2(n_471),
.Y(n_553)
);

INVx6_ASAP7_75t_L g554 ( 
.A(n_490),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g555 ( 
.A(n_487),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_499),
.A2(n_471),
.B1(n_462),
.B2(n_431),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_477),
.A2(n_237),
.B(n_364),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_507),
.A2(n_376),
.B1(n_374),
.B2(n_363),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_516),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_520),
.A2(n_517),
.B1(n_516),
.B2(n_514),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_529),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_542),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_520),
.A2(n_449),
.B1(n_459),
.B2(n_517),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_531),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_541),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_519),
.A2(n_506),
.B1(n_477),
.B2(n_508),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_527),
.B(n_451),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_546),
.A2(n_506),
.B1(n_456),
.B2(n_462),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_548),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_558),
.A2(n_506),
.B1(n_488),
.B2(n_491),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_551),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_548),
.B(n_451),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_523),
.A2(n_456),
.B1(n_365),
.B2(n_394),
.Y(n_573)
);

BUFx4f_ASAP7_75t_SL g574 ( 
.A(n_524),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_521),
.A2(n_394),
.B1(n_389),
.B2(n_498),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_551),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_545),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_538),
.A2(n_389),
.B1(n_394),
.B2(n_457),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_558),
.A2(n_496),
.B1(n_493),
.B2(n_509),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_540),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_528),
.A2(n_457),
.B1(n_423),
.B2(n_509),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_SL g582 ( 
.A1(n_532),
.A2(n_496),
.B1(n_493),
.B2(n_410),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_547),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_SL g584 ( 
.A1(n_532),
.A2(n_496),
.B1(n_493),
.B2(n_410),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_559),
.A2(n_423),
.B1(n_221),
.B2(n_364),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_535),
.A2(n_495),
.B1(n_481),
.B2(n_493),
.Y(n_586)
);

AOI222xp33_ASAP7_75t_L g587 ( 
.A1(n_534),
.A2(n_354),
.B1(n_350),
.B2(n_359),
.C1(n_411),
.C2(n_205),
.Y(n_587)
);

OAI22xp33_ASAP7_75t_L g588 ( 
.A1(n_557),
.A2(n_495),
.B1(n_475),
.B2(n_436),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_526),
.A2(n_544),
.B1(n_532),
.B2(n_550),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_534),
.A2(n_390),
.B1(n_371),
.B2(n_363),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_532),
.A2(n_221),
.B1(n_411),
.B2(n_480),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_525),
.Y(n_592)
);

OAI21xp33_ASAP7_75t_L g593 ( 
.A1(n_557),
.A2(n_371),
.B(n_415),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_541),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_550),
.A2(n_480),
.B1(n_372),
.B2(n_360),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_550),
.A2(n_372),
.B1(n_360),
.B2(n_357),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_555),
.B(n_485),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_550),
.A2(n_372),
.B1(n_360),
.B2(n_357),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_537),
.B(n_485),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_536),
.A2(n_556),
.B1(n_553),
.B2(n_537),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_537),
.A2(n_372),
.B1(n_415),
.B2(n_459),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_522),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_542),
.B(n_485),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g604 ( 
.A(n_539),
.B(n_502),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_539),
.A2(n_379),
.B1(n_497),
.B2(n_383),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_522),
.B(n_485),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_549),
.A2(n_439),
.B1(n_396),
.B2(n_497),
.Y(n_607)
);

OAI221xp5_ASAP7_75t_SL g608 ( 
.A1(n_593),
.A2(n_379),
.B1(n_359),
.B2(n_354),
.C(n_350),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_SL g609 ( 
.A1(n_567),
.A2(n_554),
.B1(n_552),
.B2(n_533),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_563),
.A2(n_533),
.B1(n_530),
.B2(n_549),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_566),
.A2(n_554),
.B1(n_552),
.B2(n_439),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_563),
.A2(n_383),
.B1(n_362),
.B2(n_494),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_567),
.A2(n_206),
.B1(n_396),
.B2(n_198),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_569),
.B(n_486),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_568),
.A2(n_206),
.B1(n_396),
.B2(n_198),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_SL g616 ( 
.A1(n_586),
.A2(n_502),
.B1(n_494),
.B2(n_486),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_604),
.A2(n_494),
.B1(n_486),
.B2(n_383),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_585),
.A2(n_206),
.B1(n_203),
.B2(n_200),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_580),
.B(n_486),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_592),
.B(n_571),
.Y(n_620)
);

NAND3xp33_ASAP7_75t_L g621 ( 
.A(n_593),
.B(n_200),
.C(n_203),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_570),
.A2(n_383),
.B1(n_362),
.B2(n_494),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_573),
.A2(n_200),
.B1(n_203),
.B2(n_440),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_SL g624 ( 
.A1(n_605),
.A2(n_543),
.B1(n_200),
.B2(n_203),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_587),
.A2(n_560),
.B1(n_564),
.B2(n_600),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_588),
.A2(n_362),
.B1(n_361),
.B2(n_356),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_564),
.A2(n_200),
.B1(n_203),
.B2(n_440),
.Y(n_627)
);

OAI221xp5_ASAP7_75t_SL g628 ( 
.A1(n_579),
.A2(n_543),
.B1(n_217),
.B2(n_413),
.C(n_203),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g629 ( 
.A(n_562),
.Y(n_629)
);

OAI221xp5_ASAP7_75t_L g630 ( 
.A1(n_591),
.A2(n_217),
.B1(n_200),
.B2(n_203),
.C(n_207),
.Y(n_630)
);

NAND3xp33_ASAP7_75t_L g631 ( 
.A(n_577),
.B(n_200),
.C(n_217),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_571),
.B(n_576),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_590),
.A2(n_217),
.B1(n_413),
.B2(n_207),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_575),
.A2(n_217),
.B1(n_207),
.B2(n_220),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_576),
.A2(n_440),
.B1(n_207),
.B2(n_217),
.Y(n_635)
);

NOR2xp67_ASAP7_75t_L g636 ( 
.A(n_565),
.B(n_43),
.Y(n_636)
);

AOI221xp5_ASAP7_75t_L g637 ( 
.A1(n_577),
.A2(n_217),
.B1(n_207),
.B2(n_225),
.C(n_220),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_572),
.B(n_440),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_561),
.A2(n_440),
.B1(n_207),
.B2(n_220),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_SL g640 ( 
.A1(n_569),
.A2(n_572),
.B1(n_561),
.B2(n_602),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_581),
.A2(n_207),
.B1(n_225),
.B2(n_220),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_583),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_583),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_602),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_620),
.B(n_562),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_642),
.B(n_565),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_SL g647 ( 
.A1(n_616),
.A2(n_589),
.B(n_574),
.Y(n_647)
);

OAI21xp33_ASAP7_75t_L g648 ( 
.A1(n_608),
.A2(n_597),
.B(n_594),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_642),
.B(n_565),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_643),
.B(n_594),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_643),
.B(n_594),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_619),
.B(n_603),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_614),
.B(n_606),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_614),
.B(n_606),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_638),
.B(n_599),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_629),
.B(n_578),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_640),
.B(n_582),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_632),
.B(n_607),
.Y(n_658)
);

OA211x2_ASAP7_75t_L g659 ( 
.A1(n_621),
.A2(n_625),
.B(n_611),
.C(n_613),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_612),
.A2(n_601),
.B1(n_598),
.B2(n_596),
.Y(n_660)
);

NAND3xp33_ASAP7_75t_L g661 ( 
.A(n_610),
.B(n_595),
.C(n_584),
.Y(n_661)
);

NAND3xp33_ASAP7_75t_L g662 ( 
.A(n_622),
.B(n_220),
.C(n_225),
.Y(n_662)
);

OAI221xp5_ASAP7_75t_SL g663 ( 
.A1(n_624),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.C(n_54),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_644),
.B(n_55),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_644),
.B(n_57),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_626),
.B(n_58),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_SL g667 ( 
.A1(n_609),
.A2(n_59),
.B(n_60),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_636),
.A2(n_225),
.B(n_220),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_636),
.B(n_62),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_617),
.B(n_63),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_633),
.B(n_64),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_631),
.B(n_66),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_653),
.B(n_627),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_SL g674 ( 
.A1(n_657),
.A2(n_630),
.B1(n_634),
.B2(n_628),
.Y(n_674)
);

AOI221xp5_ASAP7_75t_L g675 ( 
.A1(n_648),
.A2(n_623),
.B1(n_618),
.B2(n_615),
.C(n_641),
.Y(n_675)
);

NOR3xp33_ASAP7_75t_L g676 ( 
.A(n_667),
.B(n_637),
.C(n_639),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_653),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_655),
.B(n_635),
.Y(n_678)
);

NOR3xp33_ASAP7_75t_L g679 ( 
.A(n_647),
.B(n_68),
.C(n_69),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_649),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_648),
.A2(n_225),
.B1(n_220),
.B2(n_73),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_654),
.B(n_71),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_659),
.A2(n_657),
.B1(n_661),
.B2(n_666),
.Y(n_683)
);

NAND4xp75_ASAP7_75t_L g684 ( 
.A(n_659),
.B(n_658),
.C(n_656),
.D(n_652),
.Y(n_684)
);

NOR3xp33_ASAP7_75t_L g685 ( 
.A(n_661),
.B(n_72),
.C(n_75),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_L g686 ( 
.A(n_645),
.B(n_225),
.C(n_81),
.Y(n_686)
);

NAND4xp75_ASAP7_75t_L g687 ( 
.A(n_671),
.B(n_78),
.C(n_82),
.D(n_83),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_655),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_671),
.A2(n_225),
.B1(n_85),
.B2(n_86),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_654),
.B(n_84),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_680),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_688),
.Y(n_692)
);

CKINVDCx16_ASAP7_75t_R g693 ( 
.A(n_683),
.Y(n_693)
);

NAND4xp25_ASAP7_75t_SL g694 ( 
.A(n_679),
.B(n_662),
.C(n_650),
.D(n_651),
.Y(n_694)
);

NAND4xp75_ASAP7_75t_L g695 ( 
.A(n_689),
.B(n_670),
.C(n_665),
.D(n_669),
.Y(n_695)
);

XNOR2xp5_ASAP7_75t_L g696 ( 
.A(n_684),
.B(n_646),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_677),
.B(n_646),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_673),
.B(n_650),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_690),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_678),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_678),
.B(n_651),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_698),
.B(n_682),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_691),
.Y(n_703)
);

XOR2x2_ASAP7_75t_L g704 ( 
.A(n_696),
.B(n_681),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_691),
.Y(n_705)
);

XOR2x2_ASAP7_75t_L g706 ( 
.A(n_696),
.B(n_681),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_702),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_704),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_703),
.Y(n_709)
);

OA22x2_ASAP7_75t_L g710 ( 
.A1(n_704),
.A2(n_700),
.B1(n_698),
.B2(n_701),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_706),
.A2(n_693),
.B1(n_695),
.B2(n_699),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_709),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_707),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_708),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_707),
.Y(n_715)
);

OAI322xp33_ASAP7_75t_L g716 ( 
.A1(n_714),
.A2(n_710),
.A3(n_711),
.B1(n_712),
.B2(n_715),
.C1(n_713),
.C2(n_706),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_714),
.A2(n_695),
.B1(n_694),
.B2(n_685),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_712),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_718),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_716),
.A2(n_674),
.B1(n_676),
.B2(n_686),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_717),
.A2(n_692),
.B1(n_699),
.B2(n_705),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_717),
.A2(n_692),
.B1(n_697),
.B2(n_687),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_722),
.A2(n_720),
.B1(n_721),
.B2(n_719),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_SL g724 ( 
.A(n_722),
.B(n_663),
.Y(n_724)
);

OA22x2_ASAP7_75t_L g725 ( 
.A1(n_721),
.A2(n_665),
.B1(n_664),
.B2(n_668),
.Y(n_725)
);

AO22x2_ASAP7_75t_L g726 ( 
.A1(n_719),
.A2(n_662),
.B1(n_697),
.B2(n_672),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_719),
.Y(n_727)
);

NOR2x1_ASAP7_75t_L g728 ( 
.A(n_719),
.B(n_87),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_719),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_728),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_724),
.A2(n_675),
.B1(n_660),
.B2(n_90),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_727),
.Y(n_732)
);

INVxp67_ASAP7_75t_SL g733 ( 
.A(n_729),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_725),
.A2(n_675),
.B1(n_89),
.B2(n_91),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_726),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_723),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_724),
.A2(n_88),
.B1(n_92),
.B2(n_93),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_733),
.B(n_94),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_735),
.Y(n_739)
);

NOR2x1_ASAP7_75t_L g740 ( 
.A(n_732),
.B(n_95),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_730),
.Y(n_741)
);

NAND4xp25_ASAP7_75t_L g742 ( 
.A(n_731),
.B(n_97),
.C(n_99),
.D(n_101),
.Y(n_742)
);

OAI22xp33_ASAP7_75t_L g743 ( 
.A1(n_737),
.A2(n_104),
.B1(n_106),
.B2(n_108),
.Y(n_743)
);

AND4x1_ASAP7_75t_L g744 ( 
.A(n_734),
.B(n_110),
.C(n_111),
.D(n_112),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_736),
.Y(n_745)
);

OR3x2_ASAP7_75t_L g746 ( 
.A(n_741),
.B(n_739),
.C(n_742),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_740),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_745),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_738),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_744),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_743),
.B(n_113),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_745),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_752),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_748),
.Y(n_754)
);

NAND4xp25_ASAP7_75t_L g755 ( 
.A(n_749),
.B(n_115),
.C(n_117),
.D(n_119),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_747),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_746),
.A2(n_750),
.B1(n_751),
.B2(n_127),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_751),
.A2(n_124),
.B1(n_126),
.B2(n_129),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_753),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_754),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_757),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_755),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_761),
.A2(n_758),
.B1(n_756),
.B2(n_132),
.Y(n_763)
);

OA22x2_ASAP7_75t_L g764 ( 
.A1(n_760),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_764),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_765),
.A2(n_759),
.B1(n_762),
.B2(n_763),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_766),
.Y(n_767)
);

AOI221xp5_ASAP7_75t_L g768 ( 
.A1(n_767),
.A2(n_759),
.B1(n_135),
.B2(n_137),
.C(n_138),
.Y(n_768)
);

AOI211xp5_ASAP7_75t_L g769 ( 
.A1(n_768),
.A2(n_134),
.B(n_139),
.C(n_140),
.Y(n_769)
);


endmodule