module fake_netlist_5_2251_n_109 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_109);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_109;

wire n_91;
wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_96;
wire n_37;
wire n_108;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_94;
wire n_38;
wire n_105;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_99;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVxp67_ASAP7_75t_SL g22 ( 
.A(n_19),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_21),
.A2(n_27),
.B1(n_30),
.B2(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_SL g47 ( 
.A(n_35),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_43),
.B(n_27),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_29),
.Y(n_52)
);

OAI221xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_33),
.B1(n_20),
.B2(n_26),
.C(n_22),
.Y(n_53)
);

OAI221xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_33),
.B1(n_20),
.B2(n_26),
.C(n_22),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_31),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_21),
.B1(n_28),
.B2(n_25),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_46),
.B1(n_47),
.B2(n_25),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_44),
.B1(n_42),
.B2(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_44),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_55),
.B(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_42),
.B1(n_41),
.B2(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_51),
.Y(n_64)
);

AND2x4_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_51),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_62),
.B(n_58),
.C(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_55),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_56),
.B1(n_2),
.B2(n_4),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_49),
.B(n_39),
.C(n_38),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_39),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_13),
.Y(n_72)
);

OR2x6_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_39),
.Y(n_73)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_74)
);

NOR2x1p5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

AND2x4_ASAP7_75t_SL g77 ( 
.A(n_72),
.B(n_39),
.Y(n_77)
);

AND2x6_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_70),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_74),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_78),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_74),
.Y(n_85)
);

OR2x6_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_73),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_83),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_74),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_87),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_78),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_85),
.C(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_86),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_86),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_86),
.C(n_73),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_96),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_97),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_104)
);

AOI211xp5_ASAP7_75t_SL g105 ( 
.A1(n_103),
.A2(n_100),
.B(n_101),
.C(n_102),
.Y(n_105)
);

NAND5xp2_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_104),
.C(n_103),
.D(n_11),
.E(n_5),
.Y(n_106)
);

OAI222xp33_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_86),
.B1(n_73),
.B2(n_10),
.C1(n_5),
.C2(n_71),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

AOI221xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_38),
.B1(n_71),
.B2(n_78),
.C(n_73),
.Y(n_109)
);


endmodule