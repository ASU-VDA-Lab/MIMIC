module fake_netlist_5_1522_n_2408 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2408);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2408;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_544;
wire n_1007;
wire n_2369;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_2323;
wire n_2203;
wire n_1243;
wire n_1016;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_227;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_2384;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_344;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1587;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_561;
wire n_1319;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_604;
wire n_314;
wire n_368;
wire n_433;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_2339;
wire n_2093;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_2359;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_2346;
wire n_662;
wire n_459;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2399;
wire n_473;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_2400;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1205;
wire n_1044;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_2405;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_2266;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_2333;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_378;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_302;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_321;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_2269;
wire n_2309;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1400;
wire n_1342;
wire n_1214;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1422;
wire n_1077;
wire n_2364;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_323;
wire n_2287;
wire n_356;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_2282;
wire n_510;
wire n_2371;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1543;
wire n_1399;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_2286;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_2363;
wire n_916;
wire n_1081;
wire n_493;
wire n_2332;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_377;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_386;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_328;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_2278;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_2273;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_1138;
wire n_364;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;
wire n_2268;

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_135),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_66),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_128),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_3),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_85),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_27),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_31),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_9),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_58),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_132),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_176),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_221),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_74),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_155),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_187),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_138),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_217),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_45),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_170),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_19),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_210),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_86),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_41),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_102),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_122),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_29),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_220),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_41),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_100),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_72),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_87),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_180),
.Y(n_257)
);

BUFx2_ASAP7_75t_R g258 ( 
.A(n_100),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_216),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_72),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_69),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_87),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_64),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_134),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_222),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_81),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_47),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_22),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_179),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_60),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_60),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_153),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_73),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_147),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_81),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_34),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_90),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_125),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_130),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_171),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_203),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_219),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_69),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_66),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_62),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_186),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_177),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_139),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_0),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_42),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_13),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_24),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_205),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_213),
.Y(n_294)
);

BUFx8_ASAP7_75t_SL g295 ( 
.A(n_169),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_137),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_136),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_6),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_144),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_27),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_206),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_115),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_223),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_49),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_71),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_54),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_22),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_145),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_191),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_107),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_40),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_218),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_141),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_211),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_93),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_83),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_104),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_88),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_114),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_35),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_109),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_127),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_91),
.Y(n_323)
);

BUFx10_ASAP7_75t_L g324 ( 
.A(n_45),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_149),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_25),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_204),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_5),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_21),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_89),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_112),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_151),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_17),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_24),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_162),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_123),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_202),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_94),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_30),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_34),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_93),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_3),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_10),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_98),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_188),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_157),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_85),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_111),
.Y(n_348)
);

BUFx8_ASAP7_75t_SL g349 ( 
.A(n_174),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_42),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_29),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_95),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_2),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_26),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g355 ( 
.A(n_5),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_32),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_126),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_21),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_61),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_51),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_212),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_46),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_71),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_6),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_1),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_195),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_160),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_63),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_91),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_51),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_19),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_101),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_189),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_74),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_97),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_8),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_64),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_63),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_58),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_1),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_33),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_168),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_38),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_117),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_201),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_30),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_164),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_143),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_52),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_167),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_82),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_89),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_86),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_4),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_185),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_207),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_39),
.Y(n_397)
);

BUFx2_ASAP7_75t_SL g398 ( 
.A(n_175),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_2),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_52),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_55),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_116),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_158),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_121),
.Y(n_404)
);

CKINVDCx14_ASAP7_75t_R g405 ( 
.A(n_140),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_18),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_67),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_106),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_62),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_148),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_46),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_96),
.Y(n_412)
);

BUFx10_ASAP7_75t_L g413 ( 
.A(n_119),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_150),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_97),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_18),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_14),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_78),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_154),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_124),
.Y(n_420)
);

BUFx10_ASAP7_75t_L g421 ( 
.A(n_181),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_49),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_84),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_11),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_209),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_13),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_214),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_184),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_4),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_23),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_23),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_82),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_70),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_54),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_192),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_40),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_244),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_295),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_349),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_292),
.Y(n_440)
);

BUFx6f_ASAP7_75t_SL g441 ( 
.A(n_299),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_292),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_292),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_292),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_292),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_346),
.B(n_7),
.Y(n_446)
);

BUFx10_ASAP7_75t_L g447 ( 
.A(n_224),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_292),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_292),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_292),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_241),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_276),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_293),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_225),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_309),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_241),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_317),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_387),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_292),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_292),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_242),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_259),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_253),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_363),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_253),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_405),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_253),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_246),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_253),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_253),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_253),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_226),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_249),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_346),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_252),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_257),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_427),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_226),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_226),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_234),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_R g481 ( 
.A(n_240),
.B(n_103),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_268),
.B(n_7),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_234),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_234),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_229),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_229),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_256),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_280),
.B(n_8),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_256),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_256),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_290),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_240),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_241),
.Y(n_493)
);

INVxp33_ASAP7_75t_SL g494 ( 
.A(n_230),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_294),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_280),
.B(n_237),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_290),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_294),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_313),
.Y(n_499)
);

NOR2xp67_ASAP7_75t_L g500 ( 
.A(n_365),
.B(n_9),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_290),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_265),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_272),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_278),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_268),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_279),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_281),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_276),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_237),
.B(n_10),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_282),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_330),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_233),
.B(n_11),
.Y(n_512)
);

INVxp33_ASAP7_75t_SL g513 ( 
.A(n_231),
.Y(n_513)
);

CKINVDCx16_ASAP7_75t_R g514 ( 
.A(n_416),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_330),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_330),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_286),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_354),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_287),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_354),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_301),
.Y(n_521)
);

INVxp33_ASAP7_75t_SL g522 ( 
.A(n_232),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_302),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_354),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_308),
.Y(n_525)
);

NOR2xp67_ASAP7_75t_L g526 ( 
.A(n_365),
.B(n_12),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_312),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_319),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_321),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_296),
.B(n_297),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_233),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_322),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_268),
.B(n_320),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_359),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_325),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_359),
.Y(n_536)
);

CKINVDCx16_ASAP7_75t_R g537 ( 
.A(n_416),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_359),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_313),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_409),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_409),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_327),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_409),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_320),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_245),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_320),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_331),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_415),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_373),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_245),
.Y(n_550)
);

INVxp33_ASAP7_75t_L g551 ( 
.A(n_248),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_313),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_422),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_463),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_454),
.Y(n_555)
);

OAI21x1_ASAP7_75t_L g556 ( 
.A1(n_459),
.A2(n_402),
.B(n_373),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_463),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_437),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_459),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_549),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_465),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_465),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_451),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_461),
.Y(n_564)
);

CKINVDCx16_ASAP7_75t_R g565 ( 
.A(n_514),
.Y(n_565)
);

INVx5_ASAP7_75t_L g566 ( 
.A(n_549),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_467),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_496),
.B(n_296),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_533),
.B(n_415),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_467),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_468),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_469),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_469),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_453),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_470),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_470),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_471),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_471),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_440),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_473),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_530),
.B(n_297),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_452),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_508),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_492),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_440),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_455),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_442),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_442),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_443),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_533),
.B(n_415),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_475),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_443),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_444),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_R g594 ( 
.A(n_466),
.B(n_332),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_476),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_457),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_502),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_458),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_444),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_503),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_477),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_445),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_504),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_553),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_506),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_482),
.B(n_373),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_445),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_505),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_517),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_448),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_448),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_482),
.B(n_402),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_449),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_449),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_450),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_507),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_521),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_505),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_523),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_510),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_450),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_529),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_460),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_460),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_472),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_495),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_472),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_456),
.Y(n_628)
);

BUFx8_ASAP7_75t_L g629 ( 
.A(n_441),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_498),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_478),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_478),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_479),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_479),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_480),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_514),
.B(n_422),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_537),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_519),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_480),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_483),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_525),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_493),
.B(n_335),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_537),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_483),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_527),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_528),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_569),
.Y(n_647)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_606),
.Y(n_648)
);

INVx4_ASAP7_75t_SL g649 ( 
.A(n_606),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_642),
.B(n_494),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_610),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_560),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_556),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_612),
.A2(n_474),
.B1(n_446),
.B2(n_509),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_608),
.B(n_532),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_563),
.B(n_542),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_560),
.Y(n_657)
);

INVx6_ASAP7_75t_L g658 ( 
.A(n_610),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_585),
.Y(n_659)
);

BUFx10_ASAP7_75t_L g660 ( 
.A(n_555),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_569),
.B(n_539),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_563),
.B(n_547),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_558),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_642),
.B(n_513),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_563),
.B(n_451),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_612),
.B(n_451),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_569),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_585),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_560),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_618),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_588),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_560),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_588),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_590),
.B(n_456),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_612),
.B(n_499),
.Y(n_675)
);

OAI21xp33_ASAP7_75t_SL g676 ( 
.A1(n_568),
.A2(n_488),
.B(n_462),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_612),
.B(n_499),
.Y(n_677)
);

BUFx10_ASAP7_75t_L g678 ( 
.A(n_564),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_608),
.B(n_522),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_592),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_590),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_590),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_568),
.B(n_535),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_628),
.B(n_499),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_646),
.B(n_481),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_560),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_618),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_592),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_599),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_571),
.B(n_447),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_581),
.B(n_552),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_582),
.B(n_464),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_599),
.Y(n_693)
);

INVx4_ASAP7_75t_SL g694 ( 
.A(n_606),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_582),
.B(n_552),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_607),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_574),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_586),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_560),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_607),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_614),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_628),
.B(n_552),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_580),
.B(n_447),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_614),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_615),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_559),
.Y(n_706)
);

INVx6_ASAP7_75t_L g707 ( 
.A(n_610),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_615),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_627),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_559),
.Y(n_710)
);

BUFx10_ASAP7_75t_L g711 ( 
.A(n_591),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_595),
.B(n_447),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_623),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_623),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_627),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_637),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_559),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_624),
.B(n_228),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_559),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_624),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_581),
.B(n_544),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_596),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_627),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_579),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_606),
.B(n_228),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_645),
.B(n_447),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_556),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_598),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_556),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_606),
.B(n_303),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_634),
.B(n_544),
.Y(n_731)
);

AND2x2_ASAP7_75t_SL g732 ( 
.A(n_565),
.B(n_402),
.Y(n_732)
);

INVx6_ASAP7_75t_L g733 ( 
.A(n_610),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_610),
.Y(n_734)
);

OR2x2_ASAP7_75t_L g735 ( 
.A(n_583),
.B(n_546),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_610),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_606),
.B(n_546),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_579),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_606),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_627),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_L g741 ( 
.A(n_594),
.B(n_337),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_579),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_597),
.B(n_438),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_587),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_600),
.B(n_439),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_SL g746 ( 
.A1(n_565),
.A2(n_270),
.B1(n_289),
.B2(n_251),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_559),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_559),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_583),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_587),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_605),
.B(n_441),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_587),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_589),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_589),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_611),
.B(n_548),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_616),
.B(n_299),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_589),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_593),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_601),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_634),
.B(n_227),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_604),
.Y(n_761)
);

INVx4_ASAP7_75t_L g762 ( 
.A(n_613),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_639),
.B(n_548),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_620),
.B(n_441),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_639),
.B(n_484),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_640),
.B(n_227),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_640),
.B(n_484),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_604),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_613),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_611),
.B(n_348),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_627),
.Y(n_771)
);

INVx5_ASAP7_75t_L g772 ( 
.A(n_613),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_636),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_593),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_637),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_613),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_613),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_593),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_627),
.Y(n_779)
);

INVx4_ASAP7_75t_L g780 ( 
.A(n_613),
.Y(n_780)
);

AND2x6_ASAP7_75t_L g781 ( 
.A(n_611),
.B(n_235),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_611),
.B(n_235),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_602),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_621),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_567),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_638),
.B(n_299),
.Y(n_786)
);

BUFx8_ASAP7_75t_SL g787 ( 
.A(n_584),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_567),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_641),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_602),
.B(n_236),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_643),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_643),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_621),
.B(n_357),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_602),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_567),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_570),
.Y(n_796)
);

AO22x2_ASAP7_75t_L g797 ( 
.A1(n_630),
.A2(n_512),
.B1(n_300),
.B2(n_355),
.Y(n_797)
);

INVx4_ASAP7_75t_L g798 ( 
.A(n_621),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_584),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_632),
.B(n_236),
.Y(n_800)
);

AO22x2_ASAP7_75t_L g801 ( 
.A1(n_630),
.A2(n_512),
.B1(n_300),
.B2(n_355),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_554),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_570),
.Y(n_803)
);

AO21x2_ASAP7_75t_L g804 ( 
.A1(n_554),
.A2(n_250),
.B(n_239),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_570),
.Y(n_805)
);

BUFx10_ASAP7_75t_L g806 ( 
.A(n_629),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_739),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_739),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_804),
.A2(n_266),
.B1(n_262),
.B2(n_263),
.Y(n_809)
);

NOR2x1p5_ASAP7_75t_L g810 ( 
.A(n_692),
.B(n_238),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_691),
.B(n_621),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_789),
.Y(n_812)
);

OR2x6_ASAP7_75t_L g813 ( 
.A(n_791),
.B(n_626),
.Y(n_813)
);

INVx5_ASAP7_75t_L g814 ( 
.A(n_653),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_792),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_691),
.B(n_621),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_650),
.B(n_629),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_664),
.B(n_621),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_683),
.B(n_291),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_666),
.B(n_557),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_676),
.A2(n_366),
.B1(n_367),
.B2(n_361),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_732),
.B(n_629),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_667),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_648),
.B(n_629),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_647),
.A2(n_526),
.B(n_500),
.C(n_250),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_667),
.B(n_485),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_695),
.B(n_291),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_695),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_666),
.B(n_557),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_659),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_659),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_732),
.A2(n_382),
.B1(n_384),
.B2(n_372),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_804),
.A2(n_266),
.B1(n_248),
.B2(n_263),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_653),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_804),
.A2(n_782),
.B1(n_721),
.B2(n_790),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_668),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_666),
.B(n_561),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_666),
.B(n_561),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_688),
.B(n_562),
.Y(n_839)
);

INVxp33_ASAP7_75t_L g840 ( 
.A(n_768),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_R g841 ( 
.A(n_789),
.B(n_603),
.Y(n_841)
);

INVx8_ASAP7_75t_L g842 ( 
.A(n_697),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_791),
.B(n_551),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_732),
.A2(n_388),
.B1(n_395),
.B2(n_385),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_749),
.B(n_626),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_688),
.B(n_562),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_668),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_792),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_773),
.B(n_318),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_731),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_708),
.B(n_572),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_708),
.B(n_647),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_681),
.B(n_572),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_675),
.A2(n_577),
.B(n_576),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_681),
.B(n_576),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_731),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_735),
.B(n_318),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_671),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_671),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_682),
.B(n_577),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_735),
.B(n_334),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_782),
.A2(n_262),
.B1(n_283),
.B2(n_275),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_682),
.B(n_721),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_673),
.Y(n_864)
);

AND2x4_ASAP7_75t_SL g865 ( 
.A(n_806),
.B(n_609),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_763),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_654),
.A2(n_264),
.B1(n_269),
.B2(n_239),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_718),
.A2(n_531),
.B(n_545),
.C(n_486),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_673),
.B(n_578),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_680),
.B(n_578),
.Y(n_870)
);

INVxp67_ASAP7_75t_L g871 ( 
.A(n_775),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_692),
.B(n_550),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_680),
.B(n_632),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_674),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_684),
.B(n_243),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_653),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_689),
.B(n_693),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_689),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_749),
.B(n_617),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_761),
.B(n_619),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_693),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_663),
.Y(n_882)
);

OR2x6_ASAP7_75t_L g883 ( 
.A(n_799),
.B(n_398),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_696),
.B(n_632),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_661),
.A2(n_403),
.B1(n_404),
.B2(n_396),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_674),
.Y(n_886)
);

NAND2x1_ASAP7_75t_L g887 ( 
.A(n_653),
.B(n_632),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_677),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_648),
.B(n_653),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_648),
.B(n_408),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_702),
.B(n_247),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_696),
.B(n_633),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_700),
.Y(n_893)
);

NAND2x1p5_ASAP7_75t_L g894 ( 
.A(n_648),
.B(n_264),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_761),
.B(n_622),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_746),
.B(n_679),
.C(n_655),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_768),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_670),
.B(n_254),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_648),
.B(n_410),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_661),
.A2(n_414),
.B1(n_420),
.B2(n_419),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_670),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_648),
.B(n_428),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_SL g903 ( 
.A1(n_716),
.A2(n_328),
.B1(n_333),
.B2(n_306),
.Y(n_903)
);

INVx4_ASAP7_75t_L g904 ( 
.A(n_769),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_700),
.B(n_633),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_701),
.B(n_633),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_725),
.A2(n_288),
.B1(n_310),
.B2(n_274),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_802),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_701),
.B(n_704),
.Y(n_909)
);

INVx5_ASAP7_75t_L g910 ( 
.A(n_727),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_704),
.B(n_633),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_802),
.Y(n_912)
);

NOR2x1p5_ASAP7_75t_L g913 ( 
.A(n_663),
.B(n_255),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_705),
.B(n_644),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_705),
.B(n_644),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_713),
.B(n_644),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_713),
.B(n_714),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_765),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_714),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_720),
.B(n_644),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_720),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_656),
.B(n_260),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_727),
.B(n_729),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_698),
.Y(n_924)
);

AO22x1_ASAP7_75t_L g925 ( 
.A1(n_751),
.A2(n_283),
.B1(n_304),
.B2(n_275),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_662),
.B(n_267),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_764),
.B(n_299),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_785),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_785),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_756),
.B(n_271),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_687),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_727),
.B(n_314),
.Y(n_932)
);

AND2x6_ASAP7_75t_SL g933 ( 
.A(n_743),
.B(n_304),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_727),
.B(n_314),
.Y(n_934)
);

NOR2xp67_ASAP7_75t_L g935 ( 
.A(n_745),
.B(n_105),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_665),
.B(n_575),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_782),
.A2(n_345),
.B(n_425),
.C(n_390),
.Y(n_937)
);

NOR3xp33_ASAP7_75t_L g938 ( 
.A(n_799),
.B(n_277),
.C(n_273),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_727),
.B(n_336),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_729),
.B(n_336),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_786),
.B(n_685),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_770),
.B(n_575),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_730),
.A2(n_398),
.B1(n_345),
.B2(n_390),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_765),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_737),
.A2(n_782),
.B1(n_741),
.B2(n_690),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_784),
.B(n_575),
.Y(n_946)
);

BUFx8_ASAP7_75t_L g947 ( 
.A(n_787),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_784),
.B(n_575),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_703),
.A2(n_435),
.B1(n_425),
.B2(n_362),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_806),
.B(n_413),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_784),
.B(n_729),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_788),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_712),
.B(n_284),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_767),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_698),
.Y(n_955)
);

AND2x6_ASAP7_75t_SL g956 ( 
.A(n_760),
.B(n_305),
.Y(n_956)
);

AO22x1_ASAP7_75t_L g957 ( 
.A1(n_760),
.A2(n_329),
.B1(n_316),
.B2(n_311),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_769),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_729),
.B(n_575),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_726),
.B(n_285),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_760),
.Y(n_961)
);

INVx4_ASAP7_75t_L g962 ( 
.A(n_769),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_729),
.B(n_575),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_706),
.B(n_435),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_706),
.B(n_573),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_760),
.B(n_487),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_706),
.B(n_573),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_710),
.B(n_573),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_806),
.B(n_413),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_710),
.B(n_635),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_788),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_710),
.B(n_717),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_717),
.B(n_635),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_790),
.A2(n_431),
.B1(n_329),
.B2(n_380),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_790),
.A2(n_311),
.B1(n_383),
.B2(n_379),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_795),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_767),
.Y(n_977)
);

OR2x6_ASAP7_75t_L g978 ( 
.A(n_961),
.B(n_766),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_830),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_830),
.Y(n_980)
);

INVx5_ASAP7_75t_L g981 ( 
.A(n_834),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_819),
.B(n_766),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_831),
.Y(n_983)
);

AND3x1_ASAP7_75t_SL g984 ( 
.A(n_810),
.B(n_913),
.C(n_258),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_831),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_848),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_842),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_834),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_819),
.B(n_766),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_841),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_836),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_863),
.B(n_888),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_836),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_834),
.Y(n_994)
);

OAI22xp33_ASAP7_75t_L g995 ( 
.A1(n_852),
.A2(n_755),
.B1(n_759),
.B2(n_722),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_843),
.B(n_797),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_966),
.B(n_649),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_841),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_931),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_812),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_847),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_818),
.B(n_766),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_847),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_835),
.A2(n_800),
.B1(n_790),
.B2(n_781),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_815),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_834),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_858),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_901),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_875),
.B(n_800),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_858),
.Y(n_1010)
);

NAND2xp33_ASAP7_75t_SL g1011 ( 
.A(n_817),
.B(n_728),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_859),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_859),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_840),
.B(n_722),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_864),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_897),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_845),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_875),
.B(n_800),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_891),
.B(n_800),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_842),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_864),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_878),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_891),
.B(n_793),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_878),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_881),
.Y(n_1025)
);

NAND3xp33_ASAP7_75t_SL g1026 ( 
.A(n_903),
.B(n_759),
.C(n_338),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_842),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_876),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_867),
.A2(n_781),
.B1(n_738),
.B2(n_742),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_813),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_918),
.B(n_797),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_944),
.B(n_797),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_881),
.Y(n_1033)
);

NOR3xp33_ASAP7_75t_SL g1034 ( 
.A(n_882),
.B(n_307),
.C(n_298),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_922),
.B(n_724),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_R g1036 ( 
.A(n_924),
.B(n_660),
.Y(n_1036)
);

NAND3xp33_ASAP7_75t_SL g1037 ( 
.A(n_896),
.B(n_323),
.C(n_315),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_922),
.B(n_724),
.Y(n_1038)
);

CKINVDCx14_ASAP7_75t_R g1039 ( 
.A(n_955),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_966),
.B(n_649),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_813),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_947),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_893),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_876),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_876),
.Y(n_1045)
);

OR2x6_ASAP7_75t_SL g1046 ( 
.A(n_872),
.B(n_326),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_893),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_926),
.B(n_738),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_926),
.B(n_908),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_912),
.B(n_742),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_813),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_876),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_807),
.B(n_649),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_879),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_877),
.B(n_909),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_919),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_865),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_828),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_880),
.Y(n_1059)
);

AND2x6_ASAP7_75t_L g1060 ( 
.A(n_807),
.B(n_649),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_874),
.A2(n_750),
.B(n_752),
.C(n_744),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_919),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_917),
.B(n_744),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_921),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_871),
.B(n_660),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_921),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_865),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_835),
.A2(n_801),
.B1(n_797),
.B2(n_719),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_807),
.B(n_694),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_807),
.B(n_694),
.Y(n_1070)
);

AO21x2_ASAP7_75t_L g1071 ( 
.A1(n_932),
.A2(n_715),
.B(n_709),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_928),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_954),
.B(n_801),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_811),
.B(n_750),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_928),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_898),
.B(n_341),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_947),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_816),
.B(n_752),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_929),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_886),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_895),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_850),
.A2(n_781),
.B1(n_801),
.B2(n_754),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_977),
.B(n_753),
.Y(n_1083)
);

INVxp67_ASAP7_75t_SL g1084 ( 
.A(n_923),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_929),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_952),
.Y(n_1086)
);

OR2x6_ASAP7_75t_L g1087 ( 
.A(n_808),
.B(n_801),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_856),
.B(n_753),
.Y(n_1088)
);

INVx1_ASAP7_75t_SL g1089 ( 
.A(n_883),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_883),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_808),
.B(n_694),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_814),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_814),
.Y(n_1093)
);

AO22x1_ASAP7_75t_L g1094 ( 
.A1(n_849),
.A2(n_781),
.B1(n_305),
.B2(n_339),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_866),
.B(n_757),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_952),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_853),
.B(n_757),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_855),
.B(n_758),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_971),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_860),
.B(n_849),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_814),
.B(n_678),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_826),
.Y(n_1102)
);

BUFx12f_ASAP7_75t_L g1103 ( 
.A(n_956),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_823),
.B(n_827),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_827),
.B(n_758),
.Y(n_1105)
);

OR2x4_ASAP7_75t_L g1106 ( 
.A(n_941),
.B(n_316),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_839),
.B(n_774),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_814),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_808),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_808),
.B(n_694),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_910),
.B(n_678),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_971),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_976),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_976),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_930),
.A2(n_778),
.B(n_783),
.C(n_774),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_857),
.B(n_678),
.Y(n_1116)
);

INVx4_ASAP7_75t_L g1117 ( 
.A(n_910),
.Y(n_1117)
);

AOI211xp5_ASAP7_75t_L g1118 ( 
.A1(n_861),
.A2(n_339),
.B(n_344),
.C(n_340),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_820),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_910),
.Y(n_1120)
);

NAND2xp33_ASAP7_75t_SL g1121 ( 
.A(n_822),
.B(n_711),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_829),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_837),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_838),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_933),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_826),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_951),
.Y(n_1127)
);

BUFx10_ASAP7_75t_L g1128 ( 
.A(n_857),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_932),
.A2(n_783),
.B(n_794),
.C(n_778),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_887),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_846),
.B(n_794),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_851),
.B(n_717),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_873),
.Y(n_1133)
);

NOR2x1_ASAP7_75t_L g1134 ( 
.A(n_935),
.B(n_651),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_884),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_883),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_892),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_905),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_910),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_945),
.B(n_709),
.Y(n_1140)
);

INVx4_ASAP7_75t_L g1141 ( 
.A(n_904),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_957),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_825),
.B(n_715),
.Y(n_1143)
);

AND2x6_ASAP7_75t_L g1144 ( 
.A(n_959),
.B(n_652),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_861),
.B(n_711),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_906),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_R g1147 ( 
.A(n_941),
.B(n_711),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_923),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_911),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_930),
.A2(n_719),
.B(n_748),
.C(n_669),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_914),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_915),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_869),
.B(n_719),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_904),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_809),
.B(n_795),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_958),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_870),
.B(n_748),
.Y(n_1157)
);

BUFx4f_ASAP7_75t_L g1158 ( 
.A(n_894),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_925),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_916),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_938),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_920),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_809),
.B(n_748),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_833),
.A2(n_781),
.B1(n_803),
.B2(n_805),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_833),
.B(n_781),
.Y(n_1165)
);

INVxp67_ASAP7_75t_L g1166 ( 
.A(n_953),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_970),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_973),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_965),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1129),
.A2(n_963),
.B(n_939),
.Y(n_1170)
);

AOI211x1_ASAP7_75t_L g1171 ( 
.A1(n_1068),
.A2(n_907),
.B(n_939),
.C(n_934),
.Y(n_1171)
);

AOI21xp33_ASAP7_75t_L g1172 ( 
.A1(n_1116),
.A2(n_960),
.B(n_953),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_986),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1053),
.Y(n_1174)
);

INVx5_ASAP7_75t_L g1175 ( 
.A(n_1092),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1127),
.A2(n_940),
.B(n_934),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1055),
.A2(n_960),
.B(n_949),
.C(n_974),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1049),
.B(n_821),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1127),
.A2(n_940),
.B(n_942),
.Y(n_1179)
);

OA22x2_ASAP7_75t_L g1180 ( 
.A1(n_1087),
.A2(n_258),
.B1(n_844),
.B2(n_832),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_983),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1165),
.A2(n_1163),
.B(n_1018),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1100),
.B(n_885),
.Y(n_1183)
);

AOI21x1_ASAP7_75t_SL g1184 ( 
.A1(n_982),
.A2(n_964),
.B(n_972),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1117),
.A2(n_889),
.B(n_958),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_981),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1074),
.A2(n_1078),
.B(n_1130),
.Y(n_1187)
);

AOI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1002),
.A2(n_899),
.B(n_890),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_992),
.B(n_900),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1130),
.A2(n_936),
.B(n_946),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1104),
.B(n_862),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_989),
.A2(n_889),
.B1(n_862),
.B2(n_943),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1009),
.A2(n_1019),
.B(n_1023),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_981),
.Y(n_1194)
);

INVxp67_ASAP7_75t_L g1195 ( 
.A(n_1008),
.Y(n_1195)
);

INVx6_ASAP7_75t_L g1196 ( 
.A(n_986),
.Y(n_1196)
);

INVx4_ASAP7_75t_L g1197 ( 
.A(n_981),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1166),
.B(n_868),
.Y(n_1198)
);

CKINVDCx8_ASAP7_75t_R g1199 ( 
.A(n_1000),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1105),
.B(n_974),
.Y(n_1200)
);

AO22x2_ASAP7_75t_L g1201 ( 
.A1(n_1026),
.A2(n_927),
.B1(n_969),
.B2(n_950),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1122),
.B(n_975),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1130),
.A2(n_1134),
.B(n_1061),
.Y(n_1203)
);

AOI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1035),
.A2(n_902),
.B(n_890),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_SL g1205 ( 
.A1(n_1004),
.A2(n_854),
.B(n_975),
.Y(n_1205)
);

AOI22x1_ASAP7_75t_L g1206 ( 
.A1(n_1135),
.A2(n_894),
.B1(n_686),
.B2(n_652),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1053),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1134),
.A2(n_948),
.B(n_967),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1117),
.A2(n_962),
.B(n_734),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1004),
.A2(n_962),
.B1(n_824),
.B2(n_902),
.Y(n_1210)
);

AO21x2_ASAP7_75t_L g1211 ( 
.A1(n_1150),
.A2(n_824),
.B(n_968),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1122),
.B(n_781),
.Y(n_1212)
);

NAND2x1p5_ASAP7_75t_L g1213 ( 
.A(n_981),
.B(n_651),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1117),
.A2(n_1120),
.B(n_981),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1123),
.B(n_937),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1132),
.A2(n_669),
.B(n_657),
.Y(n_1216)
);

AOI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1038),
.A2(n_1048),
.B(n_980),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1120),
.A2(n_734),
.B(n_651),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_999),
.Y(n_1219)
);

AO32x2_ASAP7_75t_L g1220 ( 
.A1(n_1106),
.A2(n_777),
.A3(n_734),
.B1(n_736),
.B2(n_762),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1120),
.A2(n_981),
.B(n_1156),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1123),
.A2(n_740),
.B(n_723),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1017),
.B(n_487),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1148),
.B(n_769),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_983),
.A2(n_1012),
.B(n_1003),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1084),
.A2(n_1148),
.B1(n_1124),
.B2(n_1119),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1119),
.B(n_723),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_979),
.Y(n_1228)
);

BUFx12f_ASAP7_75t_L g1229 ( 
.A(n_1042),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1003),
.A2(n_672),
.B(n_657),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1164),
.A2(n_771),
.B(n_740),
.Y(n_1231)
);

AOI211x1_ASAP7_75t_L g1232 ( 
.A1(n_1031),
.A2(n_400),
.B(n_394),
.C(n_383),
.Y(n_1232)
);

NOR4xp25_ASAP7_75t_L g1233 ( 
.A(n_1037),
.B(n_1145),
.C(n_996),
.D(n_1032),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1133),
.B(n_1149),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1133),
.B(n_779),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_999),
.Y(n_1236)
);

NOR2x1_ASAP7_75t_SL g1237 ( 
.A(n_1092),
.B(n_769),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1118),
.A2(n_352),
.B(n_344),
.C(n_351),
.Y(n_1238)
);

OAI21xp33_ASAP7_75t_L g1239 ( 
.A1(n_1065),
.A2(n_343),
.B(n_342),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1012),
.A2(n_686),
.B(n_672),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1115),
.A2(n_699),
.A3(n_779),
.B(n_796),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1148),
.B(n_776),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1013),
.A2(n_699),
.B(n_796),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1000),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1149),
.B(n_803),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1013),
.A2(n_805),
.B(n_490),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1152),
.B(n_747),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1164),
.A2(n_762),
.B(n_736),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1054),
.B(n_261),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1155),
.A2(n_1140),
.B(n_1152),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1128),
.B(n_1054),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1015),
.A2(n_490),
.B(n_489),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1156),
.A2(n_1139),
.B(n_1063),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1148),
.B(n_776),
.Y(n_1254)
);

AOI21x1_ASAP7_75t_SL g1255 ( 
.A1(n_1140),
.A2(n_421),
.B(n_413),
.Y(n_1255)
);

NOR2x1_ASAP7_75t_SL g1256 ( 
.A(n_1092),
.B(n_1093),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1015),
.A2(n_491),
.B(n_489),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1139),
.A2(n_780),
.B(n_777),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1160),
.B(n_747),
.Y(n_1259)
);

AOI21x1_ASAP7_75t_L g1260 ( 
.A1(n_979),
.A2(n_631),
.B(n_625),
.Y(n_1260)
);

AOI21x1_ASAP7_75t_L g1261 ( 
.A1(n_980),
.A2(n_991),
.B(n_985),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1148),
.A2(n_658),
.B1(n_707),
.B2(n_733),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1005),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_985),
.Y(n_1264)
);

INVx4_ASAP7_75t_L g1265 ( 
.A(n_1028),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1005),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1030),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_997),
.B(n_777),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1092),
.A2(n_798),
.B(n_780),
.Y(n_1269)
);

AOI21x1_ASAP7_75t_L g1270 ( 
.A1(n_991),
.A2(n_1001),
.B(n_993),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1092),
.A2(n_798),
.B(n_747),
.Y(n_1271)
);

AND3x2_ASAP7_75t_L g1272 ( 
.A(n_1142),
.B(n_351),
.C(n_340),
.Y(n_1272)
);

AOI31xp67_ASAP7_75t_L g1273 ( 
.A1(n_1140),
.A2(n_625),
.A3(n_631),
.B(n_635),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1053),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1093),
.A2(n_1108),
.B(n_1069),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_993),
.A2(n_352),
.A3(n_368),
.B(n_371),
.Y(n_1276)
);

AO21x1_ASAP7_75t_L g1277 ( 
.A1(n_1140),
.A2(n_371),
.B(n_368),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1093),
.A2(n_747),
.B(n_776),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1021),
.A2(n_497),
.B(n_491),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1021),
.Y(n_1280)
);

O2A1O1Ixp5_ASAP7_75t_L g1281 ( 
.A1(n_1143),
.A2(n_374),
.B(n_379),
.C(n_380),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1093),
.A2(n_747),
.B(n_776),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1160),
.B(n_776),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1022),
.A2(n_501),
.B(n_497),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1030),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1128),
.B(n_347),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1001),
.A2(n_511),
.B(n_501),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1059),
.B(n_261),
.Y(n_1288)
);

NOR2x1_ASAP7_75t_SL g1289 ( 
.A(n_1093),
.B(n_772),
.Y(n_1289)
);

INVxp67_ASAP7_75t_SL g1290 ( 
.A(n_1028),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1162),
.B(n_658),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_997),
.B(n_511),
.Y(n_1292)
);

AO21x1_ASAP7_75t_L g1293 ( 
.A1(n_1011),
.A2(n_394),
.B(n_374),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1022),
.A2(n_516),
.B(n_515),
.Y(n_1294)
);

AO21x1_ASAP7_75t_L g1295 ( 
.A1(n_1143),
.A2(n_411),
.B(n_400),
.Y(n_1295)
);

INVx4_ASAP7_75t_L g1296 ( 
.A(n_1028),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1024),
.A2(n_516),
.B(n_515),
.Y(n_1297)
);

AO31x2_ASAP7_75t_L g1298 ( 
.A1(n_1007),
.A2(n_411),
.A3(n_417),
.B(n_418),
.Y(n_1298)
);

AOI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1007),
.A2(n_631),
.B(n_625),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1024),
.A2(n_520),
.B(n_518),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1128),
.B(n_772),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1059),
.Y(n_1302)
);

NOR2x1_ASAP7_75t_SL g1303 ( 
.A(n_1108),
.B(n_772),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1025),
.A2(n_520),
.B(n_518),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_SL g1305 ( 
.A1(n_1082),
.A2(n_418),
.B(n_417),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1057),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1010),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1025),
.A2(n_534),
.B(n_524),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_997),
.B(n_524),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1010),
.Y(n_1310)
);

AO21x1_ASAP7_75t_L g1311 ( 
.A1(n_1143),
.A2(n_433),
.B(n_436),
.Y(n_1311)
);

AO21x1_ASAP7_75t_L g1312 ( 
.A1(n_1143),
.A2(n_433),
.B(n_436),
.Y(n_1312)
);

NAND2x1p5_ASAP7_75t_L g1313 ( 
.A(n_1053),
.B(n_772),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1056),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_997),
.B(n_534),
.Y(n_1315)
);

AO21x1_ASAP7_75t_L g1316 ( 
.A1(n_1121),
.A2(n_432),
.B(n_431),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1033),
.A2(n_540),
.B(n_536),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1108),
.A2(n_772),
.B(n_566),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1147),
.B(n_772),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1081),
.B(n_536),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1040),
.B(n_538),
.Y(n_1321)
);

OAI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1106),
.A2(n_1087),
.B1(n_1082),
.B2(n_1159),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1033),
.A2(n_540),
.B(n_538),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1081),
.B(n_1076),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1043),
.A2(n_1062),
.B(n_1047),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1108),
.A2(n_1070),
.B(n_1069),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1043),
.A2(n_541),
.B(n_543),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_996),
.B(n_261),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1047),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1162),
.B(n_1135),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1108),
.A2(n_566),
.B(n_707),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_SL g1332 ( 
.A(n_990),
.B(n_413),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1056),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1064),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1186),
.Y(n_1335)
);

INVx6_ASAP7_75t_L g1336 ( 
.A(n_1175),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1250),
.B(n_1031),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1172),
.A2(n_1102),
.B1(n_1080),
.B2(n_978),
.Y(n_1338)
);

AO21x2_ASAP7_75t_L g1339 ( 
.A1(n_1193),
.A2(n_1216),
.B(n_1217),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_SL g1340 ( 
.A1(n_1295),
.A2(n_1066),
.B(n_1062),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1180),
.A2(n_1102),
.B1(n_1080),
.B2(n_1161),
.Y(n_1341)
);

O2A1O1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1177),
.A2(n_995),
.B(n_1118),
.C(n_1076),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1174),
.B(n_1032),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1261),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1244),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1243),
.A2(n_1050),
.B(n_1066),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1243),
.A2(n_1157),
.B(n_1153),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1174),
.B(n_1207),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1180),
.A2(n_1126),
.B1(n_1087),
.B2(n_1136),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1270),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1263),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1182),
.A2(n_1168),
.B(n_1131),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1230),
.A2(n_1064),
.B(n_1167),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1181),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1181),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1280),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1280),
.Y(n_1357)
);

CKINVDCx6p67_ASAP7_75t_R g1358 ( 
.A(n_1229),
.Y(n_1358)
);

INVx1_ASAP7_75t_SL g1359 ( 
.A(n_1266),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1244),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1329),
.Y(n_1361)
);

INVx2_ASAP7_75t_SL g1362 ( 
.A(n_1196),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1186),
.A2(n_1154),
.B(n_1141),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1329),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1230),
.A2(n_1169),
.B(n_1167),
.Y(n_1365)
);

INVx3_ASAP7_75t_SL g1366 ( 
.A(n_1196),
.Y(n_1366)
);

OR2x6_ASAP7_75t_L g1367 ( 
.A(n_1171),
.B(n_978),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1183),
.B(n_1073),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1189),
.B(n_1014),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1175),
.Y(n_1370)
);

AO21x2_ASAP7_75t_L g1371 ( 
.A1(n_1216),
.A2(n_1071),
.B(n_1097),
.Y(n_1371)
);

OAI211xp5_ASAP7_75t_L g1372 ( 
.A1(n_1177),
.A2(n_1051),
.B(n_1041),
.C(n_1016),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1174),
.B(n_1109),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1240),
.A2(n_1169),
.B(n_1168),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1240),
.A2(n_994),
.B(n_988),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1178),
.A2(n_1107),
.B(n_1137),
.Y(n_1376)
);

AO21x2_ASAP7_75t_L g1377 ( 
.A1(n_1187),
.A2(n_1071),
.B(n_1098),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1234),
.A2(n_1191),
.B1(n_1200),
.B2(n_1202),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1195),
.B(n_990),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1225),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_1324),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1207),
.B(n_1109),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1175),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1330),
.B(n_1073),
.Y(n_1384)
);

O2A1O1Ixp5_ASAP7_75t_L g1385 ( 
.A1(n_1178),
.A2(n_1111),
.B(n_1101),
.C(n_1094),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1198),
.B(n_998),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1293),
.A2(n_1087),
.B1(n_1089),
.B2(n_1090),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1246),
.A2(n_994),
.B(n_988),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1207),
.B(n_1155),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1186),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1175),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1219),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1228),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1187),
.A2(n_1088),
.B(n_1083),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1201),
.A2(n_1205),
.B1(n_1322),
.B2(n_1328),
.Y(n_1395)
);

NAND2x1p5_ASAP7_75t_L g1396 ( 
.A(n_1194),
.B(n_1028),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1274),
.B(n_1087),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1190),
.A2(n_1071),
.B(n_1095),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1225),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1320),
.B(n_1137),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1179),
.A2(n_1146),
.B(n_1138),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1192),
.A2(n_1146),
.B(n_1138),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1274),
.B(n_1151),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1194),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1196),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1325),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1190),
.A2(n_1079),
.B(n_1075),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1246),
.A2(n_994),
.B(n_988),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1322),
.A2(n_1106),
.B1(n_984),
.B2(n_998),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1201),
.A2(n_978),
.B1(n_1058),
.B2(n_987),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1325),
.A2(n_1045),
.B(n_1006),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1203),
.A2(n_1045),
.B(n_1006),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1264),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1219),
.Y(n_1414)
);

CKINVDCx16_ASAP7_75t_R g1415 ( 
.A(n_1229),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1307),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1236),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1203),
.A2(n_1045),
.B(n_1006),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1208),
.A2(n_1052),
.B(n_1151),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1208),
.A2(n_1052),
.B(n_1072),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1252),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1286),
.B(n_1094),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1194),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1286),
.B(n_1109),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1252),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1302),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1257),
.Y(n_1427)
);

AOI222xp33_ASAP7_75t_L g1428 ( 
.A1(n_1239),
.A2(n_423),
.B1(n_426),
.B2(n_429),
.C1(n_432),
.C2(n_261),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1197),
.A2(n_1154),
.B(n_1141),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1302),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1310),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1274),
.B(n_1072),
.Y(n_1432)
);

OR2x6_ASAP7_75t_L g1433 ( 
.A(n_1232),
.B(n_978),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1332),
.A2(n_1046),
.B1(n_1125),
.B2(n_987),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1260),
.A2(n_1052),
.B(n_1086),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1268),
.B(n_1040),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1251),
.B(n_1039),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_SL g1438 ( 
.A1(n_1199),
.A2(n_1125),
.B1(n_1103),
.B2(n_1046),
.Y(n_1438)
);

AO21x2_ASAP7_75t_L g1439 ( 
.A1(n_1222),
.A2(n_1079),
.B(n_1075),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1299),
.A2(n_1099),
.B(n_1086),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1314),
.Y(n_1441)
);

INVx5_ASAP7_75t_L g1442 ( 
.A(n_1197),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1197),
.Y(n_1443)
);

AO21x2_ASAP7_75t_L g1444 ( 
.A1(n_1233),
.A2(n_1096),
.B(n_1085),
.Y(n_1444)
);

AO21x2_ASAP7_75t_L g1445 ( 
.A1(n_1248),
.A2(n_1096),
.B(n_1085),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1333),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1215),
.A2(n_1281),
.B(n_1253),
.C(n_1210),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_SL g1448 ( 
.A(n_1199),
.B(n_1057),
.Y(n_1448)
);

OA21x2_ASAP7_75t_L g1449 ( 
.A1(n_1257),
.A2(n_1113),
.B(n_1112),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1279),
.Y(n_1450)
);

OAI21xp33_ASAP7_75t_SL g1451 ( 
.A1(n_1334),
.A2(n_1029),
.B(n_978),
.Y(n_1451)
);

OA21x2_ASAP7_75t_L g1452 ( 
.A1(n_1279),
.A2(n_1113),
.B(n_1112),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1245),
.Y(n_1453)
);

BUFx12f_ASAP7_75t_L g1454 ( 
.A(n_1267),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1204),
.A2(n_1188),
.B(n_1211),
.Y(n_1455)
);

BUFx4f_ASAP7_75t_SL g1456 ( 
.A(n_1173),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1184),
.A2(n_1114),
.B(n_1099),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1223),
.B(n_1020),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1226),
.A2(n_1154),
.B1(n_1141),
.B2(n_1028),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1211),
.A2(n_1114),
.B(n_1144),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_1306),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1284),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1212),
.A2(n_1158),
.B(n_1144),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1213),
.A2(n_1158),
.B(n_1044),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1285),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1268),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1249),
.Y(n_1467)
);

NAND2x1p5_ASAP7_75t_L g1468 ( 
.A(n_1224),
.B(n_1044),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1170),
.A2(n_1144),
.B(n_543),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1306),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1170),
.A2(n_1144),
.B(n_541),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1227),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1284),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1265),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1251),
.Y(n_1475)
);

BUFx12f_ASAP7_75t_L g1476 ( 
.A(n_1288),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1294),
.A2(n_1144),
.B(n_426),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1294),
.A2(n_1300),
.B(n_1297),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1297),
.A2(n_429),
.B(n_423),
.Y(n_1479)
);

OA21x2_ASAP7_75t_L g1480 ( 
.A1(n_1300),
.A2(n_1034),
.B(n_1144),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1304),
.A2(n_1144),
.B(n_1044),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_SL g1482 ( 
.A(n_1265),
.B(n_1067),
.Y(n_1482)
);

A2O1A1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1176),
.A2(n_1238),
.B(n_1326),
.C(n_1179),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1201),
.B(n_1036),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1292),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1292),
.B(n_1020),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1304),
.A2(n_1044),
.B(n_1158),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1213),
.A2(n_1185),
.B(n_1044),
.Y(n_1488)
);

NOR2xp67_ASAP7_75t_L g1489 ( 
.A(n_1265),
.B(n_1040),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1231),
.A2(n_1312),
.B(n_1311),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1308),
.A2(n_1060),
.B(n_658),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1292),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1308),
.A2(n_1060),
.B(n_658),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1309),
.B(n_1027),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1176),
.A2(n_1110),
.B(n_1091),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1309),
.B(n_1040),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1290),
.A2(n_1110),
.B1(n_1069),
.B2(n_1091),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1317),
.A2(n_1060),
.B(n_707),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1268),
.B(n_1069),
.Y(n_1499)
);

AO21x2_ASAP7_75t_L g1500 ( 
.A1(n_1224),
.A2(n_1254),
.B(n_1242),
.Y(n_1500)
);

O2A1O1Ixp33_ASAP7_75t_SL g1501 ( 
.A1(n_1242),
.A2(n_1060),
.B(n_421),
.C(n_1070),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1317),
.A2(n_1060),
.B(n_707),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1323),
.A2(n_1060),
.B(n_733),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1323),
.A2(n_1060),
.B(n_733),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1254),
.A2(n_1110),
.B1(n_1091),
.B2(n_1070),
.Y(n_1505)
);

OR2x6_ASAP7_75t_L g1506 ( 
.A(n_1277),
.B(n_1027),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1327),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1309),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1315),
.B(n_1070),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1327),
.A2(n_733),
.B(n_1091),
.Y(n_1510)
);

AO21x1_ASAP7_75t_L g1511 ( 
.A1(n_1301),
.A2(n_1110),
.B(n_421),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1315),
.B(n_1067),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1235),
.Y(n_1513)
);

AO31x2_ASAP7_75t_L g1514 ( 
.A1(n_1316),
.A2(n_12),
.A3(n_14),
.B(n_15),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1315),
.A2(n_421),
.B1(n_1103),
.B2(n_324),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1499),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1345),
.Y(n_1517)
);

AOI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1369),
.A2(n_1342),
.B1(n_1434),
.B2(n_1386),
.C(n_1395),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1428),
.A2(n_1305),
.B1(n_324),
.B2(n_430),
.Y(n_1519)
);

NOR2x1_ASAP7_75t_SL g1520 ( 
.A(n_1370),
.B(n_1301),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1499),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1499),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1393),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1366),
.Y(n_1524)
);

CKINVDCx20_ASAP7_75t_R g1525 ( 
.A(n_1360),
.Y(n_1525)
);

CKINVDCx11_ASAP7_75t_R g1526 ( 
.A(n_1358),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1456),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1426),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1355),
.Y(n_1529)
);

AOI21xp33_ASAP7_75t_L g1530 ( 
.A1(n_1422),
.A2(n_1291),
.B(n_1283),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1392),
.Y(n_1531)
);

A2O1A1Ixp33_ASAP7_75t_L g1532 ( 
.A1(n_1451),
.A2(n_1238),
.B(n_1275),
.C(n_1259),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1499),
.Y(n_1533)
);

INVx4_ASAP7_75t_L g1534 ( 
.A(n_1366),
.Y(n_1534)
);

AO31x2_ASAP7_75t_L g1535 ( 
.A1(n_1483),
.A2(n_1273),
.A3(n_1247),
.B(n_1220),
.Y(n_1535)
);

AOI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1476),
.A2(n_1321),
.B1(n_1077),
.B2(n_1042),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1467),
.A2(n_1319),
.B1(n_1321),
.B2(n_1296),
.Y(n_1537)
);

OR2x6_ASAP7_75t_L g1538 ( 
.A(n_1367),
.B(n_1296),
.Y(n_1538)
);

NAND2xp33_ASAP7_75t_R g1539 ( 
.A(n_1475),
.B(n_1287),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1393),
.Y(n_1540)
);

NAND4xp25_ASAP7_75t_L g1541 ( 
.A(n_1428),
.B(n_1321),
.C(n_1272),
.D(n_324),
.Y(n_1541)
);

AO21x2_ASAP7_75t_L g1542 ( 
.A1(n_1447),
.A2(n_1282),
.B(n_1278),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1402),
.A2(n_1221),
.B(n_1319),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1438),
.A2(n_324),
.B1(n_378),
.B2(n_377),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1405),
.B(n_1296),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1355),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1413),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_SL g1548 ( 
.A1(n_1438),
.A2(n_393),
.B1(n_392),
.B2(n_391),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1461),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1405),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1368),
.B(n_1276),
.Y(n_1551)
);

OAI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1515),
.A2(n_424),
.B1(n_353),
.B2(n_356),
.C(n_358),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1426),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1345),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1467),
.A2(n_350),
.B1(n_360),
.B2(n_364),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1476),
.A2(n_1077),
.B1(n_370),
.B2(n_389),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1454),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_1436),
.Y(n_1558)
);

NAND2xp33_ASAP7_75t_R g1559 ( 
.A(n_1475),
.B(n_1287),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1409),
.A2(n_369),
.B1(n_375),
.B2(n_434),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1337),
.A2(n_1378),
.B1(n_1349),
.B2(n_1341),
.Y(n_1561)
);

BUFx4f_ASAP7_75t_L g1562 ( 
.A(n_1366),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1416),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1387),
.A2(n_1206),
.B1(n_1313),
.B2(n_1262),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1381),
.B(n_1276),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1381),
.B(n_1276),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1337),
.A2(n_376),
.B1(n_381),
.B2(n_386),
.Y(n_1567)
);

NAND3x1_ASAP7_75t_L g1568 ( 
.A(n_1484),
.B(n_15),
.C(n_16),
.Y(n_1568)
);

BUFx12f_ASAP7_75t_L g1569 ( 
.A(n_1454),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1416),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1400),
.B(n_1276),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1359),
.B(n_1298),
.Y(n_1572)
);

CKINVDCx16_ASAP7_75t_R g1573 ( 
.A(n_1415),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1409),
.A2(n_397),
.B1(n_399),
.B2(n_401),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1361),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1361),
.Y(n_1576)
);

A2O1A1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1451),
.A2(n_1214),
.B(n_1209),
.C(n_1269),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1343),
.B(n_1298),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1405),
.B(n_1256),
.Y(n_1579)
);

OAI21x1_ASAP7_75t_L g1580 ( 
.A1(n_1478),
.A2(n_1255),
.B(n_1258),
.Y(n_1580)
);

OAI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1448),
.A2(n_406),
.B1(n_407),
.B2(n_412),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1384),
.B(n_1298),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1358),
.Y(n_1583)
);

AOI221x1_ASAP7_75t_L g1584 ( 
.A1(n_1338),
.A2(n_1220),
.B1(n_1271),
.B2(n_1331),
.C(n_1218),
.Y(n_1584)
);

NAND2x1p5_ASAP7_75t_L g1585 ( 
.A(n_1442),
.B(n_1287),
.Y(n_1585)
);

INVx3_ASAP7_75t_L g1586 ( 
.A(n_1436),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1431),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1343),
.B(n_1512),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1436),
.B(n_1237),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1359),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1512),
.B(n_1298),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1465),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1354),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1417),
.B(n_1241),
.Y(n_1594)
);

OAI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1478),
.A2(n_1318),
.B(n_1313),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1417),
.B(n_1241),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1367),
.A2(n_1352),
.B1(n_1490),
.B2(n_1389),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1367),
.A2(n_16),
.B1(n_17),
.B2(n_20),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_SL g1599 ( 
.A1(n_1448),
.A2(n_1303),
.B1(n_1289),
.B2(n_1220),
.Y(n_1599)
);

OR2x6_ASAP7_75t_L g1600 ( 
.A(n_1367),
.B(n_1220),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1465),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1367),
.A2(n_20),
.B1(n_25),
.B2(n_26),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1430),
.B(n_1351),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1415),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1414),
.B(n_1241),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1509),
.B(n_1241),
.Y(n_1606)
);

CKINVDCx6p67_ASAP7_75t_R g1607 ( 
.A(n_1458),
.Y(n_1607)
);

CKINVDCx20_ASAP7_75t_R g1608 ( 
.A(n_1437),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1424),
.B(n_566),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1444),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1352),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1453),
.B(n_28),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1441),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_SL g1614 ( 
.A1(n_1459),
.A2(n_215),
.B(n_208),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1354),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1458),
.Y(n_1616)
);

NAND2xp33_ASAP7_75t_R g1617 ( 
.A(n_1480),
.B(n_108),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1446),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1445),
.A2(n_566),
.B(n_200),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1444),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1362),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1446),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1356),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1490),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_1624)
);

NAND2x1p5_ASAP7_75t_L g1625 ( 
.A(n_1442),
.B(n_566),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1436),
.B(n_199),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_SL g1627 ( 
.A1(n_1372),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1490),
.A2(n_1389),
.B1(n_1433),
.B2(n_1453),
.Y(n_1628)
);

A2O1A1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1385),
.A2(n_39),
.B(n_43),
.C(n_44),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1356),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1357),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1370),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_SL g1633 ( 
.A1(n_1482),
.A2(n_43),
.B1(n_44),
.B2(n_48),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1509),
.B(n_48),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1474),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1362),
.B(n_198),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1410),
.A2(n_1379),
.B1(n_1492),
.B2(n_1508),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1470),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1357),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1492),
.B(n_50),
.Y(n_1640)
);

OAI22xp33_ASAP7_75t_SL g1641 ( 
.A1(n_1482),
.A2(n_50),
.B1(n_53),
.B2(n_55),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1364),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1508),
.A2(n_566),
.B1(n_56),
.B2(n_57),
.Y(n_1643)
);

NAND2xp33_ASAP7_75t_L g1644 ( 
.A(n_1370),
.B(n_53),
.Y(n_1644)
);

OAI222xp33_ASAP7_75t_L g1645 ( 
.A1(n_1433),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.C1(n_61),
.C2(n_65),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1513),
.B(n_59),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1486),
.A2(n_1494),
.B1(n_1506),
.B2(n_1485),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_SL g1648 ( 
.A1(n_1370),
.A2(n_118),
.B(n_196),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1364),
.Y(n_1649)
);

INVx4_ASAP7_75t_L g1650 ( 
.A(n_1370),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1432),
.Y(n_1651)
);

O2A1O1Ixp33_ASAP7_75t_SL g1652 ( 
.A1(n_1463),
.A2(n_65),
.B(n_67),
.C(n_68),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1470),
.Y(n_1653)
);

BUFx10_ASAP7_75t_L g1654 ( 
.A(n_1336),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1397),
.B(n_1348),
.Y(n_1655)
);

CKINVDCx6p67_ASAP7_75t_R g1656 ( 
.A(n_1506),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_L g1657 ( 
.A1(n_1420),
.A2(n_120),
.B(n_194),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1513),
.B(n_68),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1336),
.Y(n_1659)
);

CKINVDCx16_ASAP7_75t_R g1660 ( 
.A(n_1397),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1344),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1506),
.A2(n_566),
.B1(n_75),
.B2(n_76),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1496),
.B(n_70),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1403),
.B(n_75),
.Y(n_1664)
);

NAND2x1_ASAP7_75t_L g1665 ( 
.A(n_1336),
.B(n_129),
.Y(n_1665)
);

OAI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1376),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.C(n_79),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1403),
.B(n_77),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1344),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1433),
.A2(n_79),
.B1(n_80),
.B2(n_83),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1348),
.B(n_142),
.Y(n_1670)
);

AOI222xp33_ASAP7_75t_L g1671 ( 
.A1(n_1376),
.A2(n_80),
.B1(n_84),
.B2(n_88),
.C1(n_90),
.C2(n_92),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1506),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_1672)
);

INVx4_ASAP7_75t_L g1673 ( 
.A(n_1383),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1350),
.Y(n_1674)
);

AOI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1472),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.C(n_110),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1348),
.B(n_99),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1348),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1445),
.A2(n_193),
.B(n_131),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1506),
.A2(n_113),
.B1(n_133),
.B2(n_146),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1466),
.B(n_152),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1466),
.B(n_156),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1432),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1336),
.Y(n_1683)
);

AOI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1466),
.A2(n_159),
.B1(n_161),
.B2(n_163),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1472),
.B(n_190),
.Y(n_1685)
);

NAND2xp33_ASAP7_75t_R g1686 ( 
.A(n_1480),
.B(n_1335),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1474),
.Y(n_1687)
);

BUFx2_ASAP7_75t_L g1688 ( 
.A(n_1373),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1373),
.B(n_165),
.Y(n_1689)
);

NAND2xp33_ASAP7_75t_R g1690 ( 
.A(n_1480),
.B(n_182),
.Y(n_1690)
);

INVx4_ASAP7_75t_L g1691 ( 
.A(n_1383),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_SL g1692 ( 
.A1(n_1445),
.A2(n_166),
.B1(n_172),
.B2(n_173),
.Y(n_1692)
);

A2O1A1Ixp33_ASAP7_75t_L g1693 ( 
.A1(n_1464),
.A2(n_178),
.B(n_1495),
.C(n_1401),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1449),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1497),
.A2(n_1433),
.B1(n_1505),
.B2(n_1468),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1373),
.B(n_1382),
.Y(n_1696)
);

OA21x2_ASAP7_75t_L g1697 ( 
.A1(n_1469),
.A2(n_1471),
.B(n_1419),
.Y(n_1697)
);

INVx1_ASAP7_75t_SL g1698 ( 
.A(n_1373),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1444),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1433),
.A2(n_1511),
.B1(n_1340),
.B2(n_1382),
.Y(n_1700)
);

INVx4_ASAP7_75t_L g1701 ( 
.A(n_1383),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1382),
.B(n_1489),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1382),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1457),
.Y(n_1704)
);

OAI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1442),
.A2(n_1391),
.B1(n_1383),
.B2(n_1401),
.Y(n_1705)
);

BUFx2_ASAP7_75t_L g1706 ( 
.A(n_1474),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1518),
.B(n_1474),
.Y(n_1707)
);

OAI22xp33_ASAP7_75t_SL g1708 ( 
.A1(n_1666),
.A2(n_1468),
.B1(n_1495),
.B2(n_1514),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1671),
.A2(n_1511),
.B1(n_1340),
.B2(n_1439),
.Y(n_1709)
);

OR2x6_ASAP7_75t_L g1710 ( 
.A(n_1538),
.B(n_1469),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1541),
.A2(n_1439),
.B1(n_1394),
.B2(n_1480),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_SL g1712 ( 
.A1(n_1644),
.A2(n_1460),
.B1(n_1439),
.B2(n_1383),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1660),
.B(n_1514),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1544),
.A2(n_1468),
.B1(n_1489),
.B2(n_1391),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1523),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1616),
.B(n_1588),
.Y(n_1716)
);

AOI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1574),
.A2(n_1544),
.B1(n_1611),
.B2(n_1567),
.C(n_1552),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1540),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1667),
.B(n_1514),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1590),
.B(n_1514),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1548),
.A2(n_1500),
.B1(n_1474),
.B2(n_1460),
.Y(n_1721)
);

INVx4_ASAP7_75t_L g1722 ( 
.A(n_1562),
.Y(n_1722)
);

OAI21x1_ASAP7_75t_L g1723 ( 
.A1(n_1580),
.A2(n_1471),
.B(n_1477),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1543),
.A2(n_1488),
.B(n_1442),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1676),
.B(n_1514),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1591),
.B(n_1500),
.Y(n_1726)
);

AOI222xp33_ASAP7_75t_L g1727 ( 
.A1(n_1574),
.A2(n_1399),
.B1(n_1406),
.B2(n_1380),
.C1(n_1462),
.C2(n_1425),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1607),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1638),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1611),
.A2(n_1394),
.B1(n_1500),
.B2(n_1460),
.Y(n_1730)
);

AOI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1705),
.A2(n_1442),
.B(n_1363),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1634),
.B(n_1455),
.Y(n_1732)
);

NAND2x1p5_ASAP7_75t_L g1733 ( 
.A(n_1562),
.B(n_1442),
.Y(n_1733)
);

BUFx4f_ASAP7_75t_SL g1734 ( 
.A(n_1549),
.Y(n_1734)
);

OAI321xp33_ASAP7_75t_L g1735 ( 
.A1(n_1669),
.A2(n_1602),
.A3(n_1598),
.B1(n_1624),
.B2(n_1672),
.C(n_1629),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1603),
.B(n_1394),
.Y(n_1736)
);

A2O1A1Ixp33_ASAP7_75t_L g1737 ( 
.A1(n_1629),
.A2(n_1429),
.B(n_1487),
.C(n_1457),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1655),
.B(n_1455),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1548),
.A2(n_1394),
.B1(n_1455),
.B2(n_1339),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1572),
.B(n_1377),
.Y(n_1740)
);

OAI22x1_ASAP7_75t_L g1741 ( 
.A1(n_1647),
.A2(n_1407),
.B1(n_1380),
.B2(n_1406),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1669),
.A2(n_1339),
.B1(n_1377),
.B2(n_1398),
.Y(n_1742)
);

BUFx6f_ASAP7_75t_L g1743 ( 
.A(n_1632),
.Y(n_1743)
);

AOI211xp5_ASAP7_75t_L g1744 ( 
.A1(n_1581),
.A2(n_1501),
.B(n_1391),
.C(n_1412),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1655),
.B(n_1391),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1598),
.A2(n_1339),
.B1(n_1377),
.B2(n_1398),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1602),
.A2(n_1398),
.B1(n_1391),
.B2(n_1423),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1610),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1547),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1603),
.B(n_1335),
.Y(n_1750)
);

BUFx2_ASAP7_75t_L g1751 ( 
.A(n_1687),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1627),
.A2(n_1633),
.B1(n_1675),
.B2(n_1567),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1563),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1651),
.B(n_1682),
.Y(n_1754)
);

OAI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1560),
.A2(n_1396),
.B1(n_1423),
.B2(n_1443),
.C(n_1404),
.Y(n_1755)
);

NAND3xp33_ASAP7_75t_L g1756 ( 
.A(n_1627),
.B(n_1479),
.C(n_1407),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1561),
.A2(n_1396),
.B1(n_1423),
.B2(n_1443),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1561),
.A2(n_1396),
.B1(n_1443),
.B2(n_1404),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1570),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1565),
.B(n_1407),
.Y(n_1760)
);

OAI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1581),
.A2(n_1390),
.B1(n_1404),
.B2(n_1399),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1566),
.B(n_1479),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1587),
.Y(n_1763)
);

BUFx2_ASAP7_75t_L g1764 ( 
.A(n_1524),
.Y(n_1764)
);

OAI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1519),
.A2(n_1390),
.B1(n_1507),
.B2(n_1425),
.C(n_1421),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1677),
.B(n_1479),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1688),
.B(n_1479),
.Y(n_1767)
);

AOI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1608),
.A2(n_1371),
.B1(n_1507),
.B2(n_1427),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1573),
.A2(n_1371),
.B1(n_1421),
.B2(n_1462),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1663),
.B(n_1412),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1624),
.A2(n_1371),
.B1(n_1407),
.B2(n_1449),
.Y(n_1771)
);

A2O1A1Ixp33_ASAP7_75t_L g1772 ( 
.A1(n_1693),
.A2(n_1487),
.B(n_1419),
.C(n_1418),
.Y(n_1772)
);

INVx2_ASAP7_75t_SL g1773 ( 
.A(n_1527),
.Y(n_1773)
);

CKINVDCx11_ASAP7_75t_R g1774 ( 
.A(n_1525),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1528),
.B(n_1553),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1633),
.A2(n_1449),
.B1(n_1452),
.B2(n_1427),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1613),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1531),
.B(n_1374),
.Y(n_1778)
);

OAI211xp5_ASAP7_75t_L g1779 ( 
.A1(n_1519),
.A2(n_1450),
.B(n_1473),
.C(n_1420),
.Y(n_1779)
);

OAI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1555),
.A2(n_1450),
.B1(n_1473),
.B2(n_1449),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_SL g1781 ( 
.A1(n_1641),
.A2(n_1481),
.B1(n_1452),
.B2(n_1374),
.Y(n_1781)
);

OAI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1555),
.A2(n_1452),
.B1(n_1418),
.B2(n_1346),
.C(n_1347),
.Y(n_1782)
);

OAI21x1_ASAP7_75t_L g1783 ( 
.A1(n_1657),
.A2(n_1595),
.B(n_1435),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1640),
.A2(n_1452),
.B1(n_1346),
.B2(n_1353),
.Y(n_1784)
);

OAI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1536),
.A2(n_1411),
.B1(n_1388),
.B2(n_1408),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1592),
.Y(n_1786)
);

CKINVDCx11_ASAP7_75t_R g1787 ( 
.A(n_1526),
.Y(n_1787)
);

AOI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1692),
.A2(n_1347),
.B1(n_1510),
.B2(n_1353),
.Y(n_1788)
);

OAI21xp5_ASAP7_75t_SL g1789 ( 
.A1(n_1645),
.A2(n_1411),
.B(n_1510),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1618),
.Y(n_1790)
);

A2O1A1Ixp33_ASAP7_75t_L g1791 ( 
.A1(n_1693),
.A2(n_1408),
.B(n_1388),
.C(n_1504),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1637),
.A2(n_1440),
.B1(n_1375),
.B2(n_1435),
.Y(n_1792)
);

AOI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1652),
.A2(n_1365),
.B1(n_1440),
.B2(n_1375),
.C(n_1504),
.Y(n_1793)
);

AOI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1604),
.A2(n_1365),
.B1(n_1491),
.B2(n_1493),
.Y(n_1794)
);

AOI222xp33_ASAP7_75t_L g1795 ( 
.A1(n_1643),
.A2(n_1491),
.B1(n_1493),
.B2(n_1498),
.C1(n_1502),
.C2(n_1503),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1593),
.Y(n_1796)
);

OAI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1539),
.A2(n_1498),
.B1(n_1502),
.B2(n_1503),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_SL g1798 ( 
.A1(n_1640),
.A2(n_1662),
.B1(n_1695),
.B2(n_1679),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1692),
.A2(n_1586),
.B1(n_1558),
.B2(n_1516),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1696),
.B(n_1517),
.Y(n_1800)
);

NAND3xp33_ASAP7_75t_SL g1801 ( 
.A(n_1684),
.B(n_1678),
.C(n_1646),
.Y(n_1801)
);

BUFx6f_ASAP7_75t_L g1802 ( 
.A(n_1632),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1653),
.A2(n_1601),
.B1(n_1531),
.B2(n_1524),
.Y(n_1803)
);

OAI21x1_ASAP7_75t_L g1804 ( 
.A1(n_1619),
.A2(n_1585),
.B(n_1704),
.Y(n_1804)
);

AOI221xp5_ASAP7_75t_L g1805 ( 
.A1(n_1652),
.A2(n_1530),
.B1(n_1658),
.B2(n_1612),
.C(n_1664),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1698),
.B(n_1703),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1578),
.B(n_1516),
.Y(n_1807)
);

A2O1A1Ixp33_ASAP7_75t_L g1808 ( 
.A1(n_1532),
.A2(n_1577),
.B(n_1599),
.C(n_1653),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1528),
.A2(n_1553),
.B1(n_1626),
.B2(n_1551),
.Y(n_1809)
);

OAI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1556),
.A2(n_1532),
.B1(n_1577),
.B2(n_1617),
.C(n_1690),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1626),
.A2(n_1571),
.B1(n_1526),
.B2(n_1582),
.Y(n_1811)
);

NAND3xp33_ASAP7_75t_L g1812 ( 
.A(n_1617),
.B(n_1690),
.C(n_1685),
.Y(n_1812)
);

OAI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1700),
.A2(n_1599),
.B1(n_1597),
.B2(n_1628),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1631),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1568),
.A2(n_1670),
.B1(n_1583),
.B2(n_1554),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1594),
.B(n_1596),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1700),
.A2(n_1597),
.B1(n_1628),
.B2(n_1534),
.Y(n_1817)
);

OA21x2_ASAP7_75t_L g1818 ( 
.A1(n_1584),
.A2(n_1699),
.B(n_1694),
.Y(n_1818)
);

NAND3xp33_ASAP7_75t_L g1819 ( 
.A(n_1539),
.B(n_1559),
.C(n_1537),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1557),
.A2(n_1569),
.B1(n_1586),
.B2(n_1558),
.Y(n_1820)
);

AOI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1670),
.A2(n_1689),
.B1(n_1521),
.B2(n_1522),
.Y(n_1821)
);

OAI211xp5_ASAP7_75t_L g1822 ( 
.A1(n_1614),
.A2(n_1648),
.B(n_1605),
.C(n_1622),
.Y(n_1822)
);

BUFx6f_ASAP7_75t_L g1823 ( 
.A(n_1632),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1534),
.A2(n_1656),
.B1(n_1621),
.B2(n_1702),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1521),
.A2(n_1522),
.B1(n_1533),
.B2(n_1689),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1533),
.A2(n_1636),
.B1(n_1538),
.B2(n_1606),
.Y(n_1826)
);

HB1xp67_ASAP7_75t_L g1827 ( 
.A(n_1610),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_SL g1828 ( 
.A1(n_1564),
.A2(n_1600),
.B1(n_1520),
.B2(n_1636),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1538),
.A2(n_1550),
.B1(n_1589),
.B2(n_1579),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1576),
.B(n_1642),
.Y(n_1830)
);

INVxp67_ASAP7_75t_L g1831 ( 
.A(n_1623),
.Y(n_1831)
);

AND2x6_ASAP7_75t_L g1832 ( 
.A(n_1681),
.B(n_1589),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1661),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1615),
.B(n_1630),
.Y(n_1834)
);

AOI21xp33_ASAP7_75t_L g1835 ( 
.A1(n_1559),
.A2(n_1609),
.B(n_1542),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1579),
.A2(n_1683),
.B1(n_1659),
.B2(n_1680),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1681),
.A2(n_1609),
.B1(n_1639),
.B2(n_1649),
.Y(n_1837)
);

AO31x2_ASAP7_75t_L g1838 ( 
.A1(n_1694),
.A2(n_1668),
.A3(n_1674),
.B(n_1630),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1615),
.Y(n_1839)
);

CKINVDCx20_ASAP7_75t_R g1840 ( 
.A(n_1706),
.Y(n_1840)
);

AOI222xp33_ASAP7_75t_L g1841 ( 
.A1(n_1705),
.A2(n_1620),
.B1(n_1529),
.B2(n_1546),
.C1(n_1575),
.C2(n_1545),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1545),
.B(n_1635),
.Y(n_1842)
);

AOI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1665),
.A2(n_1635),
.B1(n_1691),
.B2(n_1673),
.Y(n_1843)
);

AOI32xp33_ASAP7_75t_L g1844 ( 
.A1(n_1650),
.A2(n_1701),
.A3(n_1691),
.B1(n_1673),
.B2(n_1620),
.Y(n_1844)
);

OAI21x1_ASAP7_75t_L g1845 ( 
.A1(n_1585),
.A2(n_1697),
.B(n_1529),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1654),
.B(n_1632),
.Y(n_1846)
);

OAI211xp5_ASAP7_75t_L g1847 ( 
.A1(n_1546),
.A2(n_1575),
.B(n_1701),
.C(n_1650),
.Y(n_1847)
);

OAI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1600),
.A2(n_1686),
.B1(n_1625),
.B2(n_1697),
.Y(n_1848)
);

OAI21xp33_ASAP7_75t_L g1849 ( 
.A1(n_1600),
.A2(n_1625),
.B(n_1686),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1697),
.A2(n_1654),
.B1(n_1542),
.B2(n_1535),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1535),
.Y(n_1851)
);

BUFx4f_ASAP7_75t_SL g1852 ( 
.A(n_1535),
.Y(n_1852)
);

INVx4_ASAP7_75t_L g1853 ( 
.A(n_1562),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1544),
.A2(n_1116),
.B1(n_1386),
.B2(n_819),
.Y(n_1854)
);

OA21x2_ASAP7_75t_L g1855 ( 
.A1(n_1584),
.A2(n_1471),
.B(n_1469),
.Y(n_1855)
);

AOI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1518),
.A2(n_819),
.B1(n_1116),
.B2(n_1386),
.Y(n_1856)
);

AOI221xp5_ASAP7_75t_L g1857 ( 
.A1(n_1574),
.A2(n_819),
.B1(n_1172),
.B2(n_446),
.C(n_1666),
.Y(n_1857)
);

BUFx3_ASAP7_75t_L g1858 ( 
.A(n_1638),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1518),
.A2(n_1172),
.B1(n_1026),
.B2(n_819),
.Y(n_1859)
);

A2O1A1Ixp33_ASAP7_75t_L g1860 ( 
.A1(n_1518),
.A2(n_1172),
.B(n_1116),
.C(n_819),
.Y(n_1860)
);

NAND3xp33_ASAP7_75t_L g1861 ( 
.A(n_1518),
.B(n_1172),
.C(n_819),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_SL g1862 ( 
.A1(n_1629),
.A2(n_1177),
.B(n_1116),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1523),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1588),
.B(n_1660),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_SL g1865 ( 
.A1(n_1666),
.A2(n_819),
.B1(n_1116),
.B2(n_1644),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1518),
.B(n_1369),
.Y(n_1866)
);

OR2x6_ASAP7_75t_L g1867 ( 
.A(n_1538),
.B(n_1614),
.Y(n_1867)
);

AOI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1518),
.A2(n_1172),
.B1(n_1026),
.B2(n_819),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1593),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1660),
.B(n_1572),
.Y(n_1870)
);

BUFx3_ASAP7_75t_L g1871 ( 
.A(n_1638),
.Y(n_1871)
);

OAI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1541),
.A2(n_1666),
.B1(n_1180),
.B2(n_1172),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1544),
.A2(n_1116),
.B1(n_1386),
.B2(n_819),
.Y(n_1873)
);

BUFx6f_ASAP7_75t_L g1874 ( 
.A(n_1562),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1523),
.Y(n_1875)
);

OAI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1544),
.A2(n_1116),
.B1(n_1386),
.B2(n_819),
.Y(n_1876)
);

OAI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1541),
.A2(n_1666),
.B1(n_1180),
.B2(n_1172),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1660),
.B(n_1572),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1588),
.B(n_1660),
.Y(n_1879)
);

AOI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1574),
.A2(n_819),
.B1(n_1172),
.B2(n_446),
.C(n_1666),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1518),
.A2(n_1172),
.B1(n_1026),
.B2(n_819),
.Y(n_1881)
);

AOI221xp5_ASAP7_75t_L g1882 ( 
.A1(n_1574),
.A2(n_819),
.B1(n_1172),
.B2(n_446),
.C(n_1666),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1518),
.A2(n_1172),
.B1(n_1026),
.B2(n_819),
.Y(n_1883)
);

AOI221xp5_ASAP7_75t_L g1884 ( 
.A1(n_1574),
.A2(n_819),
.B1(n_1172),
.B2(n_446),
.C(n_1666),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1838),
.Y(n_1885)
);

AOI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1862),
.A2(n_1860),
.B(n_1810),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1710),
.B(n_1738),
.Y(n_1887)
);

OR2x6_ASAP7_75t_L g1888 ( 
.A(n_1710),
.B(n_1867),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1833),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1856),
.B(n_1854),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1748),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1726),
.B(n_1732),
.Y(n_1892)
);

INVxp67_ASAP7_75t_L g1893 ( 
.A(n_1716),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1710),
.B(n_1845),
.Y(n_1894)
);

INVx2_ASAP7_75t_SL g1895 ( 
.A(n_1775),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1725),
.B(n_1807),
.Y(n_1896)
);

INVx2_ASAP7_75t_SL g1897 ( 
.A(n_1764),
.Y(n_1897)
);

AOI222xp33_ASAP7_75t_L g1898 ( 
.A1(n_1717),
.A2(n_1884),
.B1(n_1857),
.B2(n_1882),
.C1(n_1880),
.C2(n_1861),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1839),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1734),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1715),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1718),
.Y(n_1902)
);

BUFx2_ASAP7_75t_L g1903 ( 
.A(n_1748),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1719),
.B(n_1762),
.Y(n_1904)
);

INVxp67_ASAP7_75t_L g1905 ( 
.A(n_1786),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1866),
.B(n_1750),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1749),
.Y(n_1907)
);

INVx5_ASAP7_75t_SL g1908 ( 
.A(n_1867),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1736),
.B(n_1816),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1740),
.B(n_1760),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1870),
.B(n_1878),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1753),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1770),
.B(n_1759),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1827),
.B(n_1720),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1864),
.B(n_1879),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1827),
.B(n_1713),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1763),
.Y(n_1917)
);

BUFx3_ASAP7_75t_L g1918 ( 
.A(n_1840),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1769),
.B(n_1768),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1777),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1790),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1863),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1806),
.B(n_1805),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1875),
.B(n_1767),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1818),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1796),
.B(n_1814),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1873),
.B(n_1876),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1869),
.B(n_1754),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1811),
.B(n_1831),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1766),
.B(n_1813),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1811),
.B(n_1809),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1778),
.B(n_1818),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1834),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1851),
.Y(n_1934)
);

AOI21x1_ASAP7_75t_L g1935 ( 
.A1(n_1731),
.A2(n_1724),
.B(n_1785),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1809),
.B(n_1830),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1741),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1849),
.B(n_1730),
.Y(n_1938)
);

OR2x2_ASAP7_75t_L g1939 ( 
.A(n_1848),
.B(n_1817),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1852),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1730),
.B(n_1739),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1852),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1808),
.B(n_1712),
.Y(n_1943)
);

HB1xp67_ASAP7_75t_L g1944 ( 
.A(n_1803),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1842),
.B(n_1859),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1855),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1783),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1712),
.B(n_1784),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1784),
.B(n_1776),
.Y(n_1949)
);

AOI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1868),
.A2(n_1883),
.B1(n_1881),
.B2(n_1865),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1855),
.Y(n_1951)
);

AND2x4_ASAP7_75t_SL g1952 ( 
.A(n_1867),
.B(n_1874),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1800),
.B(n_1837),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1776),
.B(n_1835),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1723),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1850),
.Y(n_1956)
);

NOR2x1_ASAP7_75t_SL g1957 ( 
.A(n_1819),
.B(n_1822),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1828),
.B(n_1742),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1780),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1828),
.B(n_1746),
.Y(n_1960)
);

INVx2_ASAP7_75t_SL g1961 ( 
.A(n_1743),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1837),
.B(n_1872),
.Y(n_1962)
);

BUFx2_ASAP7_75t_L g1963 ( 
.A(n_1804),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1721),
.B(n_1841),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1782),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1848),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1826),
.B(n_1781),
.Y(n_1967)
);

INVx5_ASAP7_75t_SL g1968 ( 
.A(n_1874),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1792),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1781),
.B(n_1771),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1794),
.Y(n_1971)
);

BUFx2_ASAP7_75t_L g1972 ( 
.A(n_1829),
.Y(n_1972)
);

AO21x2_ASAP7_75t_L g1973 ( 
.A1(n_1791),
.A2(n_1737),
.B(n_1772),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1708),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1711),
.B(n_1771),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1711),
.B(n_1745),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1743),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1727),
.B(n_1709),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1709),
.B(n_1747),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1756),
.Y(n_1980)
);

HB1xp67_ASAP7_75t_L g1981 ( 
.A(n_1824),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1799),
.B(n_1798),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1789),
.B(n_1812),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1798),
.B(n_1788),
.Y(n_1984)
);

INVxp67_ASAP7_75t_SL g1985 ( 
.A(n_1761),
.Y(n_1985)
);

BUFx3_ASAP7_75t_L g1986 ( 
.A(n_1728),
.Y(n_1986)
);

NOR2x1_ASAP7_75t_L g1987 ( 
.A(n_1847),
.B(n_1801),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1779),
.B(n_1836),
.Y(n_1988)
);

OAI332xp33_ASAP7_75t_SL g1989 ( 
.A1(n_1872),
.A2(n_1877),
.A3(n_1714),
.B1(n_1761),
.B2(n_1758),
.B3(n_1757),
.C1(n_1797),
.C2(n_1787),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1797),
.Y(n_1990)
);

INVx1_ASAP7_75t_SL g1991 ( 
.A(n_1900),
.Y(n_1991)
);

AO21x2_ASAP7_75t_L g1992 ( 
.A1(n_1927),
.A2(n_1925),
.B(n_1946),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1907),
.Y(n_1993)
);

INVxp67_ASAP7_75t_SL g1994 ( 
.A(n_1914),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1907),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1917),
.Y(n_1996)
);

BUFx2_ASAP7_75t_L g1997 ( 
.A(n_1986),
.Y(n_1997)
);

AOI211xp5_ASAP7_75t_L g1998 ( 
.A1(n_1890),
.A2(n_1877),
.B(n_1735),
.C(n_1801),
.Y(n_1998)
);

OAI21xp33_ASAP7_75t_SL g1999 ( 
.A1(n_1943),
.A2(n_1815),
.B(n_1752),
.Y(n_1999)
);

AOI22xp33_ASAP7_75t_L g2000 ( 
.A1(n_1898),
.A2(n_1865),
.B1(n_1707),
.B2(n_1765),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1917),
.Y(n_2001)
);

OAI321xp33_ASAP7_75t_L g2002 ( 
.A1(n_1886),
.A2(n_1755),
.A3(n_1844),
.B1(n_1744),
.B2(n_1843),
.C(n_1820),
.Y(n_2002)
);

NAND3xp33_ASAP7_75t_L g2003 ( 
.A(n_1950),
.B(n_1820),
.C(n_1825),
.Y(n_2003)
);

NAND2xp33_ASAP7_75t_R g2004 ( 
.A(n_1943),
.B(n_1751),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1921),
.Y(n_2005)
);

AO21x2_ASAP7_75t_L g2006 ( 
.A1(n_1925),
.A2(n_1846),
.B(n_1821),
.Y(n_2006)
);

AOI221xp5_ASAP7_75t_L g2007 ( 
.A1(n_1974),
.A2(n_1773),
.B1(n_1729),
.B2(n_1871),
.C(n_1858),
.Y(n_2007)
);

BUFx3_ASAP7_75t_L g2008 ( 
.A(n_1986),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1921),
.Y(n_2009)
);

OAI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1982),
.A2(n_1722),
.B1(n_1853),
.B2(n_1874),
.Y(n_2010)
);

A2O1A1Ixp33_ASAP7_75t_L g2011 ( 
.A1(n_1987),
.A2(n_1874),
.B(n_1793),
.C(n_1832),
.Y(n_2011)
);

OA21x2_ASAP7_75t_L g2012 ( 
.A1(n_1946),
.A2(n_1795),
.B(n_1823),
.Y(n_2012)
);

AND2x4_ASAP7_75t_L g2013 ( 
.A(n_1894),
.B(n_1802),
.Y(n_2013)
);

AOI22xp33_ASAP7_75t_L g2014 ( 
.A1(n_1982),
.A2(n_1734),
.B1(n_1832),
.B2(n_1853),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1922),
.Y(n_2015)
);

BUFx3_ASAP7_75t_L g2016 ( 
.A(n_1986),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1922),
.Y(n_2017)
);

OAI22xp33_ASAP7_75t_L g2018 ( 
.A1(n_1962),
.A2(n_1722),
.B1(n_1733),
.B2(n_1802),
.Y(n_2018)
);

OAI22xp5_ASAP7_75t_L g2019 ( 
.A1(n_1984),
.A2(n_1733),
.B1(n_1823),
.B2(n_1832),
.Y(n_2019)
);

AOI221xp5_ASAP7_75t_L g2020 ( 
.A1(n_1974),
.A2(n_1774),
.B1(n_1823),
.B2(n_1832),
.C(n_1984),
.Y(n_2020)
);

OAI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1987),
.A2(n_1823),
.B(n_1983),
.Y(n_2021)
);

HB1xp67_ASAP7_75t_L g2022 ( 
.A(n_1891),
.Y(n_2022)
);

OR2x2_ASAP7_75t_L g2023 ( 
.A(n_1910),
.B(n_1909),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1902),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_1910),
.B(n_1909),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1902),
.Y(n_2026)
);

NOR4xp25_ASAP7_75t_SL g2027 ( 
.A(n_1963),
.B(n_1972),
.C(n_1980),
.D(n_1966),
.Y(n_2027)
);

OAI22xp33_ASAP7_75t_L g2028 ( 
.A1(n_1931),
.A2(n_1939),
.B1(n_1983),
.B2(n_1919),
.Y(n_2028)
);

AND2x6_ASAP7_75t_L g2029 ( 
.A(n_1908),
.B(n_1968),
.Y(n_2029)
);

OAI211xp5_ASAP7_75t_L g2030 ( 
.A1(n_1980),
.A2(n_1970),
.B(n_1948),
.C(n_1964),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1912),
.Y(n_2031)
);

BUFx2_ASAP7_75t_L g2032 ( 
.A(n_1897),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1896),
.B(n_1892),
.Y(n_2033)
);

AOI22xp33_ASAP7_75t_L g2034 ( 
.A1(n_1979),
.A2(n_1978),
.B1(n_1964),
.B2(n_1958),
.Y(n_2034)
);

NOR2x1p5_ASAP7_75t_L g2035 ( 
.A(n_1953),
.B(n_1929),
.Y(n_2035)
);

BUFx2_ASAP7_75t_L g2036 ( 
.A(n_1897),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1894),
.B(n_1887),
.Y(n_2037)
);

AOI22xp33_ASAP7_75t_SL g2038 ( 
.A1(n_1957),
.A2(n_1979),
.B1(n_1958),
.B2(n_1960),
.Y(n_2038)
);

AND2x4_ASAP7_75t_L g2039 ( 
.A(n_1894),
.B(n_1887),
.Y(n_2039)
);

HB1xp67_ASAP7_75t_L g2040 ( 
.A(n_1891),
.Y(n_2040)
);

OR2x2_ASAP7_75t_L g2041 ( 
.A(n_1892),
.B(n_1916),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1912),
.Y(n_2042)
);

AOI221x1_ASAP7_75t_SL g2043 ( 
.A1(n_1906),
.A2(n_1923),
.B1(n_1971),
.B2(n_1990),
.C(n_1937),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1904),
.B(n_1911),
.Y(n_2044)
);

NAND4xp25_ASAP7_75t_L g2045 ( 
.A(n_1945),
.B(n_1971),
.C(n_1937),
.D(n_1936),
.Y(n_2045)
);

INVxp67_ASAP7_75t_L g2046 ( 
.A(n_1895),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1912),
.Y(n_2047)
);

OR2x2_ASAP7_75t_L g2048 ( 
.A(n_1916),
.B(n_1914),
.Y(n_2048)
);

OAI22xp33_ASAP7_75t_L g2049 ( 
.A1(n_1939),
.A2(n_1919),
.B1(n_1975),
.B2(n_1978),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1920),
.Y(n_2050)
);

NOR2x1_ASAP7_75t_L g2051 ( 
.A(n_1918),
.B(n_1988),
.Y(n_2051)
);

AOI221xp5_ASAP7_75t_L g2052 ( 
.A1(n_1970),
.A2(n_1948),
.B1(n_1954),
.B2(n_1949),
.C(n_1965),
.Y(n_2052)
);

BUFx2_ASAP7_75t_L g2053 ( 
.A(n_1977),
.Y(n_2053)
);

NOR2xp33_ASAP7_75t_L g2054 ( 
.A(n_1981),
.B(n_1957),
.Y(n_2054)
);

NOR2x1_ASAP7_75t_L g2055 ( 
.A(n_1918),
.B(n_1988),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_1895),
.B(n_1903),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1920),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1889),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_SL g2059 ( 
.A1(n_1960),
.A2(n_1967),
.B1(n_1941),
.B2(n_1938),
.Y(n_2059)
);

BUFx2_ASAP7_75t_L g2060 ( 
.A(n_1977),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_R g2061 ( 
.A(n_1918),
.B(n_1977),
.Y(n_2061)
);

OAI33xp33_ASAP7_75t_L g2062 ( 
.A1(n_1932),
.A2(n_1893),
.A3(n_1934),
.B1(n_1933),
.B2(n_1990),
.B3(n_1928),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1924),
.B(n_1976),
.Y(n_2063)
);

OAI22xp33_ASAP7_75t_L g2064 ( 
.A1(n_1975),
.A2(n_1985),
.B1(n_1944),
.B2(n_1972),
.Y(n_2064)
);

OAI211xp5_ASAP7_75t_L g2065 ( 
.A1(n_1954),
.A2(n_1949),
.B(n_1941),
.C(n_1966),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1901),
.Y(n_2066)
);

OAI21x1_ASAP7_75t_L g2067 ( 
.A1(n_1935),
.A2(n_1947),
.B(n_1955),
.Y(n_2067)
);

OR2x2_ASAP7_75t_SL g2068 ( 
.A(n_1915),
.B(n_1965),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1899),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_2063),
.B(n_1925),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1994),
.B(n_1932),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_1992),
.B(n_1956),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2063),
.B(n_1956),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2033),
.B(n_1938),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_2037),
.B(n_1894),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2069),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2024),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2037),
.B(n_1973),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_2037),
.B(n_1973),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2026),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2048),
.B(n_1913),
.Y(n_2081)
);

INVx2_ASAP7_75t_SL g2082 ( 
.A(n_2039),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2039),
.B(n_1973),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2031),
.Y(n_2084)
);

BUFx2_ASAP7_75t_L g2085 ( 
.A(n_2061),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2042),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2039),
.B(n_1946),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2047),
.Y(n_2088)
);

HB1xp67_ASAP7_75t_L g2089 ( 
.A(n_2022),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_1992),
.B(n_1903),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2050),
.Y(n_2091)
);

INVx2_ASAP7_75t_SL g2092 ( 
.A(n_2013),
.Y(n_2092)
);

OR2x2_ASAP7_75t_L g2093 ( 
.A(n_2023),
.B(n_1951),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2012),
.B(n_1924),
.Y(n_2094)
);

BUFx12f_ASAP7_75t_L g2095 ( 
.A(n_1997),
.Y(n_2095)
);

HB1xp67_ASAP7_75t_L g2096 ( 
.A(n_2022),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_2025),
.B(n_1969),
.Y(n_2097)
);

OR2x2_ASAP7_75t_L g2098 ( 
.A(n_2040),
.B(n_1969),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2057),
.Y(n_2099)
);

INVx3_ASAP7_75t_L g2100 ( 
.A(n_2013),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2040),
.B(n_1969),
.Y(n_2101)
);

AND2x4_ASAP7_75t_L g2102 ( 
.A(n_2013),
.B(n_1888),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2058),
.B(n_1965),
.Y(n_2103)
);

BUFx3_ASAP7_75t_L g2104 ( 
.A(n_2029),
.Y(n_2104)
);

AND2x4_ASAP7_75t_L g2105 ( 
.A(n_2066),
.B(n_1888),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2012),
.B(n_1887),
.Y(n_2106)
);

INVx4_ASAP7_75t_L g2107 ( 
.A(n_2029),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2012),
.B(n_1976),
.Y(n_2108)
);

AOI21xp5_ASAP7_75t_L g2109 ( 
.A1(n_2011),
.A2(n_1989),
.B(n_1888),
.Y(n_2109)
);

BUFx2_ASAP7_75t_L g2110 ( 
.A(n_2061),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1993),
.Y(n_2111)
);

BUFx2_ASAP7_75t_L g2112 ( 
.A(n_2006),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2041),
.B(n_1963),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1995),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2044),
.B(n_1967),
.Y(n_2115)
);

INVxp67_ASAP7_75t_L g2116 ( 
.A(n_2051),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1996),
.Y(n_2117)
);

AND2x4_ASAP7_75t_L g2118 ( 
.A(n_2067),
.B(n_1888),
.Y(n_2118)
);

NOR2x1_ASAP7_75t_L g2119 ( 
.A(n_2055),
.B(n_1888),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2001),
.Y(n_2120)
);

AND2x4_ASAP7_75t_L g2121 ( 
.A(n_2067),
.B(n_1947),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2005),
.Y(n_2122)
);

NAND2xp33_ASAP7_75t_R g2123 ( 
.A(n_2027),
.B(n_1930),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2009),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2046),
.B(n_1885),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2015),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2017),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2006),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2056),
.Y(n_2129)
);

NOR2x1p5_ASAP7_75t_L g2130 ( 
.A(n_2003),
.B(n_1942),
.Y(n_2130)
);

INVxp67_ASAP7_75t_L g2131 ( 
.A(n_2103),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2115),
.B(n_2052),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2111),
.Y(n_2133)
);

BUFx3_ASAP7_75t_L g2134 ( 
.A(n_2095),
.Y(n_2134)
);

AOI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2130),
.A2(n_1998),
.B1(n_2000),
.B2(n_2030),
.Y(n_2135)
);

OAI33xp33_ASAP7_75t_L g2136 ( 
.A1(n_2103),
.A2(n_2028),
.A3(n_2049),
.B1(n_2064),
.B2(n_2045),
.B3(n_1905),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2100),
.B(n_2032),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_2090),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2115),
.B(n_2035),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2111),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2114),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2090),
.Y(n_2142)
);

OR2x2_ASAP7_75t_L g2143 ( 
.A(n_2071),
.B(n_2068),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_2071),
.B(n_2036),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2100),
.B(n_2075),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2114),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2114),
.Y(n_2147)
);

AOI21xp5_ASAP7_75t_L g2148 ( 
.A1(n_2109),
.A2(n_2011),
.B(n_2000),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2090),
.Y(n_2149)
);

INVxp67_ASAP7_75t_L g2150 ( 
.A(n_2130),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2100),
.B(n_2016),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2076),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2120),
.Y(n_2153)
);

OR2x2_ASAP7_75t_L g2154 ( 
.A(n_2097),
.B(n_2053),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2120),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2122),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2122),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2115),
.B(n_2059),
.Y(n_2158)
);

NOR2xp33_ASAP7_75t_SL g2159 ( 
.A(n_2107),
.B(n_2054),
.Y(n_2159)
);

OR2x2_ASAP7_75t_L g2160 ( 
.A(n_2097),
.B(n_2060),
.Y(n_2160)
);

HB1xp67_ASAP7_75t_L g2161 ( 
.A(n_2089),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2124),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2124),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2126),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2074),
.B(n_2065),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2126),
.Y(n_2166)
);

NOR2x1_ASAP7_75t_L g2167 ( 
.A(n_2119),
.B(n_2054),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2127),
.Y(n_2168)
);

INVx2_ASAP7_75t_SL g2169 ( 
.A(n_2095),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2127),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2117),
.Y(n_2171)
);

INVx2_ASAP7_75t_SL g2172 ( 
.A(n_2095),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2100),
.B(n_2008),
.Y(n_2173)
);

AO21x1_ASAP7_75t_L g2174 ( 
.A1(n_2123),
.A2(n_2004),
.B(n_2028),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2117),
.Y(n_2175)
);

OR2x2_ASAP7_75t_L g2176 ( 
.A(n_2097),
.B(n_1959),
.Y(n_2176)
);

NOR3xp33_ASAP7_75t_L g2177 ( 
.A(n_2109),
.B(n_1999),
.C(n_2049),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2117),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2077),
.Y(n_2179)
);

INVxp67_ASAP7_75t_SL g2180 ( 
.A(n_2116),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2077),
.Y(n_2181)
);

OR2x2_ASAP7_75t_L g2182 ( 
.A(n_2098),
.B(n_1959),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2080),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_SL g2184 ( 
.A(n_2119),
.B(n_2116),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2100),
.B(n_2008),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2080),
.Y(n_2186)
);

NAND3xp33_ASAP7_75t_L g2187 ( 
.A(n_2177),
.B(n_2034),
.C(n_2038),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2179),
.Y(n_2188)
);

NOR4xp25_ASAP7_75t_SL g2189 ( 
.A(n_2184),
.B(n_2004),
.C(n_2123),
.D(n_2110),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2145),
.B(n_2075),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2132),
.B(n_2043),
.Y(n_2191)
);

AND2x4_ASAP7_75t_L g2192 ( 
.A(n_2167),
.B(n_2180),
.Y(n_2192)
);

OR2x2_ASAP7_75t_L g2193 ( 
.A(n_2176),
.B(n_2108),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2133),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2152),
.Y(n_2195)
);

NAND2x1p5_ASAP7_75t_L g2196 ( 
.A(n_2184),
.B(n_2085),
.Y(n_2196)
);

AOI31xp33_ASAP7_75t_SL g2197 ( 
.A1(n_2148),
.A2(n_2150),
.A3(n_2165),
.B(n_2143),
.Y(n_2197)
);

HB1xp67_ASAP7_75t_L g2198 ( 
.A(n_2161),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2139),
.B(n_2034),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2140),
.Y(n_2200)
);

OAI31xp33_ASAP7_75t_L g2201 ( 
.A1(n_2143),
.A2(n_2108),
.A3(n_2064),
.B(n_2110),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2145),
.B(n_2075),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2158),
.B(n_2074),
.Y(n_2203)
);

OR2x2_ASAP7_75t_L g2204 ( 
.A(n_2176),
.B(n_2108),
.Y(n_2204)
);

AOI22xp5_ASAP7_75t_L g2205 ( 
.A1(n_2174),
.A2(n_2018),
.B1(n_2020),
.B2(n_2102),
.Y(n_2205)
);

AOI21xp33_ASAP7_75t_L g2206 ( 
.A1(n_2174),
.A2(n_2021),
.B(n_2072),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2151),
.B(n_2082),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2131),
.B(n_2074),
.Y(n_2208)
);

HB1xp67_ASAP7_75t_L g2209 ( 
.A(n_2144),
.Y(n_2209)
);

NAND2xp33_ASAP7_75t_SL g2210 ( 
.A(n_2169),
.B(n_2085),
.Y(n_2210)
);

INVx2_ASAP7_75t_SL g2211 ( 
.A(n_2134),
.Y(n_2211)
);

OR2x2_ASAP7_75t_L g2212 ( 
.A(n_2182),
.B(n_2098),
.Y(n_2212)
);

AOI222xp33_ASAP7_75t_L g2213 ( 
.A1(n_2136),
.A2(n_2062),
.B1(n_1930),
.B2(n_2002),
.C1(n_2007),
.C2(n_2094),
.Y(n_2213)
);

NAND2xp33_ASAP7_75t_SL g2214 ( 
.A(n_2169),
.B(n_2085),
.Y(n_2214)
);

OR2x4_ASAP7_75t_L g2215 ( 
.A(n_2144),
.B(n_2072),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2152),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2151),
.B(n_2082),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2179),
.Y(n_2218)
);

HB1xp67_ASAP7_75t_L g2219 ( 
.A(n_2153),
.Y(n_2219)
);

AND2x2_ASAP7_75t_SL g2220 ( 
.A(n_2135),
.B(n_2110),
.Y(n_2220)
);

OR2x2_ASAP7_75t_L g2221 ( 
.A(n_2182),
.B(n_2098),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2173),
.B(n_2082),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2173),
.B(n_2185),
.Y(n_2223)
);

NOR2xp33_ASAP7_75t_SL g2224 ( 
.A(n_2159),
.B(n_2107),
.Y(n_2224)
);

NAND2xp33_ASAP7_75t_SL g2225 ( 
.A(n_2172),
.B(n_2107),
.Y(n_2225)
);

OAI22xp33_ASAP7_75t_L g2226 ( 
.A1(n_2172),
.A2(n_2107),
.B1(n_2104),
.B2(n_2019),
.Y(n_2226)
);

BUFx3_ASAP7_75t_L g2227 ( 
.A(n_2134),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2186),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2155),
.B(n_2073),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_L g2230 ( 
.A(n_2185),
.B(n_1991),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2186),
.Y(n_2231)
);

CKINVDCx16_ASAP7_75t_R g2232 ( 
.A(n_2137),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2137),
.B(n_2078),
.Y(n_2233)
);

HB1xp67_ASAP7_75t_L g2234 ( 
.A(n_2156),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2157),
.B(n_2073),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2141),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2154),
.B(n_2078),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2162),
.B(n_2073),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2163),
.B(n_2113),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2164),
.B(n_2113),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_R g2241 ( 
.A(n_2154),
.B(n_2104),
.Y(n_2241)
);

OAI22xp33_ASAP7_75t_L g2242 ( 
.A1(n_2205),
.A2(n_2107),
.B1(n_2104),
.B2(n_2112),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2227),
.Y(n_2243)
);

NAND2xp33_ASAP7_75t_SL g2244 ( 
.A(n_2189),
.B(n_2094),
.Y(n_2244)
);

OR2x6_ASAP7_75t_L g2245 ( 
.A(n_2211),
.B(n_2104),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2188),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2191),
.B(n_2166),
.Y(n_2247)
);

AOI322xp5_ASAP7_75t_L g2248 ( 
.A1(n_2220),
.A2(n_2094),
.A3(n_2106),
.B1(n_2112),
.B2(n_2078),
.C1(n_2083),
.C2(n_2079),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2227),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2213),
.B(n_2168),
.Y(n_2250)
);

OAI211xp5_ASAP7_75t_SL g2251 ( 
.A1(n_2201),
.A2(n_2149),
.B(n_2142),
.C(n_2138),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_2223),
.Y(n_2252)
);

OA21x2_ASAP7_75t_L g2253 ( 
.A1(n_2206),
.A2(n_2142),
.B(n_2149),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2188),
.Y(n_2254)
);

OR2x2_ASAP7_75t_L g2255 ( 
.A(n_2203),
.B(n_2209),
.Y(n_2255)
);

AOI22xp5_ASAP7_75t_L g2256 ( 
.A1(n_2220),
.A2(n_2106),
.B1(n_2018),
.B2(n_2083),
.Y(n_2256)
);

AOI211xp5_ASAP7_75t_L g2257 ( 
.A1(n_2197),
.A2(n_2112),
.B(n_2010),
.C(n_2128),
.Y(n_2257)
);

AOI221xp5_ASAP7_75t_L g2258 ( 
.A1(n_2187),
.A2(n_2138),
.B1(n_2128),
.B2(n_2170),
.C(n_2106),
.Y(n_2258)
);

AO32x1_ASAP7_75t_L g2259 ( 
.A1(n_2211),
.A2(n_2223),
.A3(n_2092),
.B1(n_2217),
.B2(n_2222),
.Y(n_2259)
);

OR2x2_ASAP7_75t_L g2260 ( 
.A(n_2208),
.B(n_2160),
.Y(n_2260)
);

INVx1_ASAP7_75t_SL g2261 ( 
.A(n_2210),
.Y(n_2261)
);

OAI221xp5_ASAP7_75t_L g2262 ( 
.A1(n_2210),
.A2(n_2014),
.B1(n_2128),
.B2(n_2083),
.C(n_2079),
.Y(n_2262)
);

INVxp67_ASAP7_75t_L g2263 ( 
.A(n_2214),
.Y(n_2263)
);

AOI21xp5_ASAP7_75t_L g2264 ( 
.A1(n_2214),
.A2(n_2072),
.B(n_2079),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2218),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2232),
.B(n_2092),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2207),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2218),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2228),
.Y(n_2269)
);

NOR2xp67_ASAP7_75t_L g2270 ( 
.A(n_2192),
.B(n_2198),
.Y(n_2270)
);

OAI22xp5_ASAP7_75t_L g2271 ( 
.A1(n_2196),
.A2(n_2014),
.B1(n_2092),
.B2(n_2160),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2207),
.B(n_2102),
.Y(n_2272)
);

A2O1A1Ixp33_ASAP7_75t_L g2273 ( 
.A1(n_2192),
.A2(n_2118),
.B(n_2102),
.C(n_2016),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2199),
.B(n_2181),
.Y(n_2274)
);

INVxp67_ASAP7_75t_L g2275 ( 
.A(n_2192),
.Y(n_2275)
);

OAI21xp33_ASAP7_75t_L g2276 ( 
.A1(n_2196),
.A2(n_2118),
.B(n_2129),
.Y(n_2276)
);

OAI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2196),
.A2(n_1908),
.B1(n_2089),
.B2(n_2096),
.Y(n_2277)
);

OAI322xp33_ASAP7_75t_L g2278 ( 
.A1(n_2193),
.A2(n_2101),
.A3(n_2183),
.B1(n_2141),
.B2(n_2178),
.C1(n_2147),
.C2(n_2146),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2228),
.Y(n_2279)
);

OAI32xp33_ASAP7_75t_L g2280 ( 
.A1(n_2225),
.A2(n_2096),
.A3(n_2101),
.B1(n_2178),
.B2(n_2147),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2231),
.Y(n_2281)
);

AOI31xp33_ASAP7_75t_L g2282 ( 
.A1(n_2225),
.A2(n_2118),
.A3(n_2102),
.B(n_1940),
.Y(n_2282)
);

NAND2x1p5_ASAP7_75t_L g2283 ( 
.A(n_2217),
.B(n_2102),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2231),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2275),
.B(n_2243),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2283),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2246),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2266),
.B(n_2222),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2249),
.B(n_2230),
.Y(n_2289)
);

NOR2xp67_ASAP7_75t_L g2290 ( 
.A(n_2270),
.B(n_2219),
.Y(n_2290)
);

AOI222xp33_ASAP7_75t_L g2291 ( 
.A1(n_2250),
.A2(n_2226),
.B1(n_2224),
.B2(n_2234),
.C1(n_2237),
.C2(n_2200),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2247),
.B(n_2194),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_2283),
.Y(n_2293)
);

OAI22xp33_ASAP7_75t_L g2294 ( 
.A1(n_2256),
.A2(n_2215),
.B1(n_2193),
.B2(n_2204),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2254),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2265),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2268),
.Y(n_2297)
);

AND2x4_ASAP7_75t_L g2298 ( 
.A(n_2245),
.B(n_2190),
.Y(n_2298)
);

AOI22xp33_ASAP7_75t_L g2299 ( 
.A1(n_2244),
.A2(n_2241),
.B1(n_2118),
.B2(n_2237),
.Y(n_2299)
);

INVxp67_ASAP7_75t_SL g2300 ( 
.A(n_2263),
.Y(n_2300)
);

HB1xp67_ASAP7_75t_L g2301 ( 
.A(n_2252),
.Y(n_2301)
);

INVxp67_ASAP7_75t_L g2302 ( 
.A(n_2261),
.Y(n_2302)
);

OAI221xp5_ASAP7_75t_L g2303 ( 
.A1(n_2257),
.A2(n_2204),
.B1(n_2239),
.B2(n_2240),
.C(n_2221),
.Y(n_2303)
);

OAI21xp5_ASAP7_75t_L g2304 ( 
.A1(n_2242),
.A2(n_2195),
.B(n_2216),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2269),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2279),
.Y(n_2306)
);

NOR4xp25_ASAP7_75t_SL g2307 ( 
.A(n_2251),
.B(n_2215),
.C(n_2146),
.D(n_2171),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2281),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2245),
.Y(n_2309)
);

AOI22xp5_ASAP7_75t_L g2310 ( 
.A1(n_2258),
.A2(n_2215),
.B1(n_2118),
.B2(n_2202),
.Y(n_2310)
);

OAI22xp33_ASAP7_75t_L g2311 ( 
.A1(n_2261),
.A2(n_2238),
.B1(n_2229),
.B2(n_2235),
.Y(n_2311)
);

INVx2_ASAP7_75t_SL g2312 ( 
.A(n_2245),
.Y(n_2312)
);

OAI21xp5_ASAP7_75t_L g2313 ( 
.A1(n_2271),
.A2(n_2195),
.B(n_2216),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2284),
.Y(n_2314)
);

XOR2x2_ASAP7_75t_L g2315 ( 
.A(n_2290),
.B(n_2271),
.Y(n_2315)
);

INVx1_ASAP7_75t_SL g2316 ( 
.A(n_2288),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_2291),
.B(n_2277),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2300),
.B(n_2247),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2301),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2287),
.Y(n_2320)
);

INVx1_ASAP7_75t_SL g2321 ( 
.A(n_2288),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2287),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2298),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2302),
.B(n_2274),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2295),
.Y(n_2325)
);

NAND2xp33_ASAP7_75t_SL g2326 ( 
.A(n_2307),
.B(n_2277),
.Y(n_2326)
);

NOR3xp33_ASAP7_75t_SL g2327 ( 
.A(n_2285),
.B(n_2262),
.C(n_2273),
.Y(n_2327)
);

XOR2xp5_ASAP7_75t_L g2328 ( 
.A(n_2289),
.B(n_2255),
.Y(n_2328)
);

INVx1_ASAP7_75t_SL g2329 ( 
.A(n_2312),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2309),
.B(n_2274),
.Y(n_2330)
);

NOR3x1_ASAP7_75t_L g2331 ( 
.A(n_2312),
.B(n_2260),
.C(n_2259),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2295),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2296),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2298),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2296),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2297),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2297),
.Y(n_2337)
);

AOI22xp33_ASAP7_75t_L g2338 ( 
.A1(n_2294),
.A2(n_2299),
.B1(n_2310),
.B2(n_2267),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2319),
.Y(n_2339)
);

NOR3x1_ASAP7_75t_L g2340 ( 
.A(n_2317),
.B(n_2313),
.C(n_2292),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2316),
.B(n_2309),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2321),
.B(n_2298),
.Y(n_2342)
);

OAI21xp5_ASAP7_75t_L g2343 ( 
.A1(n_2317),
.A2(n_2311),
.B(n_2304),
.Y(n_2343)
);

AOI21xp5_ASAP7_75t_L g2344 ( 
.A1(n_2326),
.A2(n_2259),
.B(n_2253),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_2326),
.B(n_2282),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2319),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2329),
.B(n_2286),
.Y(n_2347)
);

AOI21xp5_ASAP7_75t_L g2348 ( 
.A1(n_2315),
.A2(n_2259),
.B(n_2253),
.Y(n_2348)
);

OR3x1_ASAP7_75t_L g2349 ( 
.A(n_2322),
.B(n_2280),
.C(n_2308),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2323),
.B(n_2305),
.Y(n_2350)
);

NAND4xp25_ASAP7_75t_L g2351 ( 
.A(n_2331),
.B(n_2248),
.C(n_2303),
.D(n_2306),
.Y(n_2351)
);

NOR2x1_ASAP7_75t_L g2352 ( 
.A(n_2320),
.B(n_2305),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2323),
.B(n_2306),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2342),
.B(n_2328),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2347),
.B(n_2328),
.Y(n_2355)
);

OAI211xp5_ASAP7_75t_L g2356 ( 
.A1(n_2345),
.A2(n_2338),
.B(n_2327),
.C(n_2318),
.Y(n_2356)
);

AOI221xp5_ASAP7_75t_L g2357 ( 
.A1(n_2343),
.A2(n_2324),
.B1(n_2330),
.B2(n_2334),
.C(n_2335),
.Y(n_2357)
);

AOI322xp5_ASAP7_75t_L g2358 ( 
.A1(n_2352),
.A2(n_2337),
.A3(n_2336),
.B1(n_2325),
.B2(n_2333),
.C1(n_2332),
.C2(n_2276),
.Y(n_2358)
);

AOI221x1_ASAP7_75t_L g2359 ( 
.A1(n_2344),
.A2(n_2348),
.B1(n_2339),
.B2(n_2346),
.C(n_2351),
.Y(n_2359)
);

OAI221xp5_ASAP7_75t_L g2360 ( 
.A1(n_2351),
.A2(n_2315),
.B1(n_2334),
.B2(n_2286),
.C(n_2293),
.Y(n_2360)
);

OAI21xp5_ASAP7_75t_L g2361 ( 
.A1(n_2341),
.A2(n_2282),
.B(n_2264),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2340),
.B(n_2350),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2353),
.Y(n_2363)
);

XNOR2xp5_ASAP7_75t_L g2364 ( 
.A(n_2349),
.B(n_2293),
.Y(n_2364)
);

NAND5xp2_ASAP7_75t_L g2365 ( 
.A(n_2343),
.B(n_2320),
.C(n_2314),
.D(n_2308),
.E(n_2272),
.Y(n_2365)
);

AOI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2345),
.A2(n_2314),
.B(n_2278),
.Y(n_2366)
);

O2A1O1Ixp33_ASAP7_75t_L g2367 ( 
.A1(n_2345),
.A2(n_2221),
.B(n_2212),
.C(n_2236),
.Y(n_2367)
);

NOR2xp33_ASAP7_75t_R g2368 ( 
.A(n_2354),
.B(n_2355),
.Y(n_2368)
);

AND2x4_ASAP7_75t_L g2369 ( 
.A(n_2359),
.B(n_2190),
.Y(n_2369)
);

NAND3xp33_ASAP7_75t_L g2370 ( 
.A(n_2356),
.B(n_2236),
.C(n_2212),
.Y(n_2370)
);

AOI322xp5_ASAP7_75t_L g2371 ( 
.A1(n_2362),
.A2(n_2233),
.A3(n_2202),
.B1(n_2113),
.B2(n_2070),
.C1(n_2125),
.C2(n_2129),
.Y(n_2371)
);

AOI22xp5_ASAP7_75t_L g2372 ( 
.A1(n_2364),
.A2(n_2233),
.B1(n_2121),
.B2(n_1952),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_SL g2373 ( 
.A(n_2361),
.B(n_2121),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2363),
.Y(n_2374)
);

NOR3x1_ASAP7_75t_L g2375 ( 
.A(n_2360),
.B(n_2101),
.C(n_2175),
.Y(n_2375)
);

OR2x2_ASAP7_75t_L g2376 ( 
.A(n_2365),
.B(n_2081),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2369),
.B(n_2357),
.Y(n_2377)
);

HB1xp67_ASAP7_75t_L g2378 ( 
.A(n_2368),
.Y(n_2378)
);

NAND4xp75_ASAP7_75t_L g2379 ( 
.A(n_2375),
.B(n_2366),
.C(n_2358),
.D(n_2367),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2376),
.B(n_2087),
.Y(n_2380)
);

AND3x4_ASAP7_75t_L g2381 ( 
.A(n_2372),
.B(n_2105),
.C(n_2121),
.Y(n_2381)
);

AND2x4_ASAP7_75t_L g2382 ( 
.A(n_2374),
.B(n_2087),
.Y(n_2382)
);

AOI21xp5_ASAP7_75t_L g2383 ( 
.A1(n_2373),
.A2(n_2121),
.B(n_1926),
.Y(n_2383)
);

OAI321xp33_ASAP7_75t_L g2384 ( 
.A1(n_2370),
.A2(n_2371),
.A3(n_1935),
.B1(n_1942),
.B2(n_1940),
.C(n_1961),
.Y(n_2384)
);

HB1xp67_ASAP7_75t_L g2385 ( 
.A(n_2369),
.Y(n_2385)
);

NAND4xp25_ASAP7_75t_L g2386 ( 
.A(n_2377),
.B(n_2105),
.C(n_2081),
.D(n_2121),
.Y(n_2386)
);

NOR2x1_ASAP7_75t_L g2387 ( 
.A(n_2379),
.B(n_2091),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2385),
.B(n_2099),
.Y(n_2388)
);

OA22x2_ASAP7_75t_L g2389 ( 
.A1(n_2381),
.A2(n_2125),
.B1(n_1952),
.B2(n_1961),
.Y(n_2389)
);

OAI221xp5_ASAP7_75t_SL g2390 ( 
.A1(n_2380),
.A2(n_2093),
.B1(n_2125),
.B2(n_2087),
.C(n_2070),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2378),
.Y(n_2391)
);

OAI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_2384),
.A2(n_2088),
.B(n_2086),
.Y(n_2392)
);

XNOR2xp5_ASAP7_75t_L g2393 ( 
.A(n_2391),
.B(n_2382),
.Y(n_2393)
);

NOR3xp33_ASAP7_75t_L g2394 ( 
.A(n_2387),
.B(n_2383),
.C(n_1977),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2389),
.Y(n_2395)
);

CKINVDCx5p33_ASAP7_75t_R g2396 ( 
.A(n_2388),
.Y(n_2396)
);

AND2x4_ASAP7_75t_L g2397 ( 
.A(n_2395),
.B(n_2392),
.Y(n_2397)
);

AND2x4_ASAP7_75t_L g2398 ( 
.A(n_2396),
.B(n_2386),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_SL g2399 ( 
.A(n_2397),
.B(n_2394),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2399),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2399),
.Y(n_2401)
);

NAND3xp33_ASAP7_75t_L g2402 ( 
.A(n_2400),
.B(n_2393),
.C(n_2397),
.Y(n_2402)
);

INVxp67_ASAP7_75t_L g2403 ( 
.A(n_2401),
.Y(n_2403)
);

AOI22xp33_ASAP7_75t_L g2404 ( 
.A1(n_2402),
.A2(n_2398),
.B1(n_2403),
.B2(n_2390),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2402),
.Y(n_2405)
);

NAND3xp33_ASAP7_75t_R g2406 ( 
.A(n_2404),
.B(n_1968),
.C(n_1952),
.Y(n_2406)
);

OAI221xp5_ASAP7_75t_R g2407 ( 
.A1(n_2406),
.A2(n_2405),
.B1(n_1908),
.B2(n_1968),
.C(n_2029),
.Y(n_2407)
);

AOI211xp5_ASAP7_75t_L g2408 ( 
.A1(n_2407),
.A2(n_2088),
.B(n_2084),
.C(n_2086),
.Y(n_2408)
);


endmodule