module fake_jpeg_7329_n_228 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_SL g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_33),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_1),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_1),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_45),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_17),
.B1(n_21),
.B2(n_31),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_49),
.B1(n_18),
.B2(n_19),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_2),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_31),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_16),
.C(n_23),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_17),
.B1(n_21),
.B2(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVxp67_ASAP7_75t_SL g84 ( 
.A(n_55),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_33),
.B1(n_32),
.B2(n_21),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_56),
.A2(n_62),
.B1(n_66),
.B2(n_27),
.Y(n_82)
);

OAI22x1_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_37),
.B1(n_34),
.B2(n_17),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_75),
.B1(n_79),
.B2(n_22),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_58),
.B(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_45),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_23),
.B(n_26),
.C(n_25),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_19),
.B1(n_34),
.B2(n_16),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_2),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_19),
.B1(n_34),
.B2(n_28),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_78),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_25),
.B1(n_22),
.B2(n_30),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

CKINVDCx12_ASAP7_75t_R g85 ( 
.A(n_77),
.Y(n_85)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_26),
.B1(n_28),
.B2(n_27),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_40),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_87),
.B1(n_88),
.B2(n_73),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_39),
.B1(n_38),
.B2(n_25),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_77),
.B1(n_64),
.B2(n_55),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_90),
.B(n_5),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_3),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_56),
.C(n_65),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_59),
.C(n_72),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_4),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_4),
.B(n_5),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_81),
.B(n_43),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_127),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_75),
.C(n_43),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_122),
.C(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_117),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_109),
.B(n_123),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_61),
.B(n_62),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_112),
.B(n_125),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_76),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_116),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_89),
.A2(n_66),
.B1(n_67),
.B2(n_54),
.Y(n_115)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_74),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_40),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_74),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_120),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_102),
.B1(n_100),
.B2(n_8),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_81),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_82),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_100),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_30),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

NAND2x1_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_4),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_14),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_128),
.B(n_103),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_99),
.B(n_91),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_138),
.B(n_145),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_114),
.A2(n_91),
.B1(n_103),
.B2(n_101),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_111),
.A2(n_90),
.B(n_95),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_151),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_87),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_146),
.C(n_147),
.Y(n_153)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_86),
.C(n_101),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_104),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_102),
.B(n_104),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_152),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_115),
.B1(n_105),
.B2(n_127),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_107),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_108),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_169),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_143),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_108),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_161),
.Y(n_172)
);

A2O1A1O1Ixp25_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_106),
.B(n_125),
.C(n_117),
.D(n_109),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_164),
.B(n_135),
.Y(n_180)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_166),
.A2(n_136),
.B1(n_148),
.B2(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_14),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_134),
.A2(n_106),
.B1(n_7),
.B2(n_8),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_170),
.A2(n_129),
.B1(n_136),
.B2(n_134),
.Y(n_173)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_6),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_173),
.B(n_179),
.Y(n_197)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_163),
.A2(n_131),
.B1(n_151),
.B2(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_154),
.A2(n_140),
.B1(n_142),
.B2(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_155),
.A2(n_146),
.B1(n_150),
.B2(n_147),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_170),
.C(n_166),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_153),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_155),
.A2(n_150),
.B1(n_132),
.B2(n_129),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_183),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_132),
.B(n_150),
.Y(n_183)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_185),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_153),
.C(n_159),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_195),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_191),
.C(n_194),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_164),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g206 ( 
.A(n_193),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_157),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_160),
.C(n_162),
.Y(n_195)
);

XOR2x1_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_182),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_SL g209 ( 
.A1(n_198),
.A2(n_172),
.B(n_171),
.Y(n_209)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_203),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_183),
.C(n_163),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_205),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_187),
.A2(n_173),
.B1(n_184),
.B2(n_176),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_190),
.B1(n_160),
.B2(n_196),
.Y(n_208)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_186),
.C(n_188),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_210),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_175),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_202),
.A2(n_175),
.B(n_185),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_213),
.B(n_9),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_215),
.A2(n_212),
.B(n_209),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_7),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_218),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_221),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_217),
.B(n_9),
.Y(n_221)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_214),
.A3(n_217),
.B1(n_222),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_11),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_224),
.C(n_11),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_12),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_12),
.Y(n_228)
);


endmodule