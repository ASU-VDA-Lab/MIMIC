module fake_netlist_6_4118_n_1538 (n_41, n_16, n_1, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_27, n_3, n_14, n_38, n_0, n_39, n_32, n_4, n_36, n_22, n_26, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_43, n_5, n_19, n_29, n_31, n_25, n_40, n_44, n_1538);

input n_41;
input n_16;
input n_1;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_39;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_43;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;
input n_40;
input n_44;

output n_1538;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_68;
wire n_726;
wire n_212;
wire n_700;
wire n_50;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_77;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_78;
wire n_1380;
wire n_442;
wire n_480;
wire n_142;
wire n_1402;
wire n_1009;
wire n_62;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_65;
wire n_230;
wire n_461;
wire n_873;
wire n_141;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_71;
wire n_229;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_45;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_112;
wire n_1280;
wire n_713;
wire n_1400;
wire n_126;
wire n_1467;
wire n_58;
wire n_976;
wire n_224;
wire n_48;
wire n_1445;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_92;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_102;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_121;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_61;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_117;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_134;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_136;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_88;
wire n_530;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_47;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_55;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_91;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_63;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_125;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_131;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_59;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_108;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_86;
wire n_104;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_72;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_79;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_145;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_118;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_107;
wire n_1228;
wire n_417;
wire n_446;
wire n_89;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_69;
wire n_293;
wire n_53;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_98;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_66;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_100;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_124;
wire n_1382;
wire n_1534;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_123;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1136;
wire n_128;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_146;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_113;
wire n_1533;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_90;
wire n_54;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_99;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_120;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_144;
wire n_1203;
wire n_820;
wire n_951;
wire n_106;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_140;
wire n_1138;
wire n_1275;
wire n_485;
wire n_67;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_73;
wire n_785;
wire n_746;
wire n_609;
wire n_101;
wire n_167;
wire n_1356;
wire n_127;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_133;
wire n_1320;
wire n_96;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_302;
wire n_380;
wire n_1535;
wire n_137;
wire n_1190;
wire n_397;
wire n_122;
wire n_1262;
wire n_218;
wire n_1213;
wire n_70;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_97;
wire n_782;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_80;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_83;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_105;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_76;
wire n_548;
wire n_94;
wire n_282;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_139;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_138;
wire n_1498;
wire n_1210;
wire n_49;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_85;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_75;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_110;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_57;
wire n_1007;
wire n_1378;
wire n_855;
wire n_52;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_84;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_143;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_114;
wire n_300;
wire n_222;
wire n_747;
wire n_74;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_111;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_56;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_119;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_129;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_109;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_82;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_93;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_366;
wire n_1509;
wire n_103;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_46;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_132;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_130;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_116;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_95;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_115;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_87;
wire n_257;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_81;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_64;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_135;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_60;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_51;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_19),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_13),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_0),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_13),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_21),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_18),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_11),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_15),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_11),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_21),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_2),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_31),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_1),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_86),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVxp33_ASAP7_75t_SL g94 ( 
.A(n_48),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

BUFx2_ASAP7_75t_SL g97 ( 
.A(n_71),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_51),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_53),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_55),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_60),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_83),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_83),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_88),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_88),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_88),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_73),
.B1(n_84),
.B2(n_57),
.Y(n_122)
);

OAI21x1_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_71),
.B(n_88),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

AND2x4_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_85),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_58),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_112),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_96),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_109),
.B(n_106),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_90),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_96),
.Y(n_143)
);

BUFx10_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_96),
.B(n_94),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_108),
.A2(n_127),
.B1(n_126),
.B2(n_118),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_85),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_112),
.B(n_106),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_112),
.B(n_104),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_126),
.B(n_64),
.Y(n_157)
);

OR2x6_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_64),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_58),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_116),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_116),
.A2(n_82),
.B1(n_69),
.B2(n_77),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_112),
.B(n_104),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_SL g173 ( 
.A(n_113),
.B(n_66),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

OR2x6_ASAP7_75t_L g175 ( 
.A(n_123),
.B(n_74),
.Y(n_175)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_123),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_112),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_126),
.B(n_100),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_130),
.Y(n_181)
);

NOR3xp33_ASAP7_75t_L g182 ( 
.A(n_113),
.B(n_107),
.C(n_78),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

CKINVDCx11_ASAP7_75t_R g186 ( 
.A(n_113),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_117),
.B(n_74),
.C(n_62),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_122),
.A2(n_56),
.B1(n_65),
.B2(n_92),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_110),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_122),
.A2(n_102),
.B1(n_92),
.B2(n_107),
.Y(n_193)
);

OR2x6_ASAP7_75t_L g194 ( 
.A(n_126),
.B(n_70),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_128),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_136),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_136),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_141),
.B(n_126),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_141),
.B(n_117),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_137),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_188),
.A2(n_98),
.B1(n_100),
.B2(n_94),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_150),
.A2(n_119),
.B1(n_118),
.B2(n_130),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_141),
.B(n_119),
.Y(n_203)
);

NAND2xp33_ASAP7_75t_L g204 ( 
.A(n_146),
.B(n_120),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_150),
.B(n_144),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_150),
.B(n_120),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_149),
.B(n_131),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_149),
.B(n_139),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_139),
.B(n_131),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_140),
.B(n_121),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_L g216 ( 
.A(n_146),
.B(n_121),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_144),
.B(n_115),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_143),
.B(n_131),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_143),
.B(n_131),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_157),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_166),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_140),
.B(n_115),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_144),
.B(n_115),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g226 ( 
.A(n_177),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_144),
.B(n_45),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_157),
.B(n_131),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_173),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_180),
.B(n_99),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_152),
.A2(n_58),
.B1(n_87),
.B2(n_47),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_144),
.B(n_80),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_174),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_157),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_162),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_146),
.B(n_46),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_157),
.B(n_131),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_152),
.B(n_131),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_160),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_146),
.B(n_75),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_146),
.B(n_68),
.Y(n_246)
);

NOR2xp67_ASAP7_75t_L g247 ( 
.A(n_138),
.B(n_32),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_160),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_193),
.B(n_56),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_195),
.Y(n_250)
);

NOR2xp67_ASAP7_75t_L g251 ( 
.A(n_138),
.B(n_39),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_152),
.B(n_131),
.Y(n_252)
);

AND2x4_ASAP7_75t_L g253 ( 
.A(n_194),
.B(n_81),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_195),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_180),
.B(n_99),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_152),
.A2(n_158),
.B1(n_146),
.B2(n_194),
.Y(n_256)
);

INVxp67_ASAP7_75t_SL g257 ( 
.A(n_177),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_152),
.B(n_131),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_163),
.B(n_61),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_177),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_152),
.B(n_125),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_158),
.B(n_102),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_146),
.A2(n_176),
.B(n_170),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_152),
.B(n_125),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_147),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_158),
.B(n_102),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_163),
.B(n_67),
.Y(n_267)
);

AOI221xp5_ASAP7_75t_L g268 ( 
.A1(n_193),
.A2(n_107),
.B1(n_52),
.B2(n_89),
.C(n_81),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_159),
.B(n_56),
.Y(n_270)
);

NAND2xp33_ASAP7_75t_L g271 ( 
.A(n_138),
.B(n_58),
.Y(n_271)
);

AND2x2_ASAP7_75t_SL g272 ( 
.A(n_177),
.B(n_62),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_152),
.B(n_125),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_177),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_177),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_182),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_152),
.B(n_125),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_182),
.B(n_62),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_177),
.Y(n_279)
);

NAND3xp33_ASAP7_75t_L g280 ( 
.A(n_158),
.B(n_68),
.C(n_62),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_152),
.B(n_125),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_183),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_L g283 ( 
.A(n_142),
.B(n_135),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_142),
.B(n_62),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_176),
.Y(n_285)
);

INVxp33_ASAP7_75t_L g286 ( 
.A(n_186),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_147),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_158),
.A2(n_70),
.B1(n_52),
.B2(n_72),
.Y(n_288)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_209),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_220),
.B(n_183),
.Y(n_290)
);

AND2x4_ASAP7_75t_L g291 ( 
.A(n_198),
.B(n_158),
.Y(n_291)
);

NAND2x1p5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_183),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_214),
.B(n_159),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_199),
.B(n_183),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_200),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_203),
.B(n_183),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_244),
.B(n_183),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_240),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_196),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_244),
.B(n_183),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_248),
.B(n_148),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_269),
.Y(n_303)
);

AND2x6_ASAP7_75t_SL g304 ( 
.A(n_259),
.B(n_54),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_226),
.A2(n_176),
.B(n_142),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_240),
.Y(n_306)
);

AND2x4_ASAP7_75t_L g307 ( 
.A(n_198),
.B(n_194),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_196),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_275),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_253),
.B(n_194),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_220),
.A2(n_153),
.B1(n_156),
.B2(n_165),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_222),
.B(n_153),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_248),
.B(n_148),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_238),
.B(n_172),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_205),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_238),
.B(n_172),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_232),
.B(n_172),
.Y(n_317)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_209),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_267),
.A2(n_194),
.B1(n_188),
.B2(n_165),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_255),
.B(n_170),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_200),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_211),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_205),
.Y(n_323)
);

BUFx8_ASAP7_75t_L g324 ( 
.A(n_262),
.Y(n_324)
);

AND2x6_ASAP7_75t_L g325 ( 
.A(n_275),
.B(n_170),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_210),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_212),
.B(n_179),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_257),
.B(n_179),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_202),
.B(n_179),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_202),
.B(n_184),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_200),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_210),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_223),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_276),
.B(n_156),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_262),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_215),
.Y(n_336)
);

BUFx4f_ASAP7_75t_L g337 ( 
.A(n_253),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_223),
.Y(n_338)
);

OR2x2_ASAP7_75t_SL g339 ( 
.A(n_249),
.B(n_186),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_266),
.Y(n_340)
);

AO22x1_ASAP7_75t_L g341 ( 
.A1(n_270),
.A2(n_79),
.B1(n_54),
.B2(n_59),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_227),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_201),
.Y(n_343)
);

AOI22x1_ASAP7_75t_L g344 ( 
.A1(n_215),
.A2(n_189),
.B1(n_184),
.B2(n_190),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_215),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_227),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_272),
.B(n_184),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_221),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_221),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_272),
.B(n_189),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_266),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_272),
.B(n_189),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_253),
.A2(n_194),
.B1(n_176),
.B2(n_187),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_224),
.B(n_194),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_229),
.B(n_190),
.Y(n_355)
);

BUFx8_ASAP7_75t_L g356 ( 
.A(n_224),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_207),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_253),
.A2(n_206),
.B1(n_208),
.B2(n_278),
.Y(n_358)
);

NOR2xp67_ASAP7_75t_L g359 ( 
.A(n_231),
.B(n_187),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_229),
.B(n_190),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_235),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_217),
.A2(n_230),
.B1(n_242),
.B2(n_234),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_221),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_288),
.B(n_175),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_225),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_288),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_235),
.Y(n_367)
);

OR2x6_ASAP7_75t_L g368 ( 
.A(n_260),
.B(n_176),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_237),
.B(n_191),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_209),
.B(n_178),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_260),
.B(n_274),
.Y(n_371)
);

A2O1A1Ixp33_ASAP7_75t_SL g372 ( 
.A1(n_197),
.A2(n_145),
.B(n_191),
.C(n_185),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_201),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_237),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_312),
.B(n_260),
.Y(n_375)
);

AO32x2_ASAP7_75t_L g376 ( 
.A1(n_321),
.A2(n_178),
.A3(n_268),
.B1(n_225),
.B2(n_197),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_312),
.A2(n_319),
.B1(n_362),
.B2(n_311),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_293),
.B(n_274),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_293),
.A2(n_334),
.B1(n_291),
.B2(n_335),
.Y(n_379)
);

BUFx5_ASAP7_75t_L g380 ( 
.A(n_325),
.Y(n_380)
);

BUFx8_ASAP7_75t_L g381 ( 
.A(n_306),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_310),
.B(n_274),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_318),
.B(n_209),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_298),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_340),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_363),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_318),
.A2(n_285),
.B(n_178),
.Y(n_387)
);

O2A1O1Ixp33_ASAP7_75t_L g388 ( 
.A1(n_334),
.A2(n_236),
.B(n_225),
.C(n_228),
.Y(n_388)
);

A2O1A1Ixp33_ASAP7_75t_L g389 ( 
.A1(n_302),
.A2(n_233),
.B(n_247),
.C(n_251),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_374),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_300),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_SL g392 ( 
.A(n_318),
.B(n_300),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_297),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_318),
.A2(n_285),
.B(n_289),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_363),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_351),
.B(n_279),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_318),
.A2(n_285),
.B(n_283),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_300),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_299),
.Y(n_399)
);

A2O1A1Ixp33_ASAP7_75t_SL g400 ( 
.A1(n_358),
.A2(n_271),
.B(n_275),
.C(n_236),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_R g401 ( 
.A(n_298),
.B(n_204),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_294),
.B(n_279),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_289),
.A2(n_285),
.B(n_296),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_306),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_322),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_363),
.Y(n_406)
);

AOI33xp33_ASAP7_75t_L g407 ( 
.A1(n_357),
.A2(n_89),
.A3(n_79),
.B1(n_72),
.B2(n_59),
.B3(n_76),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_295),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_313),
.A2(n_256),
.B1(n_275),
.B2(n_279),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_291),
.B(n_282),
.Y(n_410)
);

O2A1O1Ixp33_ASAP7_75t_L g411 ( 
.A1(n_317),
.A2(n_216),
.B(n_284),
.C(n_219),
.Y(n_411)
);

A2O1A1Ixp33_ASAP7_75t_L g412 ( 
.A1(n_359),
.A2(n_233),
.B(n_251),
.C(n_247),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_366),
.B(n_282),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_343),
.B(n_282),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_301),
.B(n_213),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_308),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_315),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_291),
.B(n_243),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_289),
.A2(n_283),
.B(n_218),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_300),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_307),
.Y(n_421)
);

AO32x1_ASAP7_75t_L g422 ( 
.A1(n_321),
.A2(n_76),
.A3(n_250),
.B1(n_265),
.B2(n_254),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_323),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_307),
.A2(n_241),
.B1(n_245),
.B2(n_281),
.Y(n_424)
);

A2O1A1Ixp33_ASAP7_75t_L g425 ( 
.A1(n_364),
.A2(n_280),
.B(n_263),
.C(n_252),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_326),
.B(n_332),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_328),
.A2(n_246),
.B(n_277),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_305),
.A2(n_258),
.B(n_273),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_333),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_338),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_327),
.A2(n_264),
.B(n_261),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_303),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_364),
.A2(n_280),
.B1(n_175),
.B2(n_250),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_342),
.B(n_265),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_370),
.A2(n_192),
.B(n_175),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_364),
.A2(n_175),
.B1(n_239),
.B2(n_254),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_295),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_331),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_346),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_347),
.A2(n_287),
.B(n_239),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_331),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_341),
.B(n_286),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_354),
.B(n_65),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_361),
.B(n_287),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_336),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_310),
.B(n_175),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_336),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_367),
.B(n_320),
.Y(n_448)
);

INVx8_ASAP7_75t_L g449 ( 
.A(n_307),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_370),
.A2(n_192),
.B(n_175),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_345),
.Y(n_451)
);

BUFx4f_ASAP7_75t_L g452 ( 
.A(n_310),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_354),
.B(n_145),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_345),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_324),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_339),
.Y(n_456)
);

BUFx12f_ASAP7_75t_L g457 ( 
.A(n_324),
.Y(n_457)
);

OAI21xp33_ASAP7_75t_SL g458 ( 
.A1(n_290),
.A2(n_192),
.B(n_191),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_371),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_356),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_348),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_343),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_348),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_349),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_349),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_373),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_292),
.A2(n_192),
.B(n_132),
.Y(n_467)
);

NAND3xp33_ASAP7_75t_SL g468 ( 
.A(n_373),
.B(n_56),
.C(n_65),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_337),
.A2(n_191),
.B1(n_185),
.B2(n_145),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_337),
.B(n_303),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_337),
.B(n_191),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_365),
.B(n_371),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_365),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_329),
.B(n_65),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_324),
.Y(n_475)
);

NOR2x1_ASAP7_75t_L g476 ( 
.A(n_290),
.B(n_185),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_304),
.B(n_350),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_355),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_303),
.B(n_185),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_371),
.B(n_145),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_360),
.Y(n_481)
);

AO31x2_ASAP7_75t_L g482 ( 
.A1(n_377),
.A2(n_330),
.A3(n_352),
.B(n_369),
.Y(n_482)
);

OAI21x1_ASAP7_75t_L g483 ( 
.A1(n_394),
.A2(n_344),
.B(n_292),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_390),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_399),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_416),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_403),
.A2(n_316),
.B(n_314),
.Y(n_487)
);

AOI21x1_ASAP7_75t_SL g488 ( 
.A1(n_375),
.A2(n_372),
.B(n_356),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_435),
.A2(n_353),
.B(n_145),
.Y(n_489)
);

O2A1O1Ixp5_ASAP7_75t_L g490 ( 
.A1(n_412),
.A2(n_372),
.B(n_185),
.C(n_192),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_450),
.A2(n_155),
.B(n_147),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_378),
.B(n_414),
.Y(n_492)
);

OR2x6_ASAP7_75t_L g493 ( 
.A(n_449),
.B(n_446),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_356),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_389),
.A2(n_368),
.B(n_309),
.Y(n_495)
);

AOI21x1_ASAP7_75t_L g496 ( 
.A1(n_415),
.A2(n_368),
.B(n_154),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_414),
.A2(n_303),
.B1(n_368),
.B2(n_309),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_397),
.A2(n_154),
.B(n_151),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_421),
.B(n_368),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_428),
.A2(n_151),
.B(n_154),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_383),
.A2(n_419),
.B(n_411),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_381),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_411),
.A2(n_309),
.B(n_132),
.Y(n_503)
);

NOR2xp67_ASAP7_75t_L g504 ( 
.A(n_404),
.B(n_309),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_383),
.A2(n_135),
.B(n_133),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_477),
.B(n_169),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_409),
.A2(n_325),
.B(n_169),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_391),
.Y(n_508)
);

OA21x2_ASAP7_75t_L g509 ( 
.A1(n_440),
.A2(n_155),
.B(n_169),
.Y(n_509)
);

AOI21xp33_ASAP7_75t_L g510 ( 
.A1(n_378),
.A2(n_68),
.B(n_2),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_413),
.B(n_325),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_379),
.B(n_168),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_400),
.A2(n_135),
.B(n_128),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_405),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_467),
.A2(n_168),
.B(n_167),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_431),
.A2(n_325),
.B(n_168),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_408),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_387),
.A2(n_167),
.B(n_164),
.Y(n_518)
);

AOI221xp5_ASAP7_75t_SL g519 ( 
.A1(n_443),
.A2(n_68),
.B1(n_164),
.B2(n_155),
.C(n_151),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_385),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_400),
.A2(n_133),
.B(n_135),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_437),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_385),
.B(n_167),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_462),
.B(n_68),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_466),
.B(n_1),
.Y(n_525)
);

NOR2xp67_ASAP7_75t_SL g526 ( 
.A(n_457),
.B(n_125),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_413),
.B(n_325),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_478),
.B(n_325),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_393),
.A2(n_134),
.B1(n_133),
.B2(n_132),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_427),
.A2(n_164),
.B(n_134),
.Y(n_530)
);

CKINVDCx8_ASAP7_75t_R g531 ( 
.A(n_455),
.Y(n_531)
);

NAND2x1p5_ASAP7_75t_L g532 ( 
.A(n_392),
.B(n_134),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_417),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_402),
.A2(n_134),
.B(n_133),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_436),
.A2(n_132),
.B(n_128),
.Y(n_535)
);

AO31x2_ASAP7_75t_L g536 ( 
.A1(n_433),
.A2(n_128),
.A3(n_4),
.B(n_5),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_381),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_476),
.A2(n_125),
.B(n_4),
.Y(n_538)
);

AND2x6_ASAP7_75t_L g539 ( 
.A(n_382),
.B(n_125),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_384),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_438),
.Y(n_541)
);

OAI21x1_ASAP7_75t_L g542 ( 
.A1(n_388),
.A2(n_3),
.B(n_7),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_393),
.A2(n_3),
.B(n_8),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_401),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_423),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_481),
.B(n_8),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_468),
.A2(n_9),
.B(n_12),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_448),
.B(n_9),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_396),
.B(n_12),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_388),
.A2(n_14),
.B(n_15),
.Y(n_550)
);

AO32x2_ASAP7_75t_L g551 ( 
.A1(n_376),
.A2(n_14),
.A3(n_16),
.B1(n_18),
.B2(n_22),
.Y(n_551)
);

AO31x2_ASAP7_75t_L g552 ( 
.A1(n_425),
.A2(n_16),
.A3(n_22),
.B(n_23),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_418),
.A2(n_24),
.B(n_25),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_453),
.A2(n_469),
.B(n_444),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_458),
.A2(n_25),
.B(n_27),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_474),
.B(n_28),
.Y(n_556)
);

OAI21x1_ASAP7_75t_L g557 ( 
.A1(n_471),
.A2(n_29),
.B(n_479),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_429),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_396),
.B(n_382),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_446),
.B(n_426),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_391),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_418),
.A2(n_410),
.B(n_424),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_430),
.B(n_439),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_459),
.B(n_472),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_461),
.Y(n_565)
);

AO32x2_ASAP7_75t_L g566 ( 
.A1(n_376),
.A2(n_422),
.A3(n_407),
.B1(n_398),
.B2(n_468),
.Y(n_566)
);

AOI21x1_ASAP7_75t_L g567 ( 
.A1(n_470),
.A2(n_471),
.B(n_434),
.Y(n_567)
);

AO31x2_ASAP7_75t_L g568 ( 
.A1(n_376),
.A2(n_464),
.A3(n_463),
.B(n_473),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_421),
.B(n_442),
.Y(n_569)
);

OAI21x1_ASAP7_75t_L g570 ( 
.A1(n_479),
.A2(n_470),
.B(n_445),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_441),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_447),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_452),
.A2(n_480),
.B(n_449),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_452),
.A2(n_449),
.B(n_459),
.Y(n_574)
);

A2O1A1Ixp33_ASAP7_75t_L g575 ( 
.A1(n_386),
.A2(n_406),
.B(n_395),
.C(n_454),
.Y(n_575)
);

OA21x2_ASAP7_75t_L g576 ( 
.A1(n_451),
.A2(n_465),
.B(n_376),
.Y(n_576)
);

NOR2xp67_ASAP7_75t_L g577 ( 
.A(n_460),
.B(n_398),
.Y(n_577)
);

AO22x1_ASAP7_75t_L g578 ( 
.A1(n_456),
.A2(n_460),
.B1(n_475),
.B2(n_420),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_420),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_401),
.B(n_391),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_422),
.A2(n_380),
.B(n_432),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_422),
.A2(n_391),
.B(n_432),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g583 ( 
.A1(n_380),
.A2(n_344),
.B(n_394),
.Y(n_583)
);

OAI21x1_ASAP7_75t_L g584 ( 
.A1(n_380),
.A2(n_344),
.B(n_394),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_432),
.B(n_380),
.Y(n_585)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_380),
.A2(n_344),
.B(n_394),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_432),
.B(n_380),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_405),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_384),
.Y(n_589)
);

BUFx8_ASAP7_75t_L g590 ( 
.A(n_455),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_378),
.B(n_414),
.Y(n_591)
);

OAI21x1_ASAP7_75t_L g592 ( 
.A1(n_394),
.A2(n_344),
.B(n_403),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_390),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_377),
.A2(n_257),
.B(n_226),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_378),
.B(n_414),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_499),
.B(n_493),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_494),
.A2(n_569),
.B1(n_556),
.B2(n_595),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_544),
.Y(n_598)
);

OA21x2_ASAP7_75t_L g599 ( 
.A1(n_519),
.A2(n_542),
.B(n_501),
.Y(n_599)
);

A2O1A1Ixp33_ASAP7_75t_L g600 ( 
.A1(n_492),
.A2(n_595),
.B(n_591),
.C(n_550),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_563),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_563),
.Y(n_602)
);

AO21x2_ASAP7_75t_L g603 ( 
.A1(n_581),
.A2(n_555),
.B(n_582),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_514),
.B(n_588),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_539),
.Y(n_605)
);

NAND2x1p5_ASAP7_75t_L g606 ( 
.A(n_495),
.B(n_489),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_520),
.Y(n_607)
);

OAI21x1_ASAP7_75t_L g608 ( 
.A1(n_583),
.A2(n_584),
.B(n_586),
.Y(n_608)
);

NOR2xp67_ASAP7_75t_L g609 ( 
.A(n_540),
.B(n_589),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_539),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_524),
.Y(n_611)
);

A2O1A1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_492),
.A2(n_591),
.B(n_555),
.C(n_562),
.Y(n_612)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_483),
.A2(n_592),
.B(n_534),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_539),
.Y(n_614)
);

OAI21x1_ASAP7_75t_L g615 ( 
.A1(n_495),
.A2(n_521),
.B(n_513),
.Y(n_615)
);

AOI21x1_ASAP7_75t_L g616 ( 
.A1(n_496),
.A2(n_521),
.B(n_503),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_517),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_499),
.B(n_493),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_560),
.A2(n_559),
.B1(n_497),
.B2(n_493),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_560),
.B(n_548),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_568),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_548),
.B(n_506),
.Y(n_622)
);

NAND2xp33_ASAP7_75t_L g623 ( 
.A(n_539),
.B(n_497),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_503),
.A2(n_487),
.B(n_491),
.Y(n_624)
);

OAI21x1_ASAP7_75t_L g625 ( 
.A1(n_530),
.A2(n_500),
.B(n_490),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_508),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_484),
.Y(n_627)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_535),
.A2(n_498),
.B(n_518),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_574),
.B(n_573),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_485),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g631 ( 
.A1(n_516),
.A2(n_570),
.B(n_515),
.Y(n_631)
);

AOI21x1_ASAP7_75t_L g632 ( 
.A1(n_594),
.A2(n_562),
.B(n_567),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_486),
.Y(n_633)
);

NAND2x1p5_ASAP7_75t_L g634 ( 
.A(n_557),
.B(n_554),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_523),
.Y(n_635)
);

CKINVDCx16_ASAP7_75t_R g636 ( 
.A(n_502),
.Y(n_636)
);

HB1xp67_ASAP7_75t_SL g637 ( 
.A(n_590),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_559),
.A2(n_527),
.B1(n_511),
.B2(n_531),
.Y(n_638)
);

O2A1O1Ixp33_ASAP7_75t_L g639 ( 
.A1(n_547),
.A2(n_510),
.B(n_553),
.C(n_546),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_564),
.B(n_546),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_568),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g642 ( 
.A1(n_516),
.A2(n_488),
.B(n_538),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_533),
.Y(n_643)
);

AND2x4_ASAP7_75t_SL g644 ( 
.A(n_580),
.B(n_561),
.Y(n_644)
);

BUFx2_ASAP7_75t_R g645 ( 
.A(n_537),
.Y(n_645)
);

OAI21x1_ASAP7_75t_L g646 ( 
.A1(n_581),
.A2(n_507),
.B(n_505),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_564),
.B(n_482),
.Y(n_647)
);

AO21x2_ASAP7_75t_L g648 ( 
.A1(n_594),
.A2(n_507),
.B(n_527),
.Y(n_648)
);

OA21x2_ASAP7_75t_L g649 ( 
.A1(n_543),
.A2(n_510),
.B(n_553),
.Y(n_649)
);

OAI21x1_ASAP7_75t_L g650 ( 
.A1(n_505),
.A2(n_509),
.B(n_587),
.Y(n_650)
);

OAI21x1_ASAP7_75t_L g651 ( 
.A1(n_509),
.A2(n_587),
.B(n_585),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_539),
.Y(n_652)
);

OA21x2_ASAP7_75t_L g653 ( 
.A1(n_543),
.A2(n_511),
.B(n_512),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_549),
.A2(n_590),
.B1(n_525),
.B2(n_593),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_568),
.Y(n_655)
);

AOI221xp5_ASAP7_75t_L g656 ( 
.A1(n_549),
.A2(n_545),
.B1(n_558),
.B2(n_578),
.C(n_565),
.Y(n_656)
);

AO21x2_ASAP7_75t_L g657 ( 
.A1(n_575),
.A2(n_528),
.B(n_585),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g658 ( 
.A1(n_529),
.A2(n_576),
.B(n_528),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_571),
.B(n_572),
.Y(n_659)
);

AOI222xp33_ASAP7_75t_L g660 ( 
.A1(n_577),
.A2(n_541),
.B1(n_522),
.B2(n_504),
.C1(n_526),
.C2(n_529),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_579),
.A2(n_561),
.B1(n_508),
.B2(n_576),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_508),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_566),
.B(n_552),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_566),
.Y(n_664)
);

NAND2x1p5_ASAP7_75t_L g665 ( 
.A(n_482),
.B(n_552),
.Y(n_665)
);

O2A1O1Ixp33_ASAP7_75t_SL g666 ( 
.A1(n_551),
.A2(n_566),
.B(n_552),
.C(n_536),
.Y(n_666)
);

NAND3xp33_ASAP7_75t_L g667 ( 
.A(n_536),
.B(n_551),
.C(n_482),
.Y(n_667)
);

OAI21x1_ASAP7_75t_L g668 ( 
.A1(n_532),
.A2(n_536),
.B(n_551),
.Y(n_668)
);

OAI21x1_ASAP7_75t_L g669 ( 
.A1(n_532),
.A2(n_584),
.B(n_583),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_510),
.A2(n_312),
.B1(n_319),
.B2(n_293),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_594),
.A2(n_377),
.B(n_318),
.Y(n_671)
);

OAI21x1_ASAP7_75t_L g672 ( 
.A1(n_583),
.A2(n_586),
.B(n_584),
.Y(n_672)
);

INVx6_ASAP7_75t_L g673 ( 
.A(n_493),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_517),
.Y(n_674)
);

OAI21x1_ASAP7_75t_L g675 ( 
.A1(n_583),
.A2(n_586),
.B(n_584),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_568),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_563),
.Y(n_677)
);

OAI21x1_ASAP7_75t_L g678 ( 
.A1(n_583),
.A2(n_586),
.B(n_584),
.Y(n_678)
);

OAI21x1_ASAP7_75t_L g679 ( 
.A1(n_583),
.A2(n_586),
.B(n_584),
.Y(n_679)
);

OA21x2_ASAP7_75t_L g680 ( 
.A1(n_519),
.A2(n_542),
.B(n_501),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_539),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_492),
.B(n_591),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_539),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_594),
.A2(n_377),
.B(n_318),
.Y(n_684)
);

O2A1O1Ixp33_ASAP7_75t_SL g685 ( 
.A1(n_492),
.A2(n_312),
.B(n_595),
.C(n_591),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_492),
.B(n_591),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_510),
.A2(n_312),
.B1(n_319),
.B2(n_293),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_517),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_517),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_580),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_517),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_594),
.A2(n_377),
.B(n_318),
.Y(n_692)
);

CKINVDCx11_ASAP7_75t_R g693 ( 
.A(n_531),
.Y(n_693)
);

OAI21x1_ASAP7_75t_L g694 ( 
.A1(n_583),
.A2(n_586),
.B(n_584),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_517),
.Y(n_695)
);

BUFx2_ASAP7_75t_R g696 ( 
.A(n_589),
.Y(n_696)
);

OAI21x1_ASAP7_75t_SL g697 ( 
.A1(n_495),
.A2(n_581),
.B(n_562),
.Y(n_697)
);

AO21x2_ASAP7_75t_L g698 ( 
.A1(n_501),
.A2(n_377),
.B(n_581),
.Y(n_698)
);

AOI21x1_ASAP7_75t_SL g699 ( 
.A1(n_629),
.A2(n_663),
.B(n_640),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_598),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_620),
.B(n_622),
.Y(n_701)
);

NOR2xp67_ASAP7_75t_L g702 ( 
.A(n_690),
.B(n_604),
.Y(n_702)
);

CKINVDCx12_ASAP7_75t_R g703 ( 
.A(n_696),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_670),
.A2(n_687),
.B1(n_597),
.B2(n_654),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_682),
.A2(n_611),
.B1(n_686),
.B2(n_690),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_647),
.B(n_698),
.Y(n_706)
);

CKINVDCx6p67_ASAP7_75t_R g707 ( 
.A(n_693),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_663),
.B(n_647),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_653),
.B(n_648),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_607),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_686),
.A2(n_612),
.B1(n_600),
.B2(n_656),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_627),
.Y(n_712)
);

O2A1O1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_639),
.A2(n_685),
.B(n_638),
.C(n_692),
.Y(n_713)
);

NOR2xp67_ASAP7_75t_L g714 ( 
.A(n_609),
.B(n_617),
.Y(n_714)
);

OA21x2_ASAP7_75t_L g715 ( 
.A1(n_615),
.A2(n_625),
.B(n_675),
.Y(n_715)
);

OA21x2_ASAP7_75t_L g716 ( 
.A1(n_615),
.A2(n_625),
.B(n_675),
.Y(n_716)
);

AOI21x1_ASAP7_75t_SL g717 ( 
.A1(n_629),
.A2(n_659),
.B(n_596),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_629),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_653),
.B(n_648),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_630),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_601),
.B(n_602),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_698),
.B(n_665),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_651),
.Y(n_723)
);

O2A1O1Ixp5_ASAP7_75t_L g724 ( 
.A1(n_671),
.A2(n_684),
.B(n_632),
.C(n_667),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_596),
.B(n_618),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_653),
.B(n_648),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_623),
.A2(n_698),
.B(n_603),
.Y(n_727)
);

O2A1O1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_623),
.A2(n_619),
.B(n_635),
.C(n_649),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_607),
.Y(n_729)
);

NOR2xp67_ASAP7_75t_L g730 ( 
.A(n_617),
.B(n_674),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_L g731 ( 
.A(n_674),
.B(n_688),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_653),
.B(n_677),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_662),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_665),
.B(n_621),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_693),
.Y(n_735)
);

BUFx4f_ASAP7_75t_L g736 ( 
.A(n_673),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_596),
.B(n_618),
.Y(n_737)
);

AND2x4_ASAP7_75t_L g738 ( 
.A(n_618),
.B(n_633),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_659),
.B(n_688),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_662),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_626),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_643),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_651),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_621),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_626),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_689),
.B(n_695),
.Y(n_746)
);

O2A1O1Ixp5_ASAP7_75t_L g747 ( 
.A1(n_632),
.A2(n_616),
.B(n_681),
.C(n_614),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_641),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_673),
.A2(n_637),
.B1(n_598),
.B2(n_645),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_641),
.Y(n_750)
);

OA21x2_ASAP7_75t_L g751 ( 
.A1(n_608),
.A2(n_678),
.B(n_694),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_644),
.B(n_691),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_673),
.A2(n_644),
.B1(n_636),
.B2(n_661),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_668),
.B(n_665),
.Y(n_754)
);

OA21x2_ASAP7_75t_L g755 ( 
.A1(n_608),
.A2(n_679),
.B(n_694),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_673),
.A2(n_683),
.B1(n_652),
.B2(n_605),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_689),
.B(n_691),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_695),
.B(n_626),
.Y(n_758)
);

BUFx12f_ASAP7_75t_L g759 ( 
.A(n_626),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_655),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_649),
.B(n_660),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_655),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_649),
.B(n_657),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_676),
.Y(n_764)
);

NOR2xp67_ASAP7_75t_L g765 ( 
.A(n_626),
.B(n_652),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_657),
.B(n_681),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_649),
.B(n_657),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_676),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_668),
.B(n_664),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_605),
.A2(n_614),
.B1(n_683),
.B2(n_610),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_605),
.A2(n_614),
.B1(n_683),
.B2(n_610),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_646),
.A2(n_652),
.B(n_681),
.C(n_610),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_664),
.B(n_666),
.Y(n_773)
);

OA22x2_ASAP7_75t_L g774 ( 
.A1(n_697),
.A2(n_646),
.B1(n_642),
.B2(n_658),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_SL g775 ( 
.A1(n_603),
.A2(n_599),
.B(n_680),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_658),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_650),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_634),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_606),
.B(n_697),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_606),
.A2(n_634),
.B1(n_599),
.B2(n_680),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_642),
.B(n_669),
.Y(n_781)
);

NOR2x1_ASAP7_75t_SL g782 ( 
.A(n_616),
.B(n_606),
.Y(n_782)
);

AOI21x1_ASAP7_75t_SL g783 ( 
.A1(n_634),
.A2(n_599),
.B(n_680),
.Y(n_783)
);

CKINVDCx16_ASAP7_75t_R g784 ( 
.A(n_650),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_672),
.Y(n_785)
);

OA21x2_ASAP7_75t_L g786 ( 
.A1(n_672),
.A2(n_679),
.B(n_678),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_631),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_631),
.B(n_624),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_624),
.B(n_669),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_613),
.B(n_628),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_744),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_744),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_781),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_706),
.B(n_613),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_750),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_750),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_708),
.B(n_769),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_718),
.B(n_781),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_708),
.B(n_769),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_762),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_732),
.B(n_709),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_762),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_732),
.B(n_709),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_764),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_718),
.B(n_781),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_764),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_701),
.B(n_711),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_718),
.B(n_766),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_706),
.B(n_763),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_723),
.Y(n_810)
);

AO21x2_ASAP7_75t_L g811 ( 
.A1(n_775),
.A2(n_727),
.B(n_767),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_723),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_748),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_760),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_768),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_734),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_743),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_719),
.B(n_726),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_710),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_719),
.B(n_726),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_734),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_754),
.B(n_776),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_785),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_777),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_766),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_754),
.B(n_766),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_751),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_722),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_751),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_778),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_784),
.B(n_774),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_722),
.B(n_761),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_774),
.B(n_787),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_712),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_720),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_788),
.B(n_789),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_778),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_751),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_779),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_788),
.B(n_789),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_742),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_755),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_755),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_772),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_790),
.B(n_772),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_773),
.B(n_780),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_790),
.B(n_782),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_755),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_786),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_786),
.B(n_716),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_721),
.B(n_739),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_786),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_710),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_715),
.B(n_716),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_715),
.B(n_716),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_757),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_715),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_746),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_757),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_738),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_705),
.B(n_729),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_757),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_728),
.B(n_713),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_747),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_736),
.Y(n_865)
);

INVx5_ASAP7_75t_L g866 ( 
.A(n_758),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_724),
.B(n_738),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_813),
.Y(n_868)
);

AOI221xp5_ASAP7_75t_L g869 ( 
.A1(n_807),
.A2(n_704),
.B1(n_749),
.B2(n_753),
.C(n_738),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_818),
.B(n_758),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_818),
.B(n_758),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_818),
.B(n_820),
.Y(n_872)
);

INVx5_ASAP7_75t_SL g873 ( 
.A(n_865),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_813),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_837),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_822),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_813),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_818),
.B(n_737),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_809),
.B(n_741),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_820),
.B(n_725),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_820),
.B(n_725),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_828),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_832),
.B(n_731),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_828),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_807),
.A2(n_737),
.B1(n_725),
.B2(n_707),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_828),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_820),
.B(n_737),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_814),
.Y(n_888)
);

BUFx8_ASAP7_75t_L g889 ( 
.A(n_865),
.Y(n_889)
);

CKINVDCx11_ASAP7_75t_R g890 ( 
.A(n_819),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_803),
.B(n_730),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_814),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_810),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_810),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_803),
.B(n_801),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_814),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_803),
.B(n_752),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_803),
.B(n_752),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_812),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_837),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_793),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_801),
.B(n_752),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_793),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_815),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_801),
.B(n_756),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_815),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_815),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_791),
.Y(n_908)
);

INVxp67_ASAP7_75t_SL g909 ( 
.A(n_812),
.Y(n_909)
);

NOR2x1_ASAP7_75t_L g910 ( 
.A(n_863),
.B(n_714),
.Y(n_910)
);

OR2x6_ASAP7_75t_L g911 ( 
.A(n_867),
.B(n_771),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_836),
.B(n_770),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_824),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_836),
.B(n_745),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_822),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_791),
.Y(n_916)
);

AO31x2_ASAP7_75t_L g917 ( 
.A1(n_864),
.A2(n_783),
.A3(n_699),
.B(n_717),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_863),
.A2(n_707),
.B1(n_736),
.B2(n_702),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_809),
.B(n_745),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_836),
.B(n_745),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_809),
.B(n_745),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_836),
.B(n_840),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_865),
.A2(n_703),
.B1(n_700),
.B2(n_736),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_791),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_824),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_795),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_795),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_R g928 ( 
.A(n_865),
.B(n_703),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_795),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_SL g930 ( 
.A1(n_865),
.A2(n_735),
.B(n_733),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_796),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_824),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_840),
.B(n_765),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_840),
.B(n_733),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_840),
.B(n_740),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_832),
.B(n_740),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_822),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_796),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_837),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_846),
.A2(n_844),
.B(n_864),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_839),
.A2(n_700),
.B1(n_735),
.B2(n_759),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_822),
.B(n_759),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_824),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_832),
.B(n_821),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_816),
.B(n_821),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_792),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_845),
.B(n_799),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_845),
.B(n_799),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_792),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_845),
.B(n_799),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_823),
.Y(n_951)
);

NAND5xp2_ASAP7_75t_SL g952 ( 
.A(n_941),
.B(n_831),
.C(n_867),
.D(n_845),
.E(n_833),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_945),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_890),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_945),
.Y(n_955)
);

AO21x2_ASAP7_75t_L g956 ( 
.A1(n_940),
.A2(n_864),
.B(n_849),
.Y(n_956)
);

AOI222xp33_ASAP7_75t_L g957 ( 
.A1(n_869),
.A2(n_844),
.B1(n_831),
.B2(n_867),
.C1(n_839),
.C2(n_851),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_869),
.A2(n_861),
.B1(n_846),
.B2(n_865),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_868),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_910),
.A2(n_844),
.B(n_867),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_923),
.A2(n_865),
.B1(n_860),
.B2(n_808),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_878),
.B(n_799),
.Y(n_962)
);

NAND3xp33_ASAP7_75t_L g963 ( 
.A(n_940),
.B(n_846),
.C(n_861),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_910),
.B(n_860),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_913),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_SL g966 ( 
.A1(n_928),
.A2(n_831),
.B1(n_865),
.B2(n_860),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_913),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_923),
.A2(n_865),
.B1(n_860),
.B2(n_808),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_878),
.B(n_797),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_868),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_885),
.A2(n_861),
.B1(n_831),
.B2(n_858),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_918),
.A2(n_808),
.B1(n_805),
.B2(n_798),
.Y(n_972)
);

AO21x2_ASAP7_75t_L g973 ( 
.A1(n_909),
.A2(n_849),
.B(n_848),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_878),
.B(n_797),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_875),
.Y(n_975)
);

AOI221xp5_ASAP7_75t_L g976 ( 
.A1(n_883),
.A2(n_851),
.B1(n_816),
.B2(n_821),
.C(n_858),
.Y(n_976)
);

AOI211xp5_ASAP7_75t_L g977 ( 
.A1(n_930),
.A2(n_819),
.B(n_853),
.C(n_847),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_874),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_883),
.B(n_797),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_880),
.B(n_826),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_947),
.A2(n_833),
.B(n_853),
.C(n_825),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_880),
.B(n_797),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_874),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_875),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_936),
.A2(n_847),
.B(n_858),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_877),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_936),
.A2(n_862),
.B1(n_811),
.B2(n_835),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_889),
.A2(n_862),
.B1(n_811),
.B2(n_835),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_880),
.B(n_826),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_944),
.B(n_862),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_881),
.B(n_826),
.Y(n_991)
);

INVx5_ASAP7_75t_L g992 ( 
.A(n_901),
.Y(n_992)
);

NAND3xp33_ASAP7_75t_L g993 ( 
.A(n_911),
.B(n_794),
.C(n_944),
.Y(n_993)
);

OA21x2_ASAP7_75t_L g994 ( 
.A1(n_909),
.A2(n_849),
.B(n_843),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_911),
.A2(n_811),
.B(n_794),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_877),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_888),
.Y(n_997)
);

NAND3xp33_ASAP7_75t_SL g998 ( 
.A(n_944),
.B(n_847),
.C(n_879),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_888),
.Y(n_999)
);

NAND2xp33_ASAP7_75t_SL g1000 ( 
.A(n_942),
.B(n_841),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_892),
.Y(n_1001)
);

OAI211xp5_ASAP7_75t_L g1002 ( 
.A1(n_879),
.A2(n_833),
.B(n_816),
.C(n_856),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_889),
.A2(n_862),
.B1(n_811),
.B2(n_834),
.Y(n_1003)
);

NAND2xp33_ASAP7_75t_R g1004 ( 
.A(n_911),
.B(n_847),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_893),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_889),
.A2(n_811),
.B1(n_834),
.B2(n_835),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_881),
.B(n_826),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_919),
.B(n_856),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_881),
.B(n_859),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_892),
.Y(n_1010)
);

OAI211xp5_ASAP7_75t_L g1011 ( 
.A1(n_919),
.A2(n_833),
.B(n_825),
.C(n_841),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_889),
.A2(n_811),
.B1(n_841),
.B2(n_834),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_896),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_945),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_893),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_911),
.A2(n_808),
.B1(n_805),
.B2(n_798),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_887),
.B(n_825),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_896),
.Y(n_1018)
);

AOI221x1_ASAP7_75t_L g1019 ( 
.A1(n_908),
.A2(n_806),
.B1(n_796),
.B2(n_800),
.C(n_859),
.Y(n_1019)
);

NAND4xp25_ASAP7_75t_L g1020 ( 
.A(n_919),
.B(n_794),
.C(n_837),
.D(n_806),
.Y(n_1020)
);

NOR5xp2_ASAP7_75t_SL g1021 ( 
.A(n_911),
.B(n_830),
.C(n_852),
.D(n_838),
.E(n_793),
.Y(n_1021)
);

NOR3xp33_ASAP7_75t_L g1022 ( 
.A(n_921),
.B(n_830),
.C(n_859),
.Y(n_1022)
);

OAI221xp5_ASAP7_75t_L g1023 ( 
.A1(n_911),
.A2(n_830),
.B1(n_859),
.B2(n_793),
.C(n_866),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_889),
.A2(n_905),
.B1(n_873),
.B2(n_947),
.Y(n_1024)
);

AOI33xp33_ASAP7_75t_L g1025 ( 
.A1(n_904),
.A2(n_806),
.A3(n_800),
.B1(n_854),
.B2(n_855),
.B3(n_792),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_905),
.A2(n_808),
.B1(n_859),
.B2(n_866),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_921),
.B(n_905),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_921),
.B(n_872),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_891),
.B(n_887),
.Y(n_1029)
);

OA21x2_ASAP7_75t_L g1030 ( 
.A1(n_893),
.A2(n_829),
.B(n_827),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_875),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_873),
.A2(n_866),
.B1(n_942),
.B2(n_939),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_904),
.Y(n_1033)
);

AOI221xp5_ASAP7_75t_L g1034 ( 
.A1(n_947),
.A2(n_859),
.B1(n_808),
.B2(n_800),
.C(n_798),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_900),
.Y(n_1035)
);

NAND3xp33_ASAP7_75t_L g1036 ( 
.A(n_882),
.B(n_830),
.C(n_866),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_887),
.B(n_866),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_894),
.Y(n_1038)
);

OAI221xp5_ASAP7_75t_SL g1039 ( 
.A1(n_876),
.A2(n_850),
.B1(n_792),
.B2(n_802),
.C(n_804),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_934),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_906),
.Y(n_1041)
);

OAI211xp5_ASAP7_75t_SL g1042 ( 
.A1(n_906),
.A2(n_817),
.B(n_857),
.C(n_852),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_907),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_900),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_870),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_873),
.A2(n_866),
.B1(n_805),
.B2(n_798),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_873),
.A2(n_805),
.B1(n_798),
.B2(n_866),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_870),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_870),
.B(n_866),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_959),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_954),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_1000),
.Y(n_1052)
);

OA21x2_ASAP7_75t_L g1053 ( 
.A1(n_995),
.A2(n_848),
.B(n_827),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_970),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_976),
.B(n_979),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_957),
.B(n_948),
.Y(n_1056)
);

OA21x2_ASAP7_75t_L g1057 ( 
.A1(n_1019),
.A2(n_848),
.B(n_827),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_978),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_983),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_975),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_986),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_996),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_960),
.A2(n_838),
.B(n_852),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_973),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_997),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_1027),
.Y(n_1066)
);

NOR2x1_ASAP7_75t_SL g1067 ( 
.A(n_964),
.B(n_901),
.Y(n_1067)
);

NOR2x1p5_ASAP7_75t_L g1068 ( 
.A(n_1020),
.B(n_900),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_963),
.B(n_948),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_973),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1037),
.B(n_948),
.Y(n_1071)
);

INVx5_ASAP7_75t_L g1072 ( 
.A(n_992),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_999),
.Y(n_1073)
);

NAND3xp33_ASAP7_75t_L g1074 ( 
.A(n_958),
.B(n_882),
.C(n_884),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_985),
.B(n_950),
.Y(n_1075)
);

OA21x2_ASAP7_75t_L g1076 ( 
.A1(n_1036),
.A2(n_987),
.B(n_993),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1001),
.Y(n_1077)
);

AND2x2_ASAP7_75t_SL g1078 ( 
.A(n_1025),
.B(n_901),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_994),
.Y(n_1079)
);

NAND2x1_ASAP7_75t_L g1080 ( 
.A(n_994),
.B(n_901),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_994),
.Y(n_1081)
);

INVx4_ASAP7_75t_SL g1082 ( 
.A(n_975),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_1008),
.B(n_984),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1030),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1030),
.Y(n_1085)
);

OR2x6_ASAP7_75t_L g1086 ( 
.A(n_964),
.B(n_901),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_962),
.B(n_950),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1010),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1013),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1018),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_1028),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_992),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_953),
.Y(n_1093)
);

AND2x6_ASAP7_75t_SL g1094 ( 
.A(n_1017),
.B(n_1029),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1030),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1049),
.B(n_950),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1005),
.Y(n_1097)
);

NOR2x1p5_ASAP7_75t_L g1098 ( 
.A(n_998),
.B(n_939),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1005),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_955),
.B(n_1014),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1033),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1015),
.Y(n_1102)
);

OA21x2_ASAP7_75t_L g1103 ( 
.A1(n_987),
.A2(n_843),
.B(n_848),
.Y(n_1103)
);

OA21x2_ASAP7_75t_L g1104 ( 
.A1(n_988),
.A2(n_827),
.B(n_843),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_992),
.B(n_922),
.Y(n_1105)
);

INVxp67_ASAP7_75t_R g1106 ( 
.A(n_1032),
.Y(n_1106)
);

INVx4_ASAP7_75t_SL g1107 ( 
.A(n_975),
.Y(n_1107)
);

BUFx8_ASAP7_75t_L g1108 ( 
.A(n_975),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1041),
.Y(n_1109)
);

INVx5_ASAP7_75t_L g1110 ( 
.A(n_992),
.Y(n_1110)
);

OA21x2_ASAP7_75t_L g1111 ( 
.A1(n_988),
.A2(n_829),
.B(n_843),
.Y(n_1111)
);

INVx5_ASAP7_75t_L g1112 ( 
.A(n_1035),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1015),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1043),
.Y(n_1114)
);

OA21x2_ASAP7_75t_L g1115 ( 
.A1(n_1003),
.A2(n_842),
.B(n_829),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_965),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_1035),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1038),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_969),
.B(n_871),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_1044),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_965),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_967),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_974),
.B(n_871),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_977),
.B(n_901),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_967),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_1038),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_1031),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_956),
.Y(n_1128)
);

INVx4_ASAP7_75t_SL g1129 ( 
.A(n_1031),
.Y(n_1129)
);

OR2x2_ASAP7_75t_L g1130 ( 
.A(n_990),
.B(n_872),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_956),
.Y(n_1131)
);

OAI21xp33_ASAP7_75t_SL g1132 ( 
.A1(n_1124),
.A2(n_1025),
.B(n_958),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1055),
.B(n_1017),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1079),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1059),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1059),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1079),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1061),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_1052),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1068),
.A2(n_952),
.B1(n_971),
.B2(n_1023),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_1069),
.B(n_1039),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1081),
.Y(n_1142)
);

OAI222xp33_ASAP7_75t_L g1143 ( 
.A1(n_1056),
.A2(n_968),
.B1(n_961),
.B2(n_971),
.C1(n_972),
.C2(n_966),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1106),
.B(n_980),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1106),
.B(n_980),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1105),
.B(n_922),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1061),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1072),
.B(n_1016),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_1080),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1062),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1105),
.B(n_922),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_1117),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1081),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1105),
.B(n_872),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1066),
.B(n_981),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1062),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1052),
.B(n_1098),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1065),
.Y(n_1158)
);

AND4x1_ASAP7_75t_L g1159 ( 
.A(n_1074),
.B(n_1006),
.C(n_1012),
.D(n_1003),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1071),
.B(n_895),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1071),
.B(n_895),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_1112),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_1116),
.B(n_981),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1127),
.B(n_982),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1084),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_1112),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1096),
.B(n_1129),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1127),
.B(n_871),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_1121),
.B(n_1122),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_1117),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1065),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1083),
.A2(n_1024),
.B1(n_1006),
.B2(n_1012),
.Y(n_1172)
);

NAND5xp2_ASAP7_75t_L g1173 ( 
.A(n_1075),
.B(n_1024),
.C(n_1047),
.D(n_1034),
.E(n_1026),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1073),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1096),
.B(n_895),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1073),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1084),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1072),
.B(n_1022),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1077),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1129),
.B(n_989),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1129),
.B(n_991),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1077),
.Y(n_1182)
);

INVxp67_ASAP7_75t_SL g1183 ( 
.A(n_1067),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1078),
.B(n_902),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1085),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_1072),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1088),
.Y(n_1187)
);

INVx5_ASAP7_75t_SL g1188 ( 
.A(n_1060),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_1072),
.B(n_901),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_1060),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1072),
.B(n_1022),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_1112),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1088),
.Y(n_1193)
);

NAND5xp2_ASAP7_75t_L g1194 ( 
.A(n_1094),
.B(n_1026),
.C(n_1002),
.D(n_1011),
.E(n_942),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1089),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1089),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1085),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1051),
.B(n_1007),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1120),
.B(n_1046),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1129),
.B(n_1009),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1122),
.B(n_876),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1112),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1095),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1078),
.B(n_1067),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1095),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_1141),
.B(n_1125),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1141),
.B(n_1125),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1152),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1187),
.Y(n_1209)
);

INVx2_ASAP7_75t_SL g1210 ( 
.A(n_1167),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1135),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1134),
.Y(n_1212)
);

NAND2x1p5_ASAP7_75t_L g1213 ( 
.A(n_1186),
.B(n_1110),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1167),
.B(n_1082),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1134),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1135),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1186),
.B(n_1082),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1157),
.B(n_1082),
.Y(n_1218)
);

NAND2x1p5_ASAP7_75t_L g1219 ( 
.A(n_1186),
.B(n_1110),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1157),
.B(n_1082),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1134),
.Y(n_1221)
);

INVxp67_ASAP7_75t_L g1222 ( 
.A(n_1170),
.Y(n_1222)
);

INVx2_ASAP7_75t_SL g1223 ( 
.A(n_1186),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1133),
.B(n_1051),
.Y(n_1224)
);

AOI21xp33_ASAP7_75t_SL g1225 ( 
.A1(n_1199),
.A2(n_1076),
.B(n_1086),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1169),
.B(n_1076),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1136),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1198),
.B(n_1120),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1137),
.Y(n_1229)
);

INVx1_ASAP7_75t_SL g1230 ( 
.A(n_1139),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1169),
.B(n_1076),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1139),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1136),
.Y(n_1233)
);

NOR2x1_ASAP7_75t_L g1234 ( 
.A(n_1190),
.B(n_1120),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1138),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1190),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1201),
.B(n_1076),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1132),
.B(n_1091),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1132),
.B(n_1050),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1138),
.Y(n_1240)
);

NOR2x1_ASAP7_75t_L g1241 ( 
.A(n_1194),
.B(n_1092),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1140),
.B(n_1054),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1137),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1147),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1147),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1200),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1137),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1150),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1159),
.B(n_1058),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1162),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1144),
.B(n_1107),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1150),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1144),
.B(n_1107),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1156),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1145),
.B(n_1107),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1145),
.B(n_1107),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1156),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1158),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1159),
.B(n_1090),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1142),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1204),
.B(n_1086),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1158),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1230),
.B(n_1171),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1214),
.B(n_1218),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1232),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1211),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1222),
.B(n_1160),
.Y(n_1267)
);

NAND2xp33_ASAP7_75t_SL g1268 ( 
.A(n_1249),
.B(n_1204),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1214),
.B(n_1188),
.Y(n_1269)
);

INVx4_ASAP7_75t_L g1270 ( 
.A(n_1217),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1211),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_1218),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1220),
.Y(n_1273)
);

AND2x4_ASAP7_75t_L g1274 ( 
.A(n_1234),
.B(n_1251),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1213),
.A2(n_1189),
.B(n_1149),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1208),
.B(n_1160),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1241),
.B(n_1161),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1227),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1224),
.B(n_1161),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1246),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1220),
.B(n_1188),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_1253),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1251),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1253),
.B(n_1256),
.Y(n_1284)
);

NOR2x1_ASAP7_75t_L g1285 ( 
.A(n_1217),
.B(n_1251),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1246),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1228),
.B(n_1143),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1256),
.B(n_1188),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1255),
.B(n_1188),
.Y(n_1289)
);

NAND2xp33_ASAP7_75t_R g1290 ( 
.A(n_1217),
.B(n_1092),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1210),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1242),
.B(n_1173),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1206),
.B(n_1207),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1227),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1210),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_1255),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_1255),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1250),
.Y(n_1298)
);

NOR2x1_ASAP7_75t_L g1299 ( 
.A(n_1226),
.B(n_1231),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1248),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1259),
.A2(n_1173),
.B1(n_1148),
.B2(n_1172),
.Y(n_1301)
);

NOR2x1_ASAP7_75t_L g1302 ( 
.A(n_1226),
.B(n_1231),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1248),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1209),
.B(n_1175),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1261),
.B(n_1188),
.Y(n_1305)
);

INVx1_ASAP7_75t_SL g1306 ( 
.A(n_1206),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1213),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1239),
.B(n_1236),
.Y(n_1308)
);

INVx1_ASAP7_75t_SL g1309 ( 
.A(n_1207),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1252),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1238),
.A2(n_1148),
.B1(n_1180),
.B2(n_1181),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1225),
.A2(n_1155),
.B1(n_1184),
.B2(n_1183),
.Y(n_1312)
);

INVx3_ASAP7_75t_SL g1313 ( 
.A(n_1223),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1223),
.B(n_1162),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1261),
.A2(n_1148),
.B1(n_1180),
.B2(n_1181),
.Y(n_1315)
);

AOI322xp5_ASAP7_75t_L g1316 ( 
.A1(n_1292),
.A2(n_1128),
.A3(n_1148),
.B1(n_1258),
.B2(n_1257),
.C1(n_1233),
.C2(n_1235),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1264),
.B(n_1200),
.Y(n_1317)
);

OAI221xp5_ASAP7_75t_L g1318 ( 
.A1(n_1301),
.A2(n_1213),
.B1(n_1219),
.B2(n_1237),
.C(n_1155),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1272),
.B(n_1216),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1287),
.A2(n_1237),
.B(n_1219),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1306),
.B(n_1240),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1264),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1273),
.B(n_1282),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1268),
.A2(n_1178),
.B1(n_1191),
.B2(n_1219),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1270),
.B(n_1164),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1298),
.B(n_1309),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1312),
.A2(n_1191),
.B1(n_1178),
.B2(n_1192),
.Y(n_1327)
);

AND2x2_ASAP7_75t_SL g1328 ( 
.A(n_1274),
.B(n_1178),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1293),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1284),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1308),
.A2(n_1163),
.B1(n_1086),
.B2(n_1110),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1268),
.A2(n_1192),
.B(n_1166),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1293),
.Y(n_1333)
);

XOR2x2_ASAP7_75t_L g1334 ( 
.A(n_1285),
.B(n_1189),
.Y(n_1334)
);

AOI311xp33_ASAP7_75t_L g1335 ( 
.A1(n_1265),
.A2(n_1262),
.A3(n_1254),
.B(n_1252),
.C(n_1244),
.Y(n_1335)
);

INVxp67_ASAP7_75t_L g1336 ( 
.A(n_1284),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1299),
.A2(n_1202),
.B(n_1166),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1302),
.Y(n_1338)
);

OAI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1277),
.A2(n_1163),
.B1(n_1004),
.B2(n_1086),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1311),
.A2(n_1110),
.B1(n_1112),
.B2(n_1149),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1266),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1270),
.B(n_1202),
.Y(n_1342)
);

O2A1O1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1296),
.A2(n_1245),
.B(n_1254),
.C(n_1262),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1276),
.B(n_1201),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1269),
.B(n_1146),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1266),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1271),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1269),
.B(n_1146),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1283),
.Y(n_1349)
);

OAI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1290),
.A2(n_1004),
.B1(n_1110),
.B2(n_1189),
.Y(n_1350)
);

OAI21xp33_ASAP7_75t_L g1351 ( 
.A1(n_1279),
.A2(n_1191),
.B(n_1178),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1283),
.Y(n_1352)
);

O2A1O1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1297),
.A2(n_1191),
.B(n_1247),
.C(n_1243),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1315),
.A2(n_1149),
.B1(n_1115),
.B2(n_1111),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1274),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1280),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1288),
.A2(n_1281),
.B(n_1274),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1305),
.A2(n_1154),
.B1(n_1151),
.B2(n_1108),
.Y(n_1358)
);

NAND3xp33_ASAP7_75t_L g1359 ( 
.A(n_1270),
.B(n_1260),
.C(n_1247),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1313),
.A2(n_1263),
.B1(n_1291),
.B2(n_1295),
.Y(n_1360)
);

O2A1O1Ixp5_ASAP7_75t_SL g1361 ( 
.A1(n_1271),
.A2(n_1149),
.B(n_1179),
.C(n_1171),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1313),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1291),
.B(n_1175),
.Y(n_1363)
);

AOI32xp33_ASAP7_75t_L g1364 ( 
.A1(n_1281),
.A2(n_1131),
.A3(n_1154),
.B1(n_1151),
.B2(n_1092),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1305),
.A2(n_1103),
.B1(n_1115),
.B2(n_1111),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1330),
.B(n_1295),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1356),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1318),
.A2(n_1288),
.B1(n_1267),
.B2(n_1304),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1352),
.B(n_1263),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1328),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1349),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1362),
.B(n_1280),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1336),
.B(n_1286),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1355),
.B(n_1286),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1322),
.B(n_1314),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1329),
.B(n_1314),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1338),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1324),
.A2(n_1307),
.B1(n_1289),
.B2(n_1314),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1326),
.B(n_1303),
.Y(n_1379)
);

NAND2x1_ASAP7_75t_L g1380 ( 
.A(n_1317),
.B(n_1289),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1333),
.B(n_1307),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1360),
.B(n_1278),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1360),
.B(n_1278),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1327),
.A2(n_1358),
.B1(n_1320),
.B2(n_1323),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1341),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1346),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1345),
.B(n_1275),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1337),
.B(n_1275),
.Y(n_1388)
);

OAI221xp5_ASAP7_75t_L g1389 ( 
.A1(n_1357),
.A2(n_1310),
.B1(n_1300),
.B2(n_1294),
.C(n_1260),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1337),
.Y(n_1390)
);

INVxp67_ASAP7_75t_SL g1391 ( 
.A(n_1353),
.Y(n_1391)
);

NAND2xp33_ASAP7_75t_SL g1392 ( 
.A(n_1321),
.B(n_1294),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1348),
.B(n_1300),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1342),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1316),
.B(n_1310),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1347),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1325),
.B(n_1212),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1334),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1319),
.B(n_1174),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1321),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1343),
.B(n_1174),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_1344),
.Y(n_1402)
);

O2A1O1Ixp5_ASAP7_75t_SL g1403 ( 
.A1(n_1395),
.A2(n_1340),
.B(n_1331),
.C(n_1335),
.Y(n_1403)
);

OA22x2_ASAP7_75t_L g1404 ( 
.A1(n_1395),
.A2(n_1351),
.B1(n_1340),
.B2(n_1354),
.Y(n_1404)
);

NOR2xp67_ASAP7_75t_L g1405 ( 
.A(n_1369),
.B(n_1359),
.Y(n_1405)
);

OAI32xp33_ASAP7_75t_L g1406 ( 
.A1(n_1390),
.A2(n_1331),
.A3(n_1354),
.B1(n_1363),
.B2(n_1361),
.Y(n_1406)
);

AOI221xp5_ASAP7_75t_L g1407 ( 
.A1(n_1391),
.A2(n_1339),
.B1(n_1332),
.B2(n_1350),
.C(n_1364),
.Y(n_1407)
);

OAI322xp33_ASAP7_75t_L g1408 ( 
.A1(n_1382),
.A2(n_1215),
.A3(n_1243),
.B1(n_1229),
.B2(n_1221),
.C1(n_1212),
.C2(n_1131),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_R g1409 ( 
.A(n_1392),
.B(n_1108),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1393),
.B(n_1176),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1368),
.A2(n_1365),
.B1(n_1060),
.B2(n_1168),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1369),
.B(n_1060),
.Y(n_1412)
);

AOI221xp5_ASAP7_75t_L g1413 ( 
.A1(n_1392),
.A2(n_1229),
.B1(n_1221),
.B2(n_1215),
.C(n_1142),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1388),
.A2(n_1383),
.B(n_1401),
.Y(n_1414)
);

AOI221xp5_ASAP7_75t_L g1415 ( 
.A1(n_1378),
.A2(n_1142),
.B1(n_1153),
.B2(n_1203),
.C(n_1197),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1381),
.Y(n_1416)
);

NAND3xp33_ASAP7_75t_SL g1417 ( 
.A(n_1402),
.B(n_1080),
.C(n_1203),
.Y(n_1417)
);

AOI221x1_ASAP7_75t_L g1418 ( 
.A1(n_1371),
.A2(n_1176),
.B1(n_1179),
.B2(n_1182),
.C(n_1196),
.Y(n_1418)
);

NOR3x1_ASAP7_75t_L g1419 ( 
.A(n_1380),
.B(n_1182),
.C(n_1196),
.Y(n_1419)
);

AOI321xp33_ASAP7_75t_L g1420 ( 
.A1(n_1384),
.A2(n_1205),
.A3(n_1203),
.B1(n_1197),
.B2(n_1165),
.C(n_1177),
.Y(n_1420)
);

AOI221xp5_ASAP7_75t_L g1421 ( 
.A1(n_1400),
.A2(n_1153),
.B1(n_1197),
.B2(n_1205),
.C(n_1165),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1388),
.A2(n_1063),
.B(n_1195),
.Y(n_1422)
);

NAND2x1_ASAP7_75t_L g1423 ( 
.A(n_1387),
.B(n_1193),
.Y(n_1423)
);

OAI222xp33_ASAP7_75t_L g1424 ( 
.A1(n_1370),
.A2(n_1064),
.B1(n_1070),
.B2(n_1153),
.C1(n_1185),
.C2(n_1177),
.Y(n_1424)
);

AOI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1389),
.A2(n_1205),
.B1(n_1165),
.B2(n_1177),
.C(n_1185),
.Y(n_1425)
);

INVxp67_ASAP7_75t_L g1426 ( 
.A(n_1376),
.Y(n_1426)
);

OAI211xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1394),
.A2(n_1185),
.B(n_1195),
.C(n_1193),
.Y(n_1427)
);

NOR3xp33_ASAP7_75t_L g1428 ( 
.A(n_1372),
.B(n_1070),
.C(n_1064),
.Y(n_1428)
);

NAND2x1_ASAP7_75t_L g1429 ( 
.A(n_1387),
.B(n_1060),
.Y(n_1429)
);

OAI221xp5_ASAP7_75t_L g1430 ( 
.A1(n_1370),
.A2(n_1104),
.B1(n_1111),
.B2(n_1115),
.C(n_1103),
.Y(n_1430)
);

OAI211xp5_ASAP7_75t_L g1431 ( 
.A1(n_1366),
.A2(n_1115),
.B(n_1111),
.C(n_1104),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1393),
.B(n_1101),
.Y(n_1432)
);

O2A1O1Ixp5_ASAP7_75t_L g1433 ( 
.A1(n_1398),
.A2(n_1114),
.B(n_1109),
.C(n_1101),
.Y(n_1433)
);

AOI211xp5_ASAP7_75t_L g1434 ( 
.A1(n_1398),
.A2(n_1063),
.B(n_1042),
.C(n_1109),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1375),
.A2(n_1104),
.B1(n_1103),
.B2(n_1093),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1416),
.B(n_1367),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1404),
.A2(n_1397),
.B1(n_1373),
.B2(n_1377),
.Y(n_1437)
);

OAI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1414),
.A2(n_1374),
.B1(n_1379),
.B2(n_1381),
.C(n_1399),
.Y(n_1438)
);

AOI211xp5_ASAP7_75t_L g1439 ( 
.A1(n_1406),
.A2(n_1379),
.B(n_1397),
.C(n_1377),
.Y(n_1439)
);

AOI221xp5_ASAP7_75t_L g1440 ( 
.A1(n_1407),
.A2(n_1411),
.B1(n_1408),
.B2(n_1426),
.C(n_1433),
.Y(n_1440)
);

AOI21xp33_ASAP7_75t_L g1441 ( 
.A1(n_1404),
.A2(n_1396),
.B(n_1386),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_1405),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1429),
.Y(n_1443)
);

AOI221xp5_ASAP7_75t_L g1444 ( 
.A1(n_1422),
.A2(n_1385),
.B1(n_1099),
.B2(n_1097),
.C(n_1118),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1423),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1410),
.Y(n_1446)
);

AOI322xp5_ASAP7_75t_L g1447 ( 
.A1(n_1403),
.A2(n_1040),
.A3(n_915),
.B1(n_937),
.B2(n_1087),
.C1(n_933),
.C2(n_891),
.Y(n_1447)
);

A2O1A1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1420),
.A2(n_1099),
.B(n_1102),
.C(n_1097),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1419),
.Y(n_1449)
);

NOR2x1_ASAP7_75t_L g1450 ( 
.A(n_1412),
.B(n_1126),
.Y(n_1450)
);

AOI221xp5_ASAP7_75t_L g1451 ( 
.A1(n_1417),
.A2(n_1102),
.B1(n_1113),
.B2(n_1118),
.C(n_1126),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1432),
.B(n_1126),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1409),
.B(n_1113),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1435),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1418),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1427),
.Y(n_1456)
);

OAI211xp5_ASAP7_75t_SL g1457 ( 
.A1(n_1413),
.A2(n_1123),
.B(n_1119),
.C(n_1130),
.Y(n_1457)
);

AOI22x1_ASAP7_75t_L g1458 ( 
.A1(n_1424),
.A2(n_1108),
.B1(n_1100),
.B2(n_1021),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1434),
.A2(n_1104),
.B1(n_1103),
.B2(n_1100),
.Y(n_1459)
);

NOR2x1_ASAP7_75t_L g1460 ( 
.A(n_1431),
.B(n_1057),
.Y(n_1460)
);

AOI211xp5_ASAP7_75t_SL g1461 ( 
.A1(n_1428),
.A2(n_1021),
.B(n_937),
.C(n_915),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1415),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1436),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1436),
.Y(n_1464)
);

NOR2x1_ASAP7_75t_L g1465 ( 
.A(n_1443),
.B(n_1430),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1442),
.B(n_1425),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1437),
.B(n_1130),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1449),
.B(n_1421),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1445),
.Y(n_1469)
);

OAI21xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1460),
.A2(n_903),
.B(n_933),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1443),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1455),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1438),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1456),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1439),
.B(n_935),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1446),
.Y(n_1476)
);

OAI21xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1447),
.A2(n_903),
.B(n_933),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1453),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1462),
.B(n_1048),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1473),
.A2(n_1440),
.B1(n_1454),
.B2(n_1441),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1463),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1464),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1467),
.A2(n_1450),
.B1(n_1452),
.B2(n_1458),
.Y(n_1483)
);

AOI211xp5_ASAP7_75t_L g1484 ( 
.A1(n_1466),
.A2(n_1459),
.B(n_1444),
.C(n_1457),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1471),
.B(n_1451),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1469),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1465),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1472),
.B(n_1448),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1479),
.A2(n_1053),
.B1(n_1461),
.B2(n_939),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1468),
.Y(n_1490)
);

XNOR2x1_ASAP7_75t_L g1491 ( 
.A(n_1474),
.B(n_1053),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1475),
.A2(n_1053),
.B(n_1057),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1478),
.B(n_1045),
.Y(n_1493)
);

XOR2xp5_ASAP7_75t_L g1494 ( 
.A(n_1476),
.B(n_1477),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1487),
.A2(n_1470),
.B(n_1477),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1481),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1482),
.Y(n_1497)
);

OAI31xp33_ASAP7_75t_L g1498 ( 
.A1(n_1494),
.A2(n_1490),
.A3(n_1483),
.B(n_1491),
.Y(n_1498)
);

OAI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1480),
.A2(n_1053),
.B(n_903),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1485),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1486),
.B(n_1493),
.Y(n_1501)
);

NAND3x1_ASAP7_75t_L g1502 ( 
.A(n_1488),
.B(n_1489),
.C(n_1484),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1493),
.B(n_935),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1492),
.A2(n_1057),
.B(n_934),
.Y(n_1504)
);

NAND4xp75_ASAP7_75t_L g1505 ( 
.A(n_1480),
.B(n_1057),
.C(n_935),
.D(n_934),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1480),
.A2(n_873),
.B1(n_884),
.B2(n_886),
.Y(n_1506)
);

NAND2xp33_ASAP7_75t_L g1507 ( 
.A(n_1487),
.B(n_886),
.Y(n_1507)
);

AND4x1_ASAP7_75t_L g1508 ( 
.A(n_1498),
.B(n_891),
.C(n_914),
.D(n_920),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1496),
.B(n_920),
.Y(n_1509)
);

NAND4xp75_ASAP7_75t_L g1510 ( 
.A(n_1497),
.B(n_1500),
.C(n_1495),
.D(n_1499),
.Y(n_1510)
);

NAND4xp75_ASAP7_75t_L g1511 ( 
.A(n_1502),
.B(n_914),
.C(n_920),
.D(n_912),
.Y(n_1511)
);

NOR2x1_ASAP7_75t_L g1512 ( 
.A(n_1501),
.B(n_907),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1501),
.B(n_914),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1507),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1503),
.B(n_1506),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1505),
.B(n_917),
.Y(n_1516)
);

XOR2xp5_ASAP7_75t_L g1517 ( 
.A(n_1504),
.B(n_902),
.Y(n_1517)
);

OAI221xp5_ASAP7_75t_SL g1518 ( 
.A1(n_1508),
.A2(n_912),
.B1(n_898),
.B2(n_897),
.C(n_902),
.Y(n_1518)
);

AOI322xp5_ASAP7_75t_L g1519 ( 
.A1(n_1513),
.A2(n_912),
.A3(n_898),
.B1(n_897),
.B2(n_943),
.C1(n_925),
.C2(n_932),
.Y(n_1519)
);

OAI322xp33_ASAP7_75t_L g1520 ( 
.A1(n_1514),
.A2(n_938),
.A3(n_931),
.B1(n_929),
.B2(n_927),
.C1(n_926),
.C2(n_924),
.Y(n_1520)
);

AOI221xp5_ASAP7_75t_L g1521 ( 
.A1(n_1509),
.A2(n_1515),
.B1(n_1516),
.B2(n_1517),
.C(n_1510),
.Y(n_1521)
);

NAND3xp33_ASAP7_75t_L g1522 ( 
.A(n_1512),
.B(n_1511),
.C(n_929),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1521),
.Y(n_1523)
);

XNOR2xp5_ASAP7_75t_L g1524 ( 
.A(n_1522),
.B(n_898),
.Y(n_1524)
);

NAND4xp75_ASAP7_75t_L g1525 ( 
.A(n_1518),
.B(n_897),
.C(n_931),
.D(n_927),
.Y(n_1525)
);

OR2x2_ASAP7_75t_SL g1526 ( 
.A(n_1520),
.B(n_949),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1523),
.A2(n_1519),
.B1(n_866),
.B2(n_926),
.Y(n_1527)
);

OAI31xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1524),
.A2(n_938),
.A3(n_924),
.B(n_916),
.Y(n_1528)
);

CKINVDCx16_ASAP7_75t_R g1529 ( 
.A(n_1526),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1529),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1527),
.Y(n_1531)
);

INVxp67_ASAP7_75t_L g1532 ( 
.A(n_1530),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1531),
.A2(n_1525),
.B1(n_1528),
.B2(n_873),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1532),
.B(n_1533),
.Y(n_1534)
);

OAI22x1_ASAP7_75t_L g1535 ( 
.A1(n_1534),
.A2(n_866),
.B1(n_908),
.B2(n_916),
.Y(n_1535)
);

OA331x2_ASAP7_75t_L g1536 ( 
.A1(n_1535),
.A2(n_917),
.A3(n_932),
.B1(n_943),
.B2(n_925),
.B3(n_949),
.C1(n_946),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1536),
.A2(n_793),
.B1(n_946),
.B2(n_798),
.Y(n_1537)
);

AOI211xp5_ASAP7_75t_L g1538 ( 
.A1(n_1537),
.A2(n_793),
.B(n_951),
.C(n_899),
.Y(n_1538)
);


endmodule