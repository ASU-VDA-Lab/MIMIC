module fake_jpeg_8705_n_256 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_36),
.B(n_20),
.Y(n_67)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_38),
.Y(n_63)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_60),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_34),
.B(n_33),
.C(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_50),
.B(n_56),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_30),
.B1(n_34),
.B2(n_26),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_55),
.B1(n_58),
.B2(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_23),
.B1(n_32),
.B2(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_23),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_17),
.B1(n_33),
.B2(n_24),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_23),
.B1(n_20),
.B2(n_22),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_66),
.B1(n_68),
.B2(n_31),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_18),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_0),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_67),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_32),
.B1(n_20),
.B2(n_29),
.Y(n_66)
);

HAxp5_ASAP7_75t_SL g68 ( 
.A(n_38),
.B(n_25),
.CON(n_68),
.SN(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_22),
.B1(n_29),
.B2(n_18),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_38),
.A2(n_29),
.B1(n_31),
.B2(n_35),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_35),
.B1(n_27),
.B2(n_31),
.Y(n_86)
);

OAI32xp33_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_28),
.A3(n_19),
.B1(n_31),
.B2(n_35),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_72),
.A2(n_49),
.B1(n_61),
.B2(n_51),
.Y(n_116)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

AO22x1_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_46),
.B1(n_44),
.B2(n_42),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_74),
.A2(n_42),
.B1(n_40),
.B2(n_62),
.Y(n_118)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_76),
.Y(n_95)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_82),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_24),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_25),
.Y(n_84)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_70),
.B1(n_55),
.B2(n_66),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_46),
.C(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_59),
.Y(n_101)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_92),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_90),
.A2(n_94),
.B1(n_57),
.B2(n_63),
.Y(n_96)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_91),
.A2(n_64),
.B1(n_54),
.B2(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_12),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_50),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_57),
.A2(n_35),
.B1(n_27),
.B2(n_19),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_96),
.A2(n_71),
.B1(n_92),
.B2(n_85),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_105),
.B1(n_113),
.B2(n_71),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_91),
.B1(n_89),
.B2(n_73),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_83),
.B(n_81),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_75),
.A2(n_64),
.B1(n_54),
.B2(n_47),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_70),
.B1(n_59),
.B2(n_53),
.Y(n_105)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_77),
.B(n_61),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_115),
.Y(n_126)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_78),
.A2(n_49),
.B1(n_64),
.B2(n_56),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_61),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_116),
.A2(n_118),
.B1(n_86),
.B2(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_51),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_117),
.B(n_119),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_74),
.A2(n_58),
.B(n_21),
.C(n_27),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_120),
.A2(n_125),
.B1(n_130),
.B2(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_131),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_134),
.B(n_110),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_83),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_76),
.B1(n_91),
.B2(n_72),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_141),
.B1(n_143),
.B2(n_99),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_81),
.B(n_88),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_139),
.B(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_82),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_116),
.B1(n_119),
.B2(n_96),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_89),
.B1(n_79),
.B2(n_81),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_143),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_147),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_119),
.B1(n_107),
.B2(n_110),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_145),
.A2(n_159),
.B1(n_165),
.B2(n_7),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_98),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_149),
.B(n_0),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_137),
.B(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_151),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_97),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_97),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_153),
.B(n_155),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_107),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_162),
.C(n_168),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_161),
.Y(n_169)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_104),
.C(n_108),
.Y(n_162)
);

OAI32xp33_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_108),
.A3(n_84),
.B1(n_80),
.B2(n_27),
.Y(n_163)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_9),
.A3(n_15),
.B1(n_14),
.B2(n_3),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_121),
.B(n_136),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_133),
.A2(n_98),
.B1(n_109),
.B2(n_19),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_166),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_98),
.C(n_1),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_133),
.C(n_143),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_175),
.C(n_177),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_155),
.A2(n_142),
.B1(n_139),
.B2(n_131),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_174),
.A2(n_178),
.B(n_180),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_141),
.C(n_120),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_130),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_123),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_183),
.B1(n_165),
.B2(n_150),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_164),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_180)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_167),
.A2(n_6),
.B1(n_13),
.B2(n_12),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_188),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_5),
.B1(n_13),
.B2(n_11),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_152),
.B1(n_168),
.B2(n_163),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_5),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_148),
.B1(n_161),
.B2(n_160),
.Y(n_190)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_175),
.A2(n_148),
.B1(n_144),
.B2(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_162),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_202),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_166),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_196),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_176),
.B(n_151),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_203),
.B1(n_206),
.B2(n_180),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_169),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_204),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_152),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_171),
.A2(n_156),
.B1(n_157),
.B2(n_144),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_187),
.A2(n_156),
.B(n_157),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_205),
.A2(n_178),
.B(n_189),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_184),
.A2(n_145),
.B1(n_1),
.B2(n_2),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_178),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_0),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_191),
.B(n_177),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_170),
.Y(n_214)
);

XNOR2x1_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_188),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_198),
.Y(n_228)
);

OAI22x1_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_182),
.B1(n_174),
.B2(n_185),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_217),
.A2(n_201),
.B1(n_197),
.B2(n_206),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_204),
.A2(n_207),
.B(n_198),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_221),
.Y(n_225)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_202),
.C(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_227),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_200),
.C(n_194),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_210),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_201),
.B1(n_199),
.B2(n_205),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_230),
.A2(n_217),
.B1(n_219),
.B2(n_213),
.Y(n_234)
);

INVxp67_ASAP7_75t_SL g231 ( 
.A(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_234),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_222),
.A2(n_218),
.B(n_209),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_229),
.C(n_228),
.Y(n_240)
);

NAND4xp25_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_220),
.C(n_6),
.D(n_3),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_237),
.Y(n_244)
);

OAI221xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_16),
.B1(n_4),
.B2(n_6),
.C(n_9),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_238),
.A2(n_11),
.B(n_2),
.Y(n_245)
);

NOR3xp33_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_224),
.C(n_234),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_233),
.A2(n_226),
.B1(n_227),
.B2(n_11),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_242),
.B(n_236),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_1),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_245),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_235),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_249),
.C(n_232),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_248),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_252),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_226),
.C(n_244),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_243),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_2),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_255),
.B(n_253),
.Y(n_256)
);


endmodule