module fake_jpeg_29847_n_117 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_117);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_117;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx13_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_5),
.B(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_0),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_62),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_1),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_2),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_1),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_44),
.B1(n_54),
.B2(n_53),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_53),
.B1(n_46),
.B2(n_54),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_73),
.B1(n_68),
.B2(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_71),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_48),
.B1(n_4),
.B2(n_5),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_6),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_2),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_52),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_51),
.B1(n_44),
.B2(n_49),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_48),
.B1(n_3),
.B2(n_4),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_50),
.B1(n_43),
.B2(n_44),
.Y(n_73)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_3),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_85),
.Y(n_100)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_80),
.B(n_8),
.Y(n_94)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_65),
.B(n_6),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_89),
.Y(n_99)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_68),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_90),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_93),
.B1(n_29),
.B2(n_31),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_71),
.B1(n_10),
.B2(n_11),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_97),
.B1(n_98),
.B2(n_28),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_38),
.B1(n_24),
.B2(n_13),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_95),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_11),
.B(n_16),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_33),
.B(n_36),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_20),
.B1(n_22),
.B2(n_25),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_96),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_101),
.B(n_106),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_26),
.B(n_27),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_105),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_99),
.C(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_108),
.B(n_102),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

AOI21x1_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_103),
.B(n_109),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_106),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_93),
.C(n_110),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_115),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_104),
.Y(n_117)
);


endmodule