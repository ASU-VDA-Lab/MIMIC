module fake_jpeg_3605_n_601 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_601);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_601;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_55),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_58),
.Y(n_181)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_62),
.Y(n_157)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

CKINVDCx6p67_ASAP7_75t_R g150 ( 
.A(n_63),
.Y(n_150)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_52),
.Y(n_64)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_64),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_68),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_69),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_70),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_71),
.Y(n_202)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_72),
.Y(n_170)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_73),
.Y(n_178)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_75),
.Y(n_185)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g132 ( 
.A(n_76),
.Y(n_132)
);

BUFx4f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g176 ( 
.A(n_78),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_79),
.B(n_96),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_0),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_80),
.B(n_86),
.Y(n_141)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g211 ( 
.A(n_82),
.Y(n_211)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_0),
.Y(n_86)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_88),
.Y(n_195)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_89),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_92),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_93),
.Y(n_210)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_94),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_95),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_35),
.B(n_0),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_97),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_98),
.Y(n_194)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_100),
.Y(n_198)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_101),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_102),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_37),
.B(n_0),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_103),
.B(n_51),
.Y(n_167)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_20),
.Y(n_105)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_105),
.Y(n_205)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_28),
.Y(n_107)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_35),
.B(n_44),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_118),
.Y(n_156)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_39),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_39),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_112),
.B(n_114),
.Y(n_173)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_29),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_43),
.Y(n_116)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_29),
.Y(n_117)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_40),
.B(n_16),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_29),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_119),
.B(n_47),
.Y(n_175)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_120),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_19),
.Y(n_123)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_123),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_38),
.Y(n_124)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_43),
.Y(n_125)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_125),
.Y(n_184)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_41),
.B1(n_45),
.B2(n_48),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_129),
.A2(n_130),
.B1(n_144),
.B2(n_154),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_58),
.A2(n_26),
.B1(n_31),
.B2(n_50),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_75),
.A2(n_26),
.B1(n_31),
.B2(n_50),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_102),
.A2(n_41),
.B1(n_45),
.B2(n_48),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_151),
.A2(n_164),
.B1(n_169),
.B2(n_187),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_77),
.A2(n_26),
.B1(n_31),
.B2(n_50),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_103),
.A2(n_40),
.B1(n_44),
.B2(n_41),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_90),
.A2(n_50),
.B1(n_45),
.B2(n_48),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_165),
.A2(n_166),
.B1(n_182),
.B2(n_197),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_85),
.A2(n_113),
.B1(n_63),
.B2(n_21),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_175),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_124),
.A2(n_36),
.B1(n_21),
.B2(n_51),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_64),
.B(n_49),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_172),
.B(n_179),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_49),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_201),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_62),
.B(n_47),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_107),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_121),
.A2(n_25),
.B1(n_24),
.B2(n_34),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_65),
.B(n_1),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_200),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_122),
.A2(n_54),
.B1(n_53),
.B2(n_34),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_66),
.B(n_1),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_69),
.B(n_1),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_70),
.B(n_54),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_203),
.B(n_215),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_71),
.B(n_34),
.C(n_20),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_204),
.B(n_154),
.C(n_130),
.Y(n_275)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_78),
.B(n_53),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_207),
.B(n_214),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_82),
.B(n_1),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_2),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_84),
.A2(n_53),
.B(n_46),
.C(n_5),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_91),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_92),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_129),
.A2(n_98),
.B1(n_97),
.B2(n_95),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_218),
.A2(n_237),
.B1(n_269),
.B2(n_271),
.Y(n_319)
);

OAI32xp33_ASAP7_75t_L g220 ( 
.A1(n_141),
.A2(n_93),
.A3(n_46),
.B1(n_5),
.B2(n_6),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_220),
.A2(n_246),
.B(n_166),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_150),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_221),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_222),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_181),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_223),
.B(n_248),
.Y(n_299)
);

INVx11_ASAP7_75t_L g224 ( 
.A(n_150),
.Y(n_224)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_224),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_225),
.B(n_249),
.Y(n_297)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_177),
.Y(n_226)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_226),
.Y(n_293)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_228),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_156),
.B(n_2),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_229),
.B(n_234),
.Y(n_324)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_147),
.Y(n_230)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_230),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_165),
.A2(n_46),
.B1(n_3),
.B2(n_6),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_231),
.A2(n_236),
.B1(n_282),
.B2(n_157),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_150),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_232),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_175),
.A2(n_46),
.B1(n_3),
.B2(n_6),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_233),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_143),
.B(n_2),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_L g236 ( 
.A1(n_182),
.A2(n_46),
.B1(n_8),
.B2(n_9),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_159),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_138),
.Y(n_238)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_238),
.Y(n_294)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_161),
.Y(n_239)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_239),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_173),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_240),
.A2(n_244),
.B1(n_254),
.B2(n_257),
.Y(n_298)
);

BUFx2_ASAP7_75t_SL g241 ( 
.A(n_212),
.Y(n_241)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_241),
.Y(n_307)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_142),
.Y(n_242)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_242),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_173),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_244)
);

BUFx4f_ASAP7_75t_L g245 ( 
.A(n_198),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g344 ( 
.A(n_245),
.Y(n_344)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_203),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_183),
.Y(n_247)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_247),
.Y(n_312)
);

AND2x2_ASAP7_75t_SL g248 ( 
.A(n_184),
.B(n_14),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_180),
.B(n_14),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_171),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_250),
.B(n_279),
.Y(n_303)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_132),
.Y(n_251)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_251),
.Y(n_316)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_135),
.Y(n_252)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_252),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_158),
.A2(n_16),
.B1(n_131),
.B2(n_212),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_196),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_255),
.B(n_275),
.Y(n_338)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_128),
.Y(n_256)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_256),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_158),
.A2(n_136),
.B1(n_190),
.B2(n_186),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_157),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_258),
.Y(n_317)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_132),
.Y(n_259)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_259),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_207),
.B(n_191),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_260),
.B(n_261),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_145),
.B(n_149),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_176),
.Y(n_262)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_262),
.Y(n_325)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_213),
.Y(n_263)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_263),
.Y(n_328)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_127),
.Y(n_264)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_264),
.Y(n_337)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_176),
.Y(n_266)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_266),
.Y(n_347)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_160),
.Y(n_267)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_267),
.Y(n_332)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_139),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_268),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_170),
.A2(n_178),
.B1(n_152),
.B2(n_188),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_168),
.A2(n_148),
.B1(n_205),
.B2(n_162),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_211),
.Y(n_272)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_272),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_163),
.B(n_198),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_273),
.B(n_276),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_209),
.B(n_189),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_148),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_277),
.Y(n_308)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_211),
.Y(n_278)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_278),
.Y(n_336)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_195),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_209),
.B(n_189),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_280),
.B(n_140),
.Y(n_315)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_153),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_284),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_144),
.A2(n_133),
.B1(n_134),
.B2(n_192),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_194),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_283),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_206),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_196),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_287),
.Y(n_310)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_133),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_171),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_289),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_137),
.B(n_199),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_134),
.A2(n_202),
.B1(n_146),
.B2(n_192),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_290),
.A2(n_276),
.B1(n_280),
.B2(n_258),
.Y(n_333)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_194),
.Y(n_291)
);

NOR2x1_ASAP7_75t_R g305 ( 
.A(n_291),
.B(n_210),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_265),
.A2(n_274),
.B1(n_270),
.B2(n_243),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_301),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_302),
.A2(n_311),
.B1(n_313),
.B2(n_314),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_305),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_253),
.A2(n_146),
.B1(n_202),
.B2(n_155),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_253),
.A2(n_265),
.B1(n_285),
.B2(n_217),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_315),
.B(n_262),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_265),
.A2(n_155),
.B1(n_199),
.B2(n_210),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_329),
.A2(n_345),
.B1(n_259),
.B2(n_251),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_260),
.A2(n_137),
.B1(n_140),
.B2(n_282),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_330),
.A2(n_343),
.B1(n_223),
.B2(n_224),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g331 ( 
.A(n_273),
.B(n_261),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_331),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_333),
.A2(n_331),
.B1(n_334),
.B2(n_326),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_221),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_340),
.B(n_283),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_231),
.A2(n_275),
.B1(n_236),
.B2(n_249),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_217),
.A2(n_220),
.B1(n_234),
.B2(n_248),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_246),
.A2(n_219),
.B(n_227),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_346),
.A2(n_235),
.B(n_226),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_294),
.B(n_232),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_219),
.C(n_252),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_354),
.C(n_385),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_301),
.A2(n_248),
.B1(n_225),
.B2(n_219),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_352),
.A2(n_353),
.B1(n_355),
.B2(n_378),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_229),
.C(n_228),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_296),
.B(n_255),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_356),
.Y(n_405)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_357),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_334),
.A2(n_279),
.B1(n_267),
.B2(n_283),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_358),
.Y(n_417)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_310),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_359),
.B(n_363),
.Y(n_418)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_322),
.Y(n_360)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_360),
.Y(n_408)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_335),
.Y(n_361)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_361),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_362),
.B(n_364),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_314),
.B(n_239),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_339),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_338),
.A2(n_247),
.B(n_250),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_365),
.Y(n_411)
);

A2O1A1O1Ixp25_ASAP7_75t_L g366 ( 
.A1(n_341),
.A2(n_291),
.B(n_230),
.C(n_287),
.D(n_266),
.Y(n_366)
);

XOR2x1_ASAP7_75t_SL g424 ( 
.A(n_366),
.B(n_292),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_368),
.Y(n_392)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_332),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_369),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_370),
.B(n_304),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_313),
.A2(n_272),
.B1(n_278),
.B2(n_245),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_371),
.A2(n_376),
.B1(n_379),
.B2(n_383),
.Y(n_402)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_332),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_372),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_309),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_373),
.B(n_374),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_327),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_335),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_375),
.B(n_377),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_302),
.A2(n_245),
.B1(n_343),
.B2(n_345),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_297),
.B(n_324),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_311),
.A2(n_323),
.B1(n_315),
.B2(n_330),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_331),
.A2(n_323),
.B1(n_329),
.B2(n_319),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_331),
.A2(n_324),
.B1(n_299),
.B2(n_298),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_380),
.A2(n_352),
.B1(n_348),
.B2(n_365),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_336),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_381),
.Y(n_393)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_318),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_387),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_299),
.B(n_306),
.C(n_295),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_317),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_386),
.Y(n_396)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_304),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_299),
.B(n_308),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_389),
.Y(n_416)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_344),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_303),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_390),
.A2(n_366),
.B1(n_373),
.B2(n_362),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_348),
.A2(n_346),
.B1(n_295),
.B2(n_305),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_400),
.A2(n_424),
.B(n_307),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_351),
.B(n_337),
.C(n_328),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_403),
.B(n_414),
.C(n_420),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_376),
.A2(n_320),
.B1(n_317),
.B2(n_316),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_404),
.A2(n_406),
.B1(n_357),
.B2(n_360),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_349),
.A2(n_321),
.B1(n_316),
.B2(n_336),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_407),
.A2(n_413),
.B1(n_415),
.B2(n_422),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_374),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_409),
.B(n_425),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_349),
.A2(n_321),
.B1(n_347),
.B2(n_325),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_370),
.B(n_293),
.C(n_312),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_378),
.A2(n_379),
.B1(n_355),
.B2(n_384),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_384),
.B(n_293),
.C(n_312),
.Y(n_420)
);

OA21x2_ASAP7_75t_L g421 ( 
.A1(n_353),
.A2(n_344),
.B(n_307),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_421),
.B(n_389),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_364),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_426),
.B(n_382),
.Y(n_447)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_428),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_401),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_429),
.B(n_435),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_405),
.B(n_390),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_430),
.B(n_441),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_402),
.A2(n_415),
.B1(n_419),
.B2(n_404),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_432),
.A2(n_449),
.B1(n_457),
.B2(n_396),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_391),
.B(n_354),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_436),
.Y(n_467)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_399),
.Y(n_434)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_434),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_419),
.A2(n_367),
.B1(n_380),
.B2(n_388),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_391),
.B(n_426),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_403),
.B(n_385),
.C(n_361),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_437),
.B(n_439),
.C(n_410),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_402),
.A2(n_367),
.B(n_292),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_438),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_377),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_413),
.A2(n_371),
.B1(n_358),
.B2(n_375),
.Y(n_440)
);

AO21x2_ASAP7_75t_L g487 ( 
.A1(n_440),
.A2(n_442),
.B(n_445),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_397),
.B(n_318),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_411),
.A2(n_394),
.B1(n_400),
.B2(n_412),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_444),
.B(n_453),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_421),
.A2(n_386),
.B1(n_372),
.B2(n_369),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_394),
.B(n_387),
.Y(n_446)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_446),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_447),
.B(n_414),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_395),
.B(n_342),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_448),
.B(n_451),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_406),
.A2(n_421),
.B1(n_411),
.B2(n_418),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_398),
.Y(n_450)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_450),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_395),
.B(n_342),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_452),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_418),
.A2(n_386),
.B1(n_325),
.B2(n_347),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_454),
.B(n_438),
.Y(n_474)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_408),
.Y(n_455)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_455),
.Y(n_486)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_408),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_456),
.B(n_458),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_421),
.A2(n_300),
.B1(n_344),
.B2(n_392),
.Y(n_457)
);

OAI32xp33_ASAP7_75t_L g458 ( 
.A1(n_416),
.A2(n_300),
.A3(n_417),
.B1(n_424),
.B2(n_420),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_416),
.A2(n_392),
.B(n_417),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_459),
.B(n_410),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_460),
.B(n_461),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_439),
.B(n_423),
.Y(n_461)
);

AOI22x1_ASAP7_75t_L g463 ( 
.A1(n_442),
.A2(n_409),
.B1(n_425),
.B2(n_401),
.Y(n_463)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_463),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_433),
.B(n_423),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_465),
.B(n_466),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_436),
.B(n_393),
.Y(n_466)
);

XNOR2x2_ASAP7_75t_SL g468 ( 
.A(n_459),
.B(n_446),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_468),
.B(n_472),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_393),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_469),
.B(n_488),
.C(n_444),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_470),
.A2(n_474),
.B(n_434),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_443),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_477),
.B(n_479),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_443),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_445),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_480),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_437),
.B(n_398),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_435),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_484),
.A2(n_396),
.B1(n_410),
.B2(n_450),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_431),
.B(n_447),
.C(n_427),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_491),
.B(n_492),
.C(n_498),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_467),
.B(n_454),
.Y(n_492)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_493),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_470),
.Y(n_494)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_494),
.Y(n_517)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_473),
.Y(n_497)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_497),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_467),
.B(n_432),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_469),
.B(n_429),
.C(n_449),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_500),
.B(n_506),
.C(n_488),
.Y(n_529)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_489),
.Y(n_502)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_502),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_487),
.A2(n_457),
.B1(n_428),
.B2(n_458),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_503),
.B(n_513),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_475),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_504),
.B(n_507),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_456),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_505),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_466),
.B(n_455),
.C(n_452),
.Y(n_506)
);

INVx6_ASAP7_75t_L g507 ( 
.A(n_468),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_463),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_508),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_509),
.B(n_471),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_478),
.A2(n_440),
.B(n_453),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_510),
.A2(n_478),
.B(n_485),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_512),
.A2(n_487),
.B1(n_463),
.B2(n_483),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_476),
.B(n_398),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_462),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_514),
.B(n_481),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_461),
.B(n_472),
.Y(n_515)
);

XNOR2x1_ASAP7_75t_L g528 ( 
.A(n_515),
.B(n_495),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_520),
.A2(n_522),
.B(n_523),
.Y(n_538)
);

AOI21x1_ASAP7_75t_L g522 ( 
.A1(n_511),
.A2(n_485),
.B(n_487),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_511),
.A2(n_471),
.B(n_476),
.Y(n_523)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_527),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_528),
.B(n_529),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_531),
.A2(n_509),
.B(n_510),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_532),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_507),
.A2(n_487),
.B1(n_483),
.B2(n_484),
.Y(n_533)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_533),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_499),
.B(n_505),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_534),
.A2(n_490),
.B1(n_465),
.B2(n_492),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_501),
.B(n_486),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_535),
.B(n_536),
.Y(n_547)
);

FAx1_ASAP7_75t_SL g536 ( 
.A(n_500),
.B(n_490),
.CI(n_495),
.CON(n_536),
.SN(n_536)
);

INVxp33_ASAP7_75t_SL g537 ( 
.A(n_534),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_537),
.B(n_539),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_529),
.B(n_491),
.C(n_498),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_541),
.B(n_545),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_524),
.B(n_496),
.C(n_506),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_544),
.B(n_548),
.C(n_550),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_518),
.B(n_464),
.Y(n_546)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_546),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_524),
.B(n_496),
.C(n_515),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_516),
.A2(n_487),
.B1(n_512),
.B2(n_513),
.Y(n_549)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_549),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_528),
.B(n_460),
.C(n_503),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_520),
.B(n_531),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_551),
.B(n_522),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_552),
.A2(n_516),
.B1(n_542),
.B2(n_517),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_553),
.B(n_559),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_555),
.B(n_521),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_551),
.B(n_533),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_558),
.B(n_564),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_544),
.B(n_519),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_539),
.B(n_523),
.C(n_521),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_561),
.B(n_563),
.Y(n_574)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_543),
.Y(n_562)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_562),
.Y(n_575)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_549),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_547),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_547),
.B(n_518),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_566),
.B(n_527),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_565),
.A2(n_519),
.B(n_548),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_567),
.A2(n_572),
.B(n_555),
.Y(n_583)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_570),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_559),
.B(n_542),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_571),
.B(n_576),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_560),
.A2(n_538),
.B(n_552),
.Y(n_572)
);

A2O1A1Ixp33_ASAP7_75t_SL g581 ( 
.A1(n_573),
.A2(n_565),
.B(n_553),
.C(n_517),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_561),
.B(n_540),
.C(n_550),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_558),
.B(n_540),
.C(n_538),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_577),
.B(n_557),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_569),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_578),
.A2(n_584),
.B1(n_575),
.B2(n_525),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_576),
.B(n_554),
.Y(n_580)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_580),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_581),
.B(n_582),
.Y(n_590)
);

NOR2xp67_ASAP7_75t_L g582 ( 
.A(n_574),
.B(n_554),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_583),
.B(n_585),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_568),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_586),
.B(n_556),
.Y(n_587)
);

AOI21x1_ASAP7_75t_SL g593 ( 
.A1(n_587),
.A2(n_535),
.B(n_523),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_579),
.B(n_577),
.C(n_573),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_SL g594 ( 
.A1(n_589),
.A2(n_525),
.B(n_532),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_SL g595 ( 
.A1(n_591),
.A2(n_526),
.B(n_530),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_593),
.B(n_594),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_595),
.B(n_592),
.C(n_590),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_596),
.A2(n_587),
.B(n_588),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_598),
.B(n_597),
.C(n_526),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_L g600 ( 
.A1(n_599),
.A2(n_530),
.B(n_536),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_600),
.B(n_536),
.Y(n_601)
);


endmodule