module fake_aes_6391_n_724 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_724);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_724;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_472;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_60), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_50), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_22), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_59), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_31), .Y(n_84) );
BUFx2_ASAP7_75t_SL g85 ( .A(n_2), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_12), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_2), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_18), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_41), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_73), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_7), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_25), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_57), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_14), .Y(n_94) );
BUFx2_ASAP7_75t_L g95 ( .A(n_19), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_66), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_36), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_58), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_1), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_27), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_77), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_74), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_20), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_61), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_21), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_39), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_44), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_20), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_14), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_40), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_32), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_62), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_3), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_6), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_4), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_65), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_63), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_37), .Y(n_118) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_30), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_55), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_46), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_52), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_8), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_42), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g125 ( .A(n_38), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_48), .Y(n_126) );
INVx1_ASAP7_75t_SL g127 ( .A(n_49), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_69), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_34), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_95), .B(n_0), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_87), .B(n_0), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_95), .B(n_1), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_87), .B(n_3), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_84), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_99), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_89), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_89), .Y(n_138) );
INVx4_ASAP7_75t_L g139 ( .A(n_96), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_90), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_90), .Y(n_141) );
BUFx8_ASAP7_75t_L g142 ( .A(n_92), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_92), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_93), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_93), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_99), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_98), .Y(n_147) );
BUFx2_ASAP7_75t_L g148 ( .A(n_114), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_98), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_129), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_100), .Y(n_151) );
INVx5_ASAP7_75t_L g152 ( .A(n_101), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_100), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_124), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_83), .B(n_4), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_126), .B(n_5), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_80), .B(n_5), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_124), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_129), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_128), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_128), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_125), .B(n_6), .Y(n_162) );
AND2x2_ASAP7_75t_SL g163 ( .A(n_81), .B(n_79), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_104), .Y(n_164) );
BUFx8_ASAP7_75t_L g165 ( .A(n_106), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_107), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_110), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_111), .Y(n_168) );
NAND2x1p5_ASAP7_75t_L g169 ( .A(n_86), .B(n_33), .Y(n_169) );
INVxp67_ASAP7_75t_L g170 ( .A(n_86), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_112), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_82), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_148), .B(n_114), .Y(n_173) );
OR2x2_ASAP7_75t_L g174 ( .A(n_148), .B(n_123), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_139), .B(n_123), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_131), .Y(n_176) );
AND3x1_ASAP7_75t_L g177 ( .A(n_130), .B(n_94), .C(n_88), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_131), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_139), .B(n_116), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_131), .Y(n_180) );
INVx1_ASAP7_75t_SL g181 ( .A(n_136), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_139), .B(n_121), .Y(n_182) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_136), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_139), .B(n_117), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_152), .B(n_97), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_152), .B(n_97), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_171), .B(n_122), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_131), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_171), .B(n_122), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_133), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_133), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_133), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_149), .Y(n_194) );
INVx4_ASAP7_75t_SL g195 ( .A(n_160), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_152), .B(n_96), .Y(n_196) );
INVx2_ASAP7_75t_SL g197 ( .A(n_152), .Y(n_197) );
NOR2xp33_ASAP7_75t_SL g198 ( .A(n_142), .B(n_120), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_149), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_170), .B(n_118), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_146), .B(n_118), .Y(n_201) );
AND2x6_ASAP7_75t_L g202 ( .A(n_133), .B(n_94), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_149), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_130), .B(n_88), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_145), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_145), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_152), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_149), .Y(n_208) );
AND2x6_ASAP7_75t_L g209 ( .A(n_145), .B(n_91), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_145), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_170), .B(n_102), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_149), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_134), .B(n_91), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_149), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_137), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_152), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_150), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_150), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_160), .B(n_127), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_150), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_137), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_150), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_137), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_142), .Y(n_224) );
INVx6_ASAP7_75t_L g225 ( .A(n_167), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_172), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_146), .B(n_108), .Y(n_227) );
INVxp67_ASAP7_75t_SL g228 ( .A(n_132), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_134), .B(n_119), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_135), .B(n_113), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_135), .B(n_115), .Y(n_231) );
INVx4_ASAP7_75t_L g232 ( .A(n_169), .Y(n_232) );
AOI22x1_ASAP7_75t_L g233 ( .A1(n_169), .A2(n_109), .B1(n_105), .B2(n_103), .Y(n_233) );
NOR2x1p5_ASAP7_75t_L g234 ( .A(n_132), .B(n_85), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_150), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_138), .B(n_85), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_138), .B(n_7), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_141), .B(n_35), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_162), .B(n_8), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_228), .B(n_142), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_200), .B(n_142), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_181), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_237), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_177), .A2(n_163), .B1(n_162), .B2(n_165), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_205), .Y(n_245) );
AND2x6_ASAP7_75t_L g246 ( .A(n_224), .B(n_160), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_183), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_200), .B(n_165), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_225), .Y(n_249) );
BUFx2_ASAP7_75t_L g250 ( .A(n_174), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_224), .B(n_163), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_237), .Y(n_252) );
OR2x6_ASAP7_75t_L g253 ( .A(n_232), .B(n_169), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_187), .B(n_165), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_237), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_187), .B(n_165), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_213), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_189), .B(n_161), .Y(n_258) );
INVxp67_ASAP7_75t_L g259 ( .A(n_173), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_209), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_209), .Y(n_261) );
AND2x4_ASAP7_75t_SL g262 ( .A(n_232), .B(n_151), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_213), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_175), .B(n_155), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_213), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_225), .Y(n_266) );
BUFx8_ASAP7_75t_L g267 ( .A(n_201), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_202), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_232), .B(n_163), .Y(n_269) );
INVxp67_ASAP7_75t_SL g270 ( .A(n_193), .Y(n_270) );
INVx4_ASAP7_75t_L g271 ( .A(n_195), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_234), .B(n_155), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_202), .A2(n_156), .B1(n_157), .B2(n_154), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_204), .B(n_156), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_193), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_193), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_176), .Y(n_277) );
INVx5_ASAP7_75t_L g278 ( .A(n_209), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_202), .A2(n_147), .B1(n_141), .B2(n_161), .Y(n_279) );
OR2x4_ASAP7_75t_L g280 ( .A(n_227), .B(n_236), .Y(n_280) );
INVx2_ASAP7_75t_SL g281 ( .A(n_204), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_189), .B(n_151), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_178), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_180), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_202), .Y(n_285) );
BUFx4f_ASAP7_75t_L g286 ( .A(n_202), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_188), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_211), .B(n_154), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_211), .B(n_147), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_190), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_204), .B(n_164), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_191), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_226), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_209), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_231), .B(n_164), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_209), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_192), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_231), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_206), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_179), .B(n_164), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_179), .B(n_166), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_233), .B(n_153), .Y(n_302) );
BUFx4f_ASAP7_75t_L g303 ( .A(n_239), .Y(n_303) );
NAND2x1p5_ASAP7_75t_L g304 ( .A(n_231), .B(n_166), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_226), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_210), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_195), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_236), .B(n_166), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_182), .B(n_140), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_219), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_182), .B(n_140), .Y(n_311) );
AND2x6_ASAP7_75t_L g312 ( .A(n_285), .B(n_192), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_242), .Y(n_313) );
NAND2x1p5_ASAP7_75t_L g314 ( .A(n_285), .B(n_215), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_269), .A2(n_229), .B1(n_184), .B2(n_219), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_274), .B(n_229), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_247), .Y(n_317) );
BUFx12f_ASAP7_75t_L g318 ( .A(n_267), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_275), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g320 ( .A(n_293), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_246), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g322 ( .A(n_278), .B(n_195), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_245), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_305), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_276), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_262), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_246), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_240), .A2(n_185), .B(n_186), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_269), .A2(n_184), .B1(n_221), .B2(n_223), .Y(n_329) );
INVx2_ASAP7_75t_SL g330 ( .A(n_262), .Y(n_330) );
BUFx4_ASAP7_75t_R g331 ( .A(n_267), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_245), .Y(n_332) );
INVx2_ASAP7_75t_SL g333 ( .A(n_246), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_260), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_246), .Y(n_335) );
OAI22xp5_ASAP7_75t_SL g336 ( .A1(n_244), .A2(n_230), .B1(n_198), .B2(n_140), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_299), .Y(n_337) );
BUFx12f_ASAP7_75t_L g338 ( .A(n_250), .Y(n_338) );
AOI22x1_ASAP7_75t_L g339 ( .A1(n_252), .A2(n_220), .B1(n_235), .B2(n_194), .Y(n_339) );
BUFx12f_ASAP7_75t_L g340 ( .A(n_253), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_259), .B(n_143), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_306), .Y(n_342) );
INVx3_ASAP7_75t_L g343 ( .A(n_260), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_264), .B(n_196), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_297), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_264), .B(n_143), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_297), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_304), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_270), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_246), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_270), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_243), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_260), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_304), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_253), .Y(n_355) );
INVx5_ASAP7_75t_L g356 ( .A(n_260), .Y(n_356) );
NAND2x1p5_ASAP7_75t_L g357 ( .A(n_286), .B(n_216), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_261), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_298), .B(n_143), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_259), .B(n_144), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_298), .B(n_144), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_277), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_251), .A2(n_238), .B1(n_167), .B2(n_168), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_243), .Y(n_364) );
BUFx8_ASAP7_75t_L g365 ( .A(n_261), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_283), .Y(n_366) );
AND2x6_ASAP7_75t_L g367 ( .A(n_321), .B(n_261), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_336), .A2(n_251), .B1(n_272), .B2(n_281), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_341), .A2(n_255), .B1(n_279), .B2(n_273), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_341), .Y(n_370) );
NAND3xp33_ASAP7_75t_SL g371 ( .A(n_313), .B(n_254), .C(n_256), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_334), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_336), .A2(n_272), .B1(n_253), .B2(n_303), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_328), .A2(n_258), .B(n_282), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_317), .Y(n_375) );
O2A1O1Ixp33_ASAP7_75t_SL g376 ( .A1(n_333), .A2(n_302), .B(n_241), .C(n_248), .Y(n_376) );
OAI21xp5_ASAP7_75t_L g377 ( .A1(n_344), .A2(n_311), .B(n_300), .Y(n_377) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_316), .A2(n_291), .B1(n_289), .B2(n_288), .C(n_301), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_323), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g380 ( .A1(n_340), .A2(n_303), .B1(n_286), .B2(n_268), .Y(n_380) );
AOI22xp33_ASAP7_75t_SL g381 ( .A1(n_340), .A2(n_268), .B1(n_310), .B2(n_257), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_338), .Y(n_382) );
OR2x6_ASAP7_75t_L g383 ( .A(n_326), .B(n_261), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_349), .A2(n_265), .B1(n_263), .B2(n_292), .Y(n_384) );
AOI22xp33_ASAP7_75t_SL g385 ( .A1(n_355), .A2(n_295), .B1(n_301), .B2(n_300), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_360), .B(n_280), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_SL g387 ( .A1(n_333), .A2(n_302), .B(n_366), .C(n_362), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g388 ( .A1(n_362), .A2(n_311), .B(n_308), .C(n_309), .Y(n_388) );
INVxp33_ASAP7_75t_L g389 ( .A(n_348), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_360), .B(n_280), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_359), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_354), .B(n_278), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_323), .Y(n_393) );
AO21x2_ASAP7_75t_L g394 ( .A1(n_366), .A2(n_238), .B(n_158), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_346), .A2(n_287), .B1(n_290), .B2(n_284), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_332), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_354), .B(n_294), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_359), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_326), .B(n_278), .Y(n_399) );
INVx3_ASAP7_75t_L g400 ( .A(n_367), .Y(n_400) );
OAI22xp33_ASAP7_75t_L g401 ( .A1(n_375), .A2(n_355), .B1(n_338), .B2(n_318), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_385), .A2(n_318), .B1(n_337), .B2(n_315), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_379), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_386), .B(n_324), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_377), .B(n_342), .Y(n_405) );
OAI21xp33_ASAP7_75t_L g406 ( .A1(n_388), .A2(n_329), .B(n_363), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_390), .A2(n_324), .B1(n_359), .B2(n_337), .C(n_342), .Y(n_407) );
INVx4_ASAP7_75t_L g408 ( .A(n_367), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_388), .B(n_349), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_379), .B(n_342), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_373), .A2(n_359), .B1(n_330), .B2(n_320), .Y(n_411) );
INVx3_ASAP7_75t_L g412 ( .A(n_367), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_368), .A2(n_330), .B1(n_352), .B2(n_364), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_389), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_371), .A2(n_352), .B1(n_364), .B2(n_325), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_393), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_395), .A2(n_351), .B1(n_332), .B2(n_321), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_378), .A2(n_158), .B1(n_144), .B2(n_351), .C(n_361), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_393), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_370), .A2(n_364), .B1(n_325), .B2(n_319), .Y(n_420) );
AO21x2_ASAP7_75t_L g421 ( .A1(n_376), .A2(n_158), .B(n_319), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_369), .A2(n_321), .B1(n_327), .B2(n_335), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_374), .B(n_347), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_382), .A2(n_327), .B1(n_335), .B2(n_350), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_396), .Y(n_425) );
A2O1A1Ixp33_ASAP7_75t_L g426 ( .A1(n_384), .A2(n_350), .B(n_347), .C(n_345), .Y(n_426) );
AO31x2_ASAP7_75t_L g427 ( .A1(n_396), .A2(n_347), .A3(n_194), .B(n_214), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_392), .B(n_356), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_410), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_403), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_403), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_410), .B(n_394), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_419), .B(n_394), .Y(n_433) );
AO21x2_ASAP7_75t_L g434 ( .A1(n_423), .A2(n_376), .B(n_387), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_408), .B(n_372), .Y(n_435) );
OAI321xp33_ASAP7_75t_L g436 ( .A1(n_402), .A2(n_398), .A3(n_391), .B1(n_383), .B2(n_168), .C(n_167), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_407), .A2(n_389), .B1(n_159), .B2(n_153), .C(n_150), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_419), .B(n_394), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_425), .B(n_397), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_411), .A2(n_381), .B1(n_380), .B2(n_397), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_425), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_401), .A2(n_153), .B1(n_159), .B2(n_167), .C(n_168), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_405), .B(n_392), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_416), .Y(n_444) );
AOI211xp5_ASAP7_75t_SL g445 ( .A1(n_417), .A2(n_331), .B(n_387), .C(n_399), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_416), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_417), .A2(n_409), .B1(n_415), .B2(n_405), .Y(n_447) );
BUFx3_ASAP7_75t_L g448 ( .A(n_428), .Y(n_448) );
BUFx2_ASAP7_75t_L g449 ( .A(n_416), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_409), .A2(n_372), .B(n_334), .Y(n_450) );
OA21x2_ASAP7_75t_L g451 ( .A1(n_423), .A2(n_339), .B(n_214), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_408), .B(n_372), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_427), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_404), .A2(n_153), .B1(n_159), .B2(n_167), .C(n_168), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_422), .A2(n_383), .B1(n_314), .B2(n_372), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_427), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_427), .Y(n_457) );
NAND4xp25_ASAP7_75t_L g458 ( .A(n_420), .B(n_220), .C(n_235), .D(n_11), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_406), .A2(n_353), .B(n_334), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_428), .B(n_413), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_421), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_427), .Y(n_462) );
OAI22xp5_ASAP7_75t_SL g463 ( .A1(n_414), .A2(n_383), .B1(n_314), .B2(n_392), .Y(n_463) );
BUFx2_ASAP7_75t_L g464 ( .A(n_408), .Y(n_464) );
NAND4xp25_ASAP7_75t_SL g465 ( .A(n_424), .B(n_9), .C(n_10), .D(n_11), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_435), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g467 ( .A(n_442), .B(n_168), .C(n_167), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_429), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_430), .Y(n_469) );
OAI33xp33_ASAP7_75t_L g470 ( .A1(n_458), .A2(n_406), .A3(n_10), .B1(n_12), .B2(n_13), .B3(n_15), .Y(n_470) );
OAI22xp5_ASAP7_75t_SL g471 ( .A1(n_463), .A2(n_408), .B1(n_428), .B2(n_412), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_449), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_458), .A2(n_418), .B1(n_428), .B2(n_400), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_449), .B(n_427), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_432), .B(n_421), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_439), .Y(n_476) );
INVx3_ASAP7_75t_L g477 ( .A(n_435), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_431), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_431), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_441), .Y(n_480) );
AO31x2_ASAP7_75t_L g481 ( .A1(n_447), .A2(n_426), .A3(n_421), .B(n_345), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_448), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_448), .Y(n_483) );
AO21x2_ASAP7_75t_L g484 ( .A1(n_459), .A2(n_421), .B(n_322), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g485 ( .A1(n_465), .A2(n_418), .B1(n_168), .B2(n_159), .C(n_153), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_446), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_439), .B(n_153), .Y(n_487) );
INVx4_ASAP7_75t_L g488 ( .A(n_464), .Y(n_488) );
AND2x2_ASAP7_75t_SL g489 ( .A(n_464), .B(n_400), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_448), .B(n_9), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_432), .B(n_427), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_460), .A2(n_412), .B1(n_400), .B2(n_159), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_441), .B(n_159), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_444), .A2(n_412), .B(n_400), .Y(n_494) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_446), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_433), .B(n_412), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_433), .B(n_13), .Y(n_497) );
NAND2x1_ASAP7_75t_SL g498 ( .A(n_453), .B(n_399), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_438), .B(n_15), .Y(n_499) );
OAI31xp33_ASAP7_75t_L g500 ( .A1(n_445), .A2(n_314), .A3(n_399), .B(n_357), .Y(n_500) );
OAI31xp33_ASAP7_75t_L g501 ( .A1(n_445), .A2(n_357), .A3(n_294), .B(n_296), .Y(n_501) );
INVx2_ASAP7_75t_SL g502 ( .A(n_446), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_438), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_444), .B(n_16), .Y(n_504) );
INVxp67_ASAP7_75t_L g505 ( .A(n_443), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_460), .A2(n_383), .B1(n_367), .B2(n_365), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_443), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_453), .Y(n_508) );
AOI211xp5_ASAP7_75t_L g509 ( .A1(n_463), .A2(n_199), .B(n_203), .C(n_208), .Y(n_509) );
OAI21xp5_ASAP7_75t_SL g510 ( .A1(n_440), .A2(n_357), .B(n_365), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_456), .B(n_16), .Y(n_511) );
OR2x6_ASAP7_75t_L g512 ( .A(n_455), .B(n_358), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_447), .B(n_17), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_455), .A2(n_358), .B(n_353), .Y(n_514) );
BUFx3_ASAP7_75t_L g515 ( .A(n_435), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_437), .A2(n_367), .B1(n_365), .B2(n_339), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_462), .B(n_53), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g518 ( .A1(n_462), .A2(n_365), .B1(n_367), .B2(n_312), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_469), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_510), .A2(n_454), .B1(n_457), .B2(n_456), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_469), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_479), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_476), .B(n_468), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_491), .B(n_457), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_491), .B(n_461), .Y(n_525) );
BUFx2_ASAP7_75t_L g526 ( .A(n_488), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_508), .Y(n_527) );
NAND2x1_ASAP7_75t_L g528 ( .A(n_488), .B(n_452), .Y(n_528) );
OR2x6_ASAP7_75t_L g529 ( .A(n_512), .B(n_461), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_505), .B(n_17), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_482), .Y(n_531) );
NAND5xp2_ASAP7_75t_L g532 ( .A(n_509), .B(n_436), .C(n_450), .D(n_21), .E(n_19), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_488), .B(n_436), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_497), .B(n_461), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_508), .Y(n_535) );
INVx3_ASAP7_75t_R g536 ( .A(n_517), .Y(n_536) );
INVx2_ASAP7_75t_SL g537 ( .A(n_472), .Y(n_537) );
OAI221xp5_ASAP7_75t_L g538 ( .A1(n_513), .A2(n_225), .B1(n_451), .B2(n_222), .C(n_217), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_507), .B(n_18), .Y(n_539) );
BUFx2_ASAP7_75t_L g540 ( .A(n_482), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_503), .B(n_434), .Y(n_541) );
NOR3xp33_ASAP7_75t_L g542 ( .A(n_470), .B(n_217), .C(n_222), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_502), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_503), .B(n_434), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_479), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_502), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_480), .Y(n_547) );
AND2x2_ASAP7_75t_SL g548 ( .A(n_489), .B(n_452), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_474), .B(n_434), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_497), .B(n_23), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_486), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_499), .Y(n_552) );
AND2x2_ASAP7_75t_SL g553 ( .A(n_489), .B(n_435), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_475), .B(n_434), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_480), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_486), .Y(n_556) );
AND2x4_ASAP7_75t_SL g557 ( .A(n_466), .B(n_452), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_495), .Y(n_558) );
AND2x4_ASAP7_75t_SL g559 ( .A(n_466), .B(n_452), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_475), .B(n_451), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_496), .B(n_451), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_473), .A2(n_451), .B1(n_343), .B2(n_312), .Y(n_562) );
NAND3xp33_ASAP7_75t_L g563 ( .A(n_490), .B(n_199), .C(n_208), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_474), .B(n_496), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_466), .B(n_24), .Y(n_565) );
OAI33xp33_ASAP7_75t_L g566 ( .A1(n_511), .A2(n_26), .A3(n_28), .B1(n_29), .B2(n_43), .B3(n_45), .Y(n_566) );
OAI21xp5_ASAP7_75t_L g567 ( .A1(n_485), .A2(n_312), .B(n_222), .Y(n_567) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_504), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_477), .B(n_47), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_499), .B(n_208), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g571 ( .A(n_492), .B(n_511), .C(n_506), .D(n_487), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_477), .B(n_51), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_478), .B(n_212), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_512), .A2(n_343), .B1(n_312), .B2(n_356), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_504), .B(n_212), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_493), .Y(n_576) );
NAND4xp25_ASAP7_75t_L g577 ( .A(n_500), .B(n_217), .C(n_266), .D(n_249), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_498), .Y(n_578) );
NAND3xp33_ASAP7_75t_L g579 ( .A(n_517), .B(n_199), .C(n_203), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_477), .B(n_54), .Y(n_580) );
INVxp67_ASAP7_75t_L g581 ( .A(n_526), .Y(n_581) );
NAND3xp33_ASAP7_75t_SL g582 ( .A(n_533), .B(n_518), .C(n_516), .Y(n_582) );
XNOR2xp5_ASAP7_75t_L g583 ( .A(n_548), .B(n_471), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_524), .B(n_515), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_552), .B(n_483), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_548), .B(n_517), .Y(n_586) );
BUFx2_ASAP7_75t_L g587 ( .A(n_540), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_523), .Y(n_588) );
NAND2x1p5_ASAP7_75t_L g589 ( .A(n_553), .B(n_483), .Y(n_589) );
NAND2xp33_ASAP7_75t_L g590 ( .A(n_533), .B(n_467), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_524), .B(n_515), .Y(n_591) );
XNOR2x2_ASAP7_75t_L g592 ( .A(n_531), .B(n_514), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_553), .B(n_494), .Y(n_593) );
NAND2xp33_ASAP7_75t_L g594 ( .A(n_578), .B(n_498), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_564), .B(n_512), .Y(n_595) );
A2O1A1Ixp33_ASAP7_75t_L g596 ( .A1(n_550), .A2(n_501), .B(n_481), .C(n_343), .Y(n_596) );
NAND2x1_ASAP7_75t_SL g597 ( .A(n_568), .B(n_481), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_537), .B(n_481), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_537), .B(n_481), .Y(n_599) );
OAI21xp5_ASAP7_75t_L g600 ( .A1(n_579), .A2(n_312), .B(n_356), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_525), .B(n_481), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_519), .Y(n_602) );
NOR4xp25_ASAP7_75t_L g603 ( .A(n_571), .B(n_484), .C(n_343), .D(n_67), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_525), .B(n_484), .Y(n_604) );
OA21x2_ASAP7_75t_L g605 ( .A1(n_520), .A2(n_484), .B(n_207), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_529), .B(n_56), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_521), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_522), .B(n_212), .Y(n_608) );
A2O1A1Ixp33_ASAP7_75t_L g609 ( .A1(n_539), .A2(n_356), .B(n_296), .C(n_353), .Y(n_609) );
NOR3xp33_ASAP7_75t_L g610 ( .A(n_566), .B(n_271), .C(n_307), .Y(n_610) );
AND2x4_ASAP7_75t_L g611 ( .A(n_529), .B(n_64), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_557), .B(n_68), .Y(n_612) );
AOI31xp33_ASAP7_75t_L g613 ( .A1(n_530), .A2(n_70), .A3(n_71), .B(n_72), .Y(n_613) );
XNOR2x1_ASAP7_75t_L g614 ( .A(n_528), .B(n_75), .Y(n_614) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_558), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_557), .B(n_76), .Y(n_616) );
NOR2x1_ASAP7_75t_L g617 ( .A(n_532), .B(n_271), .Y(n_617) );
INVx3_ASAP7_75t_SL g618 ( .A(n_570), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_545), .B(n_218), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_547), .Y(n_620) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_563), .B(n_218), .C(n_199), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_559), .B(n_78), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_527), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_555), .Y(n_624) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_558), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_559), .B(n_218), .Y(n_626) );
OR2x2_ASAP7_75t_L g627 ( .A(n_534), .B(n_203), .Y(n_627) );
INVxp67_ASAP7_75t_L g628 ( .A(n_544), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_554), .B(n_218), .Y(n_629) );
NAND3xp33_ASAP7_75t_L g630 ( .A(n_538), .B(n_203), .C(n_208), .Y(n_630) );
NAND2x1_ASAP7_75t_SL g631 ( .A(n_536), .B(n_307), .Y(n_631) );
AOI211xp5_ASAP7_75t_SL g632 ( .A1(n_594), .A2(n_536), .B(n_549), .C(n_580), .Y(n_632) );
NAND5xp2_ASAP7_75t_L g633 ( .A(n_596), .B(n_562), .C(n_567), .D(n_574), .E(n_542), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_588), .B(n_554), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_602), .Y(n_635) );
INVx1_ASAP7_75t_SL g636 ( .A(n_587), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_607), .Y(n_637) );
XOR2x2_ASAP7_75t_L g638 ( .A(n_583), .B(n_580), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_584), .B(n_560), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_620), .Y(n_640) );
INVx3_ASAP7_75t_L g641 ( .A(n_589), .Y(n_641) );
XNOR2x1_ASAP7_75t_L g642 ( .A(n_617), .B(n_569), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_628), .B(n_541), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_624), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_615), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_615), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_628), .B(n_541), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_625), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_625), .Y(n_649) );
XOR2xp5_ASAP7_75t_L g650 ( .A(n_614), .B(n_570), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_603), .A2(n_576), .B1(n_560), .B2(n_561), .C(n_546), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_591), .B(n_561), .Y(n_652) );
NOR3xp33_ASAP7_75t_SL g653 ( .A(n_582), .B(n_577), .C(n_573), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_604), .B(n_549), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_581), .B(n_544), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_581), .B(n_543), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_618), .B(n_543), .Y(n_657) );
XNOR2x2_ASAP7_75t_L g658 ( .A(n_592), .B(n_572), .Y(n_658) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_582), .B(n_572), .C(n_569), .D(n_565), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_618), .B(n_546), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_585), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_595), .B(n_565), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_601), .B(n_535), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_586), .A2(n_529), .B1(n_535), .B2(n_556), .Y(n_664) );
XNOR2xp5_ASAP7_75t_L g665 ( .A(n_586), .B(n_529), .Y(n_665) );
INVxp67_ASAP7_75t_L g666 ( .A(n_629), .Y(n_666) );
INVxp67_ASAP7_75t_L g667 ( .A(n_590), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g668 ( .A1(n_613), .A2(n_575), .B(n_551), .C(n_197), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_L g669 ( .A1(n_609), .A2(n_575), .B(n_216), .C(n_212), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_593), .A2(n_312), .B1(n_356), .B2(n_334), .Y(n_670) );
OAI21xp5_ASAP7_75t_L g671 ( .A1(n_630), .A2(n_312), .B(n_356), .Y(n_671) );
OAI322xp33_ASAP7_75t_L g672 ( .A1(n_598), .A2(n_278), .A3(n_334), .B1(n_353), .B2(n_358), .C1(n_599), .C2(n_593), .Y(n_672) );
INVx1_ASAP7_75t_SL g673 ( .A(n_612), .Y(n_673) );
INVx2_ASAP7_75t_SL g674 ( .A(n_631), .Y(n_674) );
OAI321xp33_ASAP7_75t_L g675 ( .A1(n_589), .A2(n_596), .A3(n_622), .B1(n_616), .B2(n_600), .C(n_626), .Y(n_675) );
AOI31xp33_ASAP7_75t_L g676 ( .A1(n_606), .A2(n_353), .A3(n_358), .B(n_611), .Y(n_676) );
OAI222xp33_ASAP7_75t_L g677 ( .A1(n_606), .A2(n_358), .B1(n_611), .B2(n_627), .C1(n_623), .C2(n_619), .Y(n_677) );
XNOR2xp5_ASAP7_75t_L g678 ( .A(n_605), .B(n_610), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_597), .B(n_605), .Y(n_679) );
INVx2_ASAP7_75t_SL g680 ( .A(n_608), .Y(n_680) );
INVxp67_ASAP7_75t_L g681 ( .A(n_605), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_609), .B(n_621), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g683 ( .A1(n_610), .A2(n_613), .B(n_590), .C(n_603), .Y(n_683) );
NOR2xp33_ASAP7_75t_SL g684 ( .A(n_587), .B(n_548), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_602), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_602), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_603), .B(n_587), .Y(n_687) );
NAND3xp33_ASAP7_75t_SL g688 ( .A(n_683), .B(n_668), .C(n_667), .Y(n_688) );
XNOR2xp5_ASAP7_75t_L g689 ( .A(n_638), .B(n_642), .Y(n_689) );
AOI21xp33_ASAP7_75t_L g690 ( .A1(n_683), .A2(n_687), .B(n_678), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_686), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_668), .A2(n_675), .B(n_638), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_684), .A2(n_676), .B(n_642), .Y(n_693) );
XNOR2xp5_ASAP7_75t_L g694 ( .A(n_650), .B(n_673), .Y(n_694) );
AOI22x1_ASAP7_75t_L g695 ( .A1(n_632), .A2(n_636), .B1(n_641), .B2(n_665), .Y(n_695) );
NOR2xp33_ASAP7_75t_SL g696 ( .A(n_674), .B(n_659), .Y(n_696) );
AO22x2_ASAP7_75t_L g697 ( .A1(n_661), .A2(n_641), .B1(n_646), .B2(n_645), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_641), .A2(n_664), .B1(n_660), .B2(n_657), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_639), .B(n_652), .Y(n_699) );
O2A1O1Ixp33_ASAP7_75t_L g700 ( .A1(n_653), .A2(n_681), .B(n_669), .C(n_633), .Y(n_700) );
O2A1O1Ixp33_ASAP7_75t_SL g701 ( .A1(n_677), .A2(n_651), .B(n_658), .C(n_679), .Y(n_701) );
AND2x4_ASAP7_75t_L g702 ( .A(n_693), .B(n_685), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_690), .A2(n_634), .B1(n_635), .B2(n_637), .C(n_644), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g704 ( .A1(n_692), .A2(n_653), .B1(n_655), .B2(n_640), .C(n_656), .Y(n_704) );
AOI211xp5_ASAP7_75t_SL g705 ( .A1(n_701), .A2(n_658), .B(n_682), .C(n_672), .Y(n_705) );
OAI211xp5_ASAP7_75t_SL g706 ( .A1(n_700), .A2(n_670), .B(n_669), .C(n_666), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_691), .B(n_654), .Y(n_707) );
OAI21x1_ASAP7_75t_L g708 ( .A1(n_695), .A2(n_648), .B(n_649), .Y(n_708) );
NOR2x1p5_ASAP7_75t_L g709 ( .A(n_688), .B(n_643), .Y(n_709) );
NAND3xp33_ASAP7_75t_SL g710 ( .A(n_705), .B(n_696), .C(n_671), .Y(n_710) );
OAI311xp33_ASAP7_75t_L g711 ( .A1(n_704), .A2(n_689), .A3(n_697), .B1(n_694), .C1(n_698), .Y(n_711) );
NOR3xp33_ASAP7_75t_SL g712 ( .A(n_706), .B(n_662), .C(n_697), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_702), .A2(n_654), .B1(n_699), .B2(n_647), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_707), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_710), .A2(n_702), .B1(n_709), .B2(n_703), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_711), .A2(n_708), .B(n_663), .Y(n_716) );
XNOR2xp5_ASAP7_75t_L g717 ( .A(n_712), .B(n_680), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_717), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_715), .Y(n_719) );
XOR2xp5_ASAP7_75t_L g720 ( .A(n_718), .B(n_716), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_719), .Y(n_721) );
OR3x2_ASAP7_75t_L g722 ( .A(n_721), .B(n_719), .C(n_714), .Y(n_722) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_722), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_723), .A2(n_720), .B(n_713), .Y(n_724) );
endmodule