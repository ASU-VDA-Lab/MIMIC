module fake_jpeg_19370_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_43),
.Y(n_45)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_16),
.B1(n_20),
.B2(n_33),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_47),
.A2(n_31),
.B1(n_32),
.B2(n_18),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_23),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_39),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_33),
.B1(n_19),
.B2(n_20),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_41),
.B1(n_43),
.B2(n_19),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_33),
.B1(n_20),
.B2(n_19),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_60),
.A2(n_31),
.B1(n_32),
.B2(n_18),
.Y(n_98)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_42),
.B(n_30),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_63),
.B(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_17),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

BUFx4f_ASAP7_75t_SL g66 ( 
.A(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_64),
.B(n_41),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_34),
.C(n_39),
.Y(n_117)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_73),
.Y(n_122)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_28),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_75),
.Y(n_114)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_78),
.B(n_79),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_54),
.B(n_26),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_82),
.A2(n_89),
.B1(n_97),
.B2(n_98),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_62),
.B(n_21),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_88),
.Y(n_120)
);

AO22x2_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_40),
.B1(n_35),
.B2(n_39),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_90),
.A2(n_93),
.B(n_96),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_47),
.A2(n_38),
.B1(n_29),
.B2(n_23),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_105),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_60),
.A2(n_38),
.B1(n_29),
.B2(n_35),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_15),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_29),
.B1(n_35),
.B2(n_21),
.Y(n_94)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_95),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_15),
.Y(n_96)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_99),
.Y(n_131)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_17),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_104),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_58),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_37),
.B1(n_34),
.B2(n_24),
.Y(n_133)
);

NAND2x1_ASAP7_75t_L g107 ( 
.A(n_49),
.B(n_40),
.Y(n_107)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_40),
.C(n_39),
.Y(n_109)
);

XNOR2x1_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_112),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_40),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_117),
.B(n_129),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_65),
.A2(n_44),
.B1(n_40),
.B2(n_37),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_137),
.B1(n_93),
.B2(n_96),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_67),
.B(n_15),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_0),
.B(n_1),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_37),
.C(n_34),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_95),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_82),
.A2(n_44),
.B1(n_37),
.B2(n_34),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_138),
.Y(n_139)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

AO22x1_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_89),
.B1(n_90),
.B2(n_69),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_152),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_115),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_141),
.B(n_143),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_119),
.A2(n_97),
.B1(n_85),
.B2(n_68),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_147),
.B1(n_148),
.B2(n_151),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_SL g143 ( 
.A(n_125),
.B(n_87),
.C(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_144),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_162),
.B1(n_108),
.B2(n_127),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_146),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_89),
.B1(n_98),
.B2(n_103),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_89),
.B1(n_84),
.B2(n_99),
.Y(n_148)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_156),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_117),
.A2(n_90),
.B1(n_84),
.B2(n_77),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_72),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_136),
.A2(n_86),
.B1(n_70),
.B2(n_105),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_121),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_155),
.B(n_157),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_110),
.B(n_76),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_169),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_159),
.A2(n_164),
.B1(n_109),
.B2(n_127),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_80),
.B1(n_74),
.B2(n_96),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_167),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_80),
.B1(n_74),
.B2(n_44),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_123),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_132),
.A2(n_24),
.B1(n_25),
.B2(n_22),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_168),
.A2(n_118),
.B1(n_131),
.B2(n_114),
.Y(n_185)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_166),
.A2(n_111),
.B(n_135),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_170),
.A2(n_184),
.B(n_192),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_112),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_187),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_178),
.A2(n_182),
.B1(n_149),
.B2(n_12),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_129),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_183),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_155),
.A2(n_134),
.B1(n_130),
.B2(n_120),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_153),
.B(n_135),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_165),
.A2(n_118),
.B(n_134),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_185),
.A2(n_189),
.B1(n_199),
.B2(n_201),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_118),
.Y(n_187)
);

AOI32xp33_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_120),
.A3(n_122),
.B1(n_131),
.B2(n_114),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_142),
.A2(n_116),
.B1(n_113),
.B2(n_126),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_139),
.B(n_116),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_151),
.B(n_10),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_159),
.C(n_168),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_66),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_196),
.B(n_157),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_66),
.B(n_83),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_197),
.A2(n_200),
.B(n_170),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_145),
.A2(n_24),
.B1(n_104),
.B2(n_25),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_147),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_199)
);

XOR2x2_ASAP7_75t_L g200 ( 
.A(n_140),
.B(n_24),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_148),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_203),
.B(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_204),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_191),
.B(n_158),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_175),
.B(n_182),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_209),
.B(n_228),
.Y(n_252)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

A2O1A1O1Ixp25_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_172),
.B(n_183),
.C(n_179),
.D(n_195),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_231),
.Y(n_253)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_172),
.A2(n_144),
.B(n_140),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_217),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_222),
.Y(n_243)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_181),
.A2(n_167),
.B1(n_169),
.B2(n_141),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_218),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_164),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_220),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_192),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_226),
.B1(n_201),
.B2(n_199),
.Y(n_235)
);

OAI32xp33_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_149),
.A3(n_25),
.B1(n_22),
.B2(n_161),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_225),
.Y(n_239)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_227),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_186),
.B(n_161),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_186),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_229),
.Y(n_237)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_230),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_226),
.A2(n_177),
.B1(n_220),
.B2(n_214),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_233),
.A2(n_244),
.B1(n_245),
.B2(n_222),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_176),
.C(n_178),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_216),
.C(n_224),
.Y(n_254)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_227),
.A2(n_177),
.B1(n_208),
.B2(n_219),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_211),
.A2(n_185),
.B1(n_202),
.B2(n_180),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_223),
.A2(n_202),
.B1(n_173),
.B2(n_184),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_246),
.A2(n_247),
.B1(n_206),
.B2(n_218),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_223),
.A2(n_173),
.B1(n_1),
.B2(n_2),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_255),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_253),
.B(n_212),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_215),
.B(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_256),
.B(n_270),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_215),
.C(n_225),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_263),
.C(n_264),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_246),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_247),
.A2(n_210),
.B1(n_206),
.B2(n_221),
.Y(n_259)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_260),
.A2(n_267),
.B1(n_248),
.B2(n_240),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_205),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_272),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_205),
.C(n_213),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_217),
.C(n_25),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_236),
.Y(n_265)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_233),
.A2(n_11),
.B1(n_10),
.B2(n_2),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_22),
.C(n_11),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_251),
.C(n_245),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_242),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_251),
.B1(n_239),
.B2(n_240),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_0),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_232),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_273),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_0),
.Y(n_272)
);

INVxp67_ASAP7_75t_SL g273 ( 
.A(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_244),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_3),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_281),
.A2(n_269),
.B1(n_255),
.B2(n_2),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_237),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_284),
.B(n_285),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_260),
.B1(n_241),
.B2(n_272),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_262),
.A2(n_248),
.B1(n_249),
.B2(n_239),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_287),
.B(n_267),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_241),
.C(n_249),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_264),
.C(n_268),
.Y(n_294)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_261),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_293),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_299),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_296),
.B1(n_301),
.B2(n_278),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_281),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_285),
.C(n_289),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_280),
.C(n_277),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_275),
.A2(n_3),
.B(n_4),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_295),
.C(n_282),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_286),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_294),
.Y(n_303)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_309),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_307),
.B(n_310),
.Y(n_311)
);

AOI21x1_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_274),
.B(n_283),
.Y(n_308)
);

OA21x2_ASAP7_75t_L g315 ( 
.A1(n_308),
.A2(n_300),
.B(n_299),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_288),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_301),
.B1(n_296),
.B2(n_282),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_293),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_304),
.B(n_297),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_314),
.B(n_315),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_317),
.A2(n_318),
.B(n_302),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_310),
.C(n_277),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_313),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_320),
.A2(n_303),
.B(n_316),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_322),
.B(n_319),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_315),
.B(n_291),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_4),
.C(n_5),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_4),
.C(n_6),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_7),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_7),
.Y(n_328)
);


endmodule