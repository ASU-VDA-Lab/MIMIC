module real_jpeg_28749_n_17 (n_8, n_0, n_2, n_10, n_9, n_330, n_12, n_6, n_11, n_14, n_7, n_329, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_330;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_329;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_0),
.A2(n_33),
.B1(n_35),
.B2(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_44),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_0),
.A2(n_44),
.B1(n_99),
.B2(n_100),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_0),
.A2(n_44),
.B1(n_157),
.B2(n_158),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_35),
.Y(n_34)
);

A2O1A1O1Ixp25_ASAP7_75t_L g37 ( 
.A1(n_1),
.A2(n_34),
.B(n_35),
.C(n_38),
.D(n_42),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_1),
.B(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_1),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_1),
.A2(n_60),
.B(n_64),
.Y(n_86)
);

A2O1A1O1Ixp25_ASAP7_75t_L g98 ( 
.A1(n_1),
.A2(n_99),
.B(n_101),
.C(n_102),
.D(n_104),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_1),
.B(n_99),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_1),
.B(n_130),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_SL g155 ( 
.A1(n_1),
.A2(n_132),
.B(n_156),
.C(n_157),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_1),
.A2(n_81),
.B1(n_157),
.B2(n_158),
.Y(n_165)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_3),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_3),
.A2(n_33),
.B1(n_35),
.B2(n_154),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_3),
.A2(n_99),
.B1(n_100),
.B2(n_154),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_3),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_299)
);

BUFx12_ASAP7_75t_L g132 ( 
.A(n_4),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_217),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_5),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_5),
.A2(n_33),
.B1(n_35),
.B2(n_217),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_5),
.A2(n_99),
.B1(n_100),
.B2(n_217),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_7),
.A2(n_33),
.B1(n_35),
.B2(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_56),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_7),
.A2(n_56),
.B1(n_99),
.B2(n_100),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_7),
.A2(n_56),
.B1(n_157),
.B2(n_158),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_8),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_8),
.A2(n_33),
.B1(n_35),
.B2(n_114),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_8),
.A2(n_99),
.B1(n_100),
.B2(n_114),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_8),
.A2(n_114),
.B1(n_157),
.B2(n_158),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g158 ( 
.A(n_9),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_63),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_10),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_10),
.A2(n_33),
.B1(n_35),
.B2(n_63),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_10),
.A2(n_63),
.B1(n_99),
.B2(n_100),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_10),
.A2(n_63),
.B1(n_157),
.B2(n_158),
.Y(n_210)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_11),
.B(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_11),
.B(n_35),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_12),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_12),
.A2(n_33),
.B1(n_35),
.B2(n_199),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_12),
.A2(n_99),
.B1(n_100),
.B2(n_199),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_12),
.A2(n_157),
.B1(n_158),
.B2(n_199),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_13),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_13),
.A2(n_33),
.B1(n_35),
.B2(n_136),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_13),
.A2(n_99),
.B1(n_100),
.B2(n_136),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_13),
.A2(n_136),
.B1(n_157),
.B2(n_158),
.Y(n_289)
);

BUFx24_ASAP7_75t_L g100 ( 
.A(n_14),
.Y(n_100)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_15),
.A2(n_51),
.B1(n_99),
.B2(n_100),
.Y(n_103)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_16),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_313),
.Y(n_17)
);

OAI321xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_277),
.A3(n_306),
.B1(n_311),
.B2(n_312),
.C(n_329),
.Y(n_18)
);

AOI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_227),
.A3(n_266),
.B1(n_271),
.B2(n_276),
.C(n_330),
.Y(n_19)
);

NOR3xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_178),
.C(n_223),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_145),
.B(n_177),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_119),
.B(n_144),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_94),
.B(n_118),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_68),
.B(n_93),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_46),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_26),
.B(n_46),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_37),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_27),
.B(n_37),
.Y(n_77)
);

AOI32xp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.A3(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_28),
.B(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_29),
.B(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_35),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g117 ( 
.A(n_33),
.B(n_52),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_39),
.B(n_40),
.C(n_41),
.Y(n_38)
);

AOI32xp33_ASAP7_75t_L g115 ( 
.A1(n_35),
.A2(n_100),
.A3(n_101),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_38),
.A2(n_41),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_38),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_38),
.A2(n_41),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_38),
.A2(n_41),
.B1(n_243),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_42),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_55),
.B(n_57),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_45),
.A2(n_57),
.B(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_45),
.A2(n_141),
.B1(n_176),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_45),
.A2(n_141),
.B1(n_201),
.B2(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_45),
.A2(n_141),
.B(n_252),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_59),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_54),
.C(n_59),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_50),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_50),
.A2(n_102),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_50),
.A2(n_102),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_50),
.A2(n_102),
.B1(n_255),
.B2(n_284),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_50),
.A2(n_102),
.B(n_319),
.Y(n_318)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_55),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B(n_64),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_66),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_60),
.A2(n_113),
.B1(n_135),
.B2(n_137),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_60),
.A2(n_76),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_60),
.A2(n_76),
.B1(n_198),
.B2(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_60),
.A2(n_76),
.B(n_216),
.Y(n_245)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_72),
.B(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_67),
.A2(n_84),
.B(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_SL g137 ( 
.A(n_67),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_67),
.A2(n_73),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_78),
.B(n_92),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_77),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_77),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_85),
.B(n_91),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_80),
.B(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_89),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_81),
.A2(n_99),
.B(n_131),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_95),
.B(n_96),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_110),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_107),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_107),
.C(n_110),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_99),
.A2(n_100),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_102),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_104),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_106),
.A2(n_125),
.B(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_106),
.A2(n_186),
.B1(n_213),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_106),
.A2(n_186),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_109),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_115),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_121),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_138),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_139),
.C(n_140),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_128),
.C(n_134),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_124),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_134),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_130),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_130),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_130),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_130),
.A2(n_163),
.B1(n_191),
.B2(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_130),
.A2(n_163),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_132),
.B1(n_157),
.B2(n_158),
.Y(n_164)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_135),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B(n_143),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_146),
.B(n_147),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_161),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_149),
.B(n_150),
.C(n_161),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_155),
.B1(n_159),
.B2(n_160),
.Y(n_150)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_153),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_155),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_159),
.Y(n_182)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_169),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_171),
.C(n_174),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_165),
.B(n_166),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_163),
.B(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_163),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_167),
.A2(n_234),
.B(n_235),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_174),
.B2(n_175),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_173),
.Y(n_187)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_179),
.A2(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_203),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_180),
.B(n_203),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_195),
.C(n_202),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_184),
.C(n_194),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_189),
.B2(n_194),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B(n_188),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_189),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_192),
.B(n_193),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_192),
.A2(n_193),
.B(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_192),
.A2(n_234),
.B1(n_262),
.B2(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_192),
.A2(n_234),
.B1(n_289),
.B2(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_202),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_200),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_203)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_214),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_205),
.B(n_214),
.C(n_222),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_209),
.C(n_211),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_210),
.Y(n_235)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_218),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_224),
.B(n_225),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_247),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_228),
.B(n_247),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_239),
.C(n_246),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_229),
.B(n_239),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_238),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_230),
.Y(n_238)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_236),
.C(n_238),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_237),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_244),
.B2(n_245),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_245),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_245),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_245),
.A2(n_260),
.B(n_263),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_265),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_257),
.B1(n_258),
.B2(n_264),
.Y(n_248)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_253),
.B(n_256),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_253),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_256),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_256),
.A2(n_279),
.B1(n_280),
.B2(n_291),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_264),
.C(n_265),
.Y(n_307)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_263),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_267),
.A2(n_272),
.B(n_275),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_268),
.B(n_269),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_294),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_294),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_291),
.C(n_292),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_288),
.B2(n_290),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_283),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_287),
.C(n_288),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_284),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_285),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_287),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_287),
.B(n_298),
.C(n_302),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_288),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_290),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_297),
.C(n_305),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_292),
.A2(n_293),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_305),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_299),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_304),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_327),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_326),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_316),
.B(n_326),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_325),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_320),
.B1(n_323),
.B2(n_324),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_318),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_320),
.Y(n_323)
);


endmodule