module fake_jpeg_7878_n_267 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_267);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_267;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_218;
wire n_63;
wire n_92;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_41),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_17),
.B1(n_22),
.B2(n_33),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_45),
.A2(n_47),
.B1(n_49),
.B2(n_58),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_28),
.B1(n_26),
.B2(n_23),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_46),
.A2(n_55),
.B(n_60),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_17),
.B1(n_22),
.B2(n_33),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_18),
.B1(n_31),
.B2(n_21),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_28),
.B1(n_16),
.B2(n_26),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_20),
.B1(n_23),
.B2(n_27),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_61),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_20),
.B1(n_27),
.B2(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_31),
.B1(n_27),
.B2(n_25),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_43),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_31),
.B1(n_25),
.B2(n_21),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_21),
.B1(n_30),
.B2(n_19),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_38),
.B(n_42),
.C(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_67),
.B(n_74),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_68),
.B(n_70),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_42),
.B1(n_43),
.B2(n_38),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_69),
.A2(n_52),
.B1(n_57),
.B2(n_54),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_38),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_78),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_85),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_38),
.Y(n_80)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_15),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_48),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_44),
.A2(n_30),
.B1(n_32),
.B2(n_19),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_30),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_56),
.Y(n_90)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_65),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_90),
.B(n_108),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_2),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_104),
.B(n_67),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_100),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_95),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_79),
.Y(n_138)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_40),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_52),
.B1(n_57),
.B2(n_66),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_107),
.A2(n_109),
.B1(n_76),
.B2(n_72),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_68),
.B(n_54),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_57),
.B1(n_51),
.B2(n_49),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_110),
.Y(n_129)
);

BUFx12_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

MAJx2_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_40),
.C(n_35),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_71),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_115),
.Y(n_150)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_117),
.Y(n_160)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_118),
.B(n_124),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_87),
.B(n_80),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_120),
.A2(n_126),
.B(n_136),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_111),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_134),
.B1(n_135),
.B2(n_96),
.Y(n_144)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_95),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_130),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_91),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_98),
.Y(n_131)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_101),
.A2(n_87),
.B1(n_71),
.B2(n_75),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_101),
.A2(n_85),
.B1(n_88),
.B2(n_86),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_84),
.B(n_73),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_138),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_112),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_153),
.Y(n_173)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_145),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_132),
.A2(n_96),
.B1(n_93),
.B2(n_97),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_148),
.B1(n_135),
.B2(n_129),
.Y(n_168)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_146),
.B1(n_137),
.B2(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_119),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_93),
.B1(n_113),
.B2(n_82),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_99),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_151),
.B(n_159),
.Y(n_167)
);

NAND2xp33_ASAP7_75t_SL g151 ( 
.A(n_134),
.B(n_111),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_99),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_118),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_113),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_158),
.B(n_114),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_126),
.A2(n_35),
.B(n_40),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_161),
.B(n_163),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_32),
.B(n_19),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_164),
.B(n_129),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_119),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_133),
.A2(n_32),
.B1(n_19),
.B2(n_83),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_169),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_168),
.B(n_172),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_179),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_171),
.B(n_154),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_176),
.A2(n_140),
.B1(n_32),
.B2(n_35),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_130),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_177),
.B(n_183),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_157),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_145),
.B1(n_144),
.B2(n_161),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_155),
.B1(n_143),
.B2(n_154),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_115),
.Y(n_182)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_149),
.B(n_124),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_117),
.Y(n_185)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_128),
.Y(n_187)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_139),
.C(n_153),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_203),
.Y(n_210)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_206),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_159),
.B(n_155),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_176),
.B(n_187),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_204),
.B1(n_172),
.B2(n_168),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_202),
.B(n_207),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_185),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_171),
.B(n_15),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_186),
.B1(n_198),
.B2(n_199),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_212),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_181),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_202),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_214),
.C(n_207),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_167),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_217),
.B(n_220),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_216),
.A2(n_223),
.B1(n_191),
.B2(n_169),
.Y(n_227)
);

BUFx12_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_194),
.B(n_166),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_221),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_174),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_184),
.B1(n_170),
.B2(n_204),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_179),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_180),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_226),
.B(n_228),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_227),
.B(n_229),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_193),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_220),
.A2(n_201),
.B1(n_205),
.B2(n_196),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_232),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_92),
.B1(n_54),
.B2(n_83),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_233),
.A2(n_235),
.B1(n_209),
.B2(n_217),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_219),
.A2(n_92),
.B1(n_4),
.B2(n_5),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_224),
.B(n_214),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_240),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_217),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_2),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g250 ( 
.A(n_241),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_226),
.B(n_92),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_243),
.B(n_233),
.Y(n_245)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_242),
.A2(n_228),
.B(n_235),
.Y(n_248)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_248),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_231),
.B1(n_210),
.B2(n_5),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_244),
.A2(n_2),
.B(n_4),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_4),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_5),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_237),
.Y(n_255)
);

AOI322xp5_ASAP7_75t_L g261 ( 
.A1(n_255),
.A2(n_246),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_7),
.C2(n_12),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_251),
.A2(n_238),
.B(n_6),
.Y(n_257)
);

NOR3xp33_ASAP7_75t_SL g259 ( 
.A(n_257),
.B(n_250),
.C(n_245),
.Y(n_259)
);

O2A1O1Ixp33_ASAP7_75t_SL g263 ( 
.A1(n_259),
.A2(n_260),
.B(n_262),
.C(n_256),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_254),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_7),
.C2(n_13),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_7),
.C(n_8),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_264),
.C(n_12),
.Y(n_265)
);

AO21x2_ASAP7_75t_L g266 ( 
.A1(n_265),
.A2(n_12),
.B(n_14),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_14),
.Y(n_267)
);


endmodule