module real_aes_8844_n_254 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_254);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_254;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_626;
wire n_400;
wire n_539;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_812;
wire n_817;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_449;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_283;
wire n_314;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_259;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_797;
wire n_668;
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_0), .A2(n_75), .B1(n_338), .B2(n_383), .Y(n_460) );
AOI22xp33_ASAP7_75t_SL g574 ( .A1(n_1), .A2(n_162), .B1(n_575), .B2(n_577), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_2), .A2(n_52), .B1(n_345), .B2(n_537), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_3), .A2(n_238), .B1(n_557), .B2(n_558), .Y(n_556) );
AOI22xp33_ASAP7_75t_SL g432 ( .A1(n_4), .A2(n_187), .B1(n_433), .B2(n_434), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g805 ( .A1(n_5), .A2(n_44), .B1(n_541), .B2(n_612), .C(n_806), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_6), .Y(n_619) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_7), .A2(n_248), .B1(n_636), .B2(n_637), .Y(n_635) );
AOI22xp33_ASAP7_75t_SL g458 ( .A1(n_8), .A2(n_104), .B1(n_388), .B2(n_459), .Y(n_458) );
AOI222xp33_ASAP7_75t_L g706 ( .A1(n_9), .A2(n_35), .B1(n_117), .B2(n_627), .C1(n_665), .C2(n_707), .Y(n_706) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_10), .A2(n_40), .B1(n_388), .B2(n_731), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_11), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_12), .A2(n_125), .B1(n_378), .B2(n_546), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_13), .A2(n_194), .B1(n_607), .B2(n_609), .Y(n_606) );
AOI221xp5_ASAP7_75t_L g815 ( .A1(n_14), .A2(n_200), .B1(n_700), .B2(n_722), .C(n_816), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_15), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_16), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_17), .A2(n_43), .B1(n_436), .B2(n_537), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g299 ( .A(n_18), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_19), .A2(n_211), .B1(n_338), .B2(n_347), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_20), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_21), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_22), .A2(n_127), .B1(n_447), .B2(n_448), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_23), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_24), .A2(n_207), .B1(n_682), .B2(n_684), .C(n_685), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_25), .Y(n_493) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_26), .A2(n_50), .B1(n_699), .B2(n_700), .C(n_701), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_27), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_28), .A2(n_191), .B1(n_323), .B2(n_328), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_29), .B(n_793), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_30), .A2(n_252), .B1(n_455), .B2(n_530), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_31), .Y(n_473) );
AO22x2_ASAP7_75t_L g277 ( .A1(n_32), .A2(n_92), .B1(n_278), .B2(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g765 ( .A(n_32), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_33), .A2(n_79), .B1(n_378), .B2(n_380), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_34), .A2(n_57), .B1(n_378), .B2(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_36), .A2(n_220), .B1(n_345), .B2(n_537), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_37), .Y(n_750) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_38), .A2(n_77), .B1(n_612), .B2(n_692), .C(n_695), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_39), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_41), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_42), .A2(n_145), .B1(n_498), .B2(n_499), .Y(n_497) );
AOI22xp33_ASAP7_75t_SL g462 ( .A1(n_45), .A2(n_54), .B1(n_332), .B2(n_463), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_46), .Y(n_355) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_47), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g725 ( .A1(n_48), .A2(n_178), .B1(n_502), .B2(n_726), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_49), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_51), .A2(n_154), .B1(n_346), .B2(n_465), .Y(n_464) );
AO22x2_ASAP7_75t_L g281 ( .A1(n_53), .A2(n_95), .B1(n_278), .B2(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g766 ( .A(n_53), .Y(n_766) );
AOI22xp33_ASAP7_75t_SL g728 ( .A1(n_55), .A2(n_105), .B1(n_345), .B2(n_506), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_56), .A2(n_222), .B1(n_505), .B2(n_506), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_58), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_59), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_60), .B(n_744), .Y(n_743) );
AOI222xp33_ASAP7_75t_L g578 ( .A1(n_61), .A2(n_141), .B1(n_150), .B2(n_329), .C1(n_364), .C2(n_579), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_62), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_63), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_64), .A2(n_89), .B1(n_295), .B2(n_323), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_65), .A2(n_97), .B1(n_429), .B2(n_430), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_66), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_67), .A2(n_166), .B1(n_454), .B2(n_455), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g622 ( .A(n_68), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_69), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_70), .A2(n_88), .B1(n_410), .B2(n_595), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_71), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_72), .Y(n_786) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_73), .A2(n_121), .B1(n_386), .B2(n_387), .Y(n_437) );
AOI222xp33_ASAP7_75t_L g819 ( .A1(n_74), .A2(n_100), .B1(n_147), .B2(n_665), .C1(n_820), .C2(n_822), .Y(n_819) );
XNOR2x2_ASAP7_75t_L g553 ( .A(n_76), .B(n_554), .Y(n_553) );
AOI221xp5_ASAP7_75t_L g809 ( .A1(n_78), .A2(n_126), .B1(n_684), .B2(n_810), .C(n_811), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_80), .Y(n_542) );
AOI222xp33_ASAP7_75t_L g749 ( .A1(n_81), .A2(n_151), .B1(n_159), .B2(n_577), .C1(n_665), .C2(n_707), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_82), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_83), .Y(n_817) );
AOI22xp33_ASAP7_75t_SL g409 ( .A1(n_84), .A2(n_205), .B1(n_364), .B2(n_410), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_85), .A2(n_86), .B1(n_323), .B2(n_380), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g415 ( .A1(n_87), .A2(n_135), .B1(n_416), .B2(n_419), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_90), .A2(n_144), .B1(n_346), .B2(n_382), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_91), .A2(n_176), .B1(n_338), .B2(n_633), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_93), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_94), .A2(n_142), .B1(n_652), .B2(n_655), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_96), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_98), .A2(n_680), .B1(n_708), .B2(n_709), .Y(n_679) );
INVx1_ASAP7_75t_L g708 ( .A(n_98), .Y(n_708) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_99), .A2(n_235), .B1(n_305), .B2(n_454), .Y(n_723) );
AND2x2_ASAP7_75t_L g261 ( .A(n_101), .B(n_262), .Y(n_261) );
AOI211xp5_ASAP7_75t_L g254 ( .A1(n_102), .A2(n_255), .B(n_263), .C(n_767), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_103), .A2(n_230), .B1(n_390), .B2(n_502), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_106), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_107), .Y(n_734) );
INVx1_ASAP7_75t_L g258 ( .A(n_108), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_109), .A2(n_219), .B1(n_566), .B2(n_567), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_110), .A2(n_167), .B1(n_323), .B2(n_546), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_111), .A2(n_129), .B1(n_301), .B2(n_305), .Y(n_300) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_112), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_113), .A2(n_247), .B1(n_301), .B2(n_448), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_114), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_115), .B(n_367), .Y(n_366) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_116), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_118), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_119), .A2(n_123), .B1(n_726), .B2(n_739), .Y(n_738) );
OA22x2_ASAP7_75t_L g267 ( .A1(n_120), .A2(n_268), .B1(n_269), .B2(n_350), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_120), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g666 ( .A(n_122), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_124), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_128), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_130), .A2(n_231), .B1(n_429), .B2(n_569), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_131), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_132), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_133), .B(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_134), .B(n_416), .Y(n_450) );
INVx2_ASAP7_75t_L g262 ( .A(n_136), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_137), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_138), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g365 ( .A(n_139), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_140), .A2(n_146), .B1(n_560), .B2(n_563), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_143), .Y(n_672) );
AND2x6_ASAP7_75t_L g257 ( .A(n_148), .B(n_258), .Y(n_257) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_148), .Y(n_759) );
AO22x2_ASAP7_75t_L g287 ( .A1(n_149), .A2(n_204), .B1(n_278), .B2(n_282), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_152), .A2(n_175), .B1(n_380), .B2(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_153), .A2(n_182), .B1(n_386), .B2(n_387), .Y(n_385) );
AOI22xp33_ASAP7_75t_SL g423 ( .A1(n_155), .A2(n_209), .B1(n_347), .B2(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_156), .B(n_452), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_157), .A2(n_228), .B1(n_338), .B2(n_341), .Y(n_337) );
AOI22xp33_ASAP7_75t_SL g427 ( .A1(n_158), .A2(n_241), .B1(n_428), .B2(n_430), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_160), .A2(n_769), .B1(n_798), .B2(n_799), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_160), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_161), .A2(n_189), .B1(n_331), .B2(n_333), .Y(n_330) );
INVx1_ASAP7_75t_L g614 ( .A(n_163), .Y(n_614) );
AOI22xp33_ASAP7_75t_SL g412 ( .A1(n_164), .A2(n_208), .B1(n_413), .B2(n_414), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_165), .A2(n_217), .B1(n_390), .B2(n_391), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_168), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_169), .B(n_477), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_170), .A2(n_186), .B1(n_332), .B2(n_535), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_171), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_172), .A2(n_199), .B1(n_569), .B2(n_774), .Y(n_773) );
AO22x2_ASAP7_75t_L g285 ( .A1(n_173), .A2(n_221), .B1(n_278), .B2(n_279), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_174), .Y(n_597) );
AO22x1_ASAP7_75t_L g803 ( .A1(n_177), .A2(n_804), .B1(n_823), .B2(n_824), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_177), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_179), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_180), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_181), .Y(n_689) );
AOI22xp33_ASAP7_75t_SL g732 ( .A1(n_183), .A2(n_216), .B1(n_541), .B2(n_733), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_184), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_185), .A2(n_202), .B1(n_447), .B2(n_448), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_188), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_190), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_192), .Y(n_521) );
INVx1_ASAP7_75t_L g571 ( .A(n_193), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_195), .A2(n_227), .B1(n_499), .B2(n_541), .Y(n_605) );
AOI22xp33_ASAP7_75t_SL g717 ( .A1(n_196), .A2(n_232), .B1(n_410), .B2(n_448), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_197), .B(n_722), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_198), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_201), .B(n_579), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_203), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_204), .B(n_764), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g671 ( .A(n_206), .Y(n_671) );
OA22x2_ASAP7_75t_L g402 ( .A1(n_210), .A2(n_403), .B1(n_404), .B2(n_438), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_210), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_212), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_213), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_214), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g639 ( .A(n_215), .Y(n_639) );
CKINVDCx20_ASAP7_75t_R g686 ( .A(n_218), .Y(n_686) );
INVx1_ASAP7_75t_L g762 ( .A(n_221), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_223), .A2(n_239), .B1(n_323), .B2(n_331), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_224), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_225), .A2(n_229), .B1(n_345), .B2(n_347), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_226), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_233), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_234), .A2(n_641), .B1(n_673), .B2(n_674), .Y(n_640) );
INVx1_ASAP7_75t_L g673 ( .A(n_234), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_236), .Y(n_362) );
INVx1_ASAP7_75t_L g278 ( .A(n_237), .Y(n_278) );
INVx1_ASAP7_75t_L g280 ( .A(n_237), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_240), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_242), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_243), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_244), .Y(n_591) );
OA22x2_ASAP7_75t_L g514 ( .A1(n_245), .A2(n_515), .B1(n_516), .B2(n_517), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_245), .Y(n_515) );
AOI22x1_ASAP7_75t_L g351 ( .A1(n_246), .A2(n_352), .B1(n_393), .B2(n_394), .Y(n_351) );
INVx1_ASAP7_75t_L g393 ( .A(n_246), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_249), .A2(n_253), .B1(n_382), .B2(n_648), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_250), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_251), .Y(n_625) );
INVx1_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_258), .Y(n_758) );
OAI21xp5_ASAP7_75t_L g829 ( .A1(n_259), .A2(n_757), .B(n_830), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_260), .Y(n_259) );
INVxp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_677), .B1(n_752), .B2(n_753), .C(n_754), .Y(n_263) );
INVx1_ASAP7_75t_L g752 ( .A(n_264), .Y(n_752) );
XNOR2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_397), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_351), .B1(n_395), .B2(n_396), .Y(n_265) );
INVx1_ASAP7_75t_L g395 ( .A(n_266), .Y(n_395) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g350 ( .A(n_269), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_320), .Y(n_269) );
NOR3xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_293), .C(n_309), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_273), .B1(n_288), .B2(n_289), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_273), .A2(n_359), .B1(n_619), .B2(n_620), .Y(n_618) );
BUFx3_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g357 ( .A(n_274), .Y(n_357) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_274), .Y(n_484) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_283), .Y(n_274) );
INVx2_ASAP7_75t_L g296 ( .A(n_275), .Y(n_296) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_281), .Y(n_275) );
AND2x2_ASAP7_75t_L g292 ( .A(n_276), .B(n_281), .Y(n_292) );
AND2x2_ASAP7_75t_L g326 ( .A(n_276), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g304 ( .A(n_277), .B(n_287), .Y(n_304) );
AND2x2_ASAP7_75t_L g316 ( .A(n_277), .B(n_281), .Y(n_316) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g282 ( .A(n_280), .Y(n_282) );
INVx1_ASAP7_75t_L g308 ( .A(n_281), .Y(n_308) );
INVx2_ASAP7_75t_L g327 ( .A(n_281), .Y(n_327) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2x1p5_ASAP7_75t_L g291 ( .A(n_284), .B(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g346 ( .A(n_284), .B(n_326), .Y(n_346) );
AND2x4_ASAP7_75t_L g418 ( .A(n_284), .B(n_296), .Y(n_418) );
AND2x6_ASAP7_75t_L g421 ( .A(n_284), .B(n_292), .Y(n_421) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g298 ( .A(n_285), .Y(n_298) );
INVx1_ASAP7_75t_L g303 ( .A(n_285), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_285), .B(n_287), .Y(n_312) );
INVx1_ASAP7_75t_L g319 ( .A(n_285), .Y(n_319) );
AND2x2_ASAP7_75t_L g297 ( .A(n_286), .B(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g325 ( .A(n_287), .B(n_319), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_289), .A2(n_484), .B1(n_661), .B2(n_662), .Y(n_660) );
OA211x2_ASAP7_75t_L g741 ( .A1(n_289), .A2(n_742), .B(n_743), .C(n_745), .Y(n_741) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g359 ( .A(n_290), .Y(n_359) );
INVx2_ASAP7_75t_L g797 ( .A(n_290), .Y(n_797) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx3_ASAP7_75t_L g488 ( .A(n_291), .Y(n_488) );
AND2x4_ASAP7_75t_L g332 ( .A(n_292), .B(n_297), .Y(n_332) );
AND2x2_ASAP7_75t_L g343 ( .A(n_292), .B(n_325), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_292), .B(n_325), .Y(n_688) );
OAI21xp33_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_299), .B(n_300), .Y(n_293) );
INVx2_ASAP7_75t_SL g380 ( .A(n_294), .Y(n_380) );
INVx4_ASAP7_75t_L g731 ( .A(n_294), .Y(n_731) );
INVx3_ASAP7_75t_L g810 ( .A(n_294), .Y(n_810) );
INVx11_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx11_ASAP7_75t_L g426 ( .A(n_295), .Y(n_426) );
AND2x6_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x6_ASAP7_75t_L g329 ( .A(n_297), .B(n_316), .Y(n_329) );
AND2x2_ASAP7_75t_L g340 ( .A(n_297), .B(n_326), .Y(n_340) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_301), .Y(n_367) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_301), .Y(n_410) );
BUFx12f_ASAP7_75t_L g447 ( .A(n_301), .Y(n_447) );
AND2x4_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g335 ( .A(n_303), .B(n_327), .Y(n_335) );
AND2x4_ASAP7_75t_L g306 ( .A(n_304), .B(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g334 ( .A(n_304), .B(n_335), .Y(n_334) );
NAND2x1p5_ASAP7_75t_L g371 ( .A(n_304), .B(n_372), .Y(n_371) );
BUFx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_L g413 ( .A(n_306), .Y(n_413) );
BUFx3_ASAP7_75t_L g455 ( .A(n_306), .Y(n_455) );
INVx1_ASAP7_75t_L g576 ( .A(n_306), .Y(n_576) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x6_ASAP7_75t_L g311 ( .A(n_308), .B(n_312), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B1(n_313), .B2(n_314), .Y(n_309) );
INVx6_ASAP7_75t_SL g392 ( .A(n_311), .Y(n_392) );
INVx1_ASAP7_75t_SL g465 ( .A(n_311), .Y(n_465) );
INVx1_ASAP7_75t_L g609 ( .A(n_311), .Y(n_609) );
INVx1_ASAP7_75t_L g349 ( .A(n_312), .Y(n_349) );
BUFx2_ASAP7_75t_L g374 ( .A(n_314), .Y(n_374) );
CKINVDCx16_ASAP7_75t_R g602 ( .A(n_314), .Y(n_602) );
OR2x6_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g414 ( .A(n_316), .B(n_318), .Y(n_414) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_321), .B(n_336), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_330), .Y(n_321) );
BUFx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx3_ASAP7_75t_L g388 ( .A(n_324), .Y(n_388) );
BUFx3_ASAP7_75t_L g567 ( .A(n_324), .Y(n_567) );
BUFx3_ASAP7_75t_L g657 ( .A(n_324), .Y(n_657) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_325), .B(n_326), .Y(n_551) );
AND2x4_ASAP7_75t_L g348 ( .A(n_326), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g372 ( .A(n_327), .Y(n_372) );
INVx2_ASAP7_75t_SL g361 ( .A(n_328), .Y(n_361) );
INVx2_ASAP7_75t_L g472 ( .A(n_328), .Y(n_472) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g407 ( .A(n_329), .Y(n_407) );
BUFx3_ASAP7_75t_L g525 ( .A(n_329), .Y(n_525) );
INVx4_ASAP7_75t_L g593 ( .A(n_329), .Y(n_593) );
INVx2_ASAP7_75t_L g715 ( .A(n_329), .Y(n_715) );
BUFx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx3_ASAP7_75t_L g386 ( .A(n_332), .Y(n_386) );
INVx6_ASAP7_75t_L g503 ( .A(n_332), .Y(n_503) );
BUFx3_ASAP7_75t_L g654 ( .A(n_332), .Y(n_654) );
BUFx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx4f_ASAP7_75t_SL g364 ( .A(n_334), .Y(n_364) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_334), .Y(n_454) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_334), .Y(n_492) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_334), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_344), .Y(n_336) );
INVx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx3_ASAP7_75t_L g498 ( .A(n_339), .Y(n_498) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_340), .Y(n_379) );
BUFx2_ASAP7_75t_SL g541 ( .A(n_340), .Y(n_541) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_341), .Y(n_390) );
INVx5_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g429 ( .A(n_342), .Y(n_429) );
INVx4_ASAP7_75t_L g463 ( .A(n_342), .Y(n_463) );
INVx1_ASAP7_75t_L g535 ( .A(n_342), .Y(n_535) );
INVx3_ASAP7_75t_L g637 ( .A(n_342), .Y(n_637) );
BUFx3_ASAP7_75t_L g727 ( .A(n_342), .Y(n_727) );
INVx8_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g436 ( .A(n_346), .Y(n_436) );
BUFx3_ASAP7_75t_L g505 ( .A(n_346), .Y(n_505) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_346), .Y(n_562) );
INVx2_ASAP7_75t_L g649 ( .A(n_346), .Y(n_649) );
INVxp67_ASAP7_75t_L g783 ( .A(n_347), .Y(n_783) );
BUFx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx3_ASAP7_75t_L g383 ( .A(n_348), .Y(n_383) );
BUFx2_ASAP7_75t_SL g499 ( .A(n_348), .Y(n_499) );
BUFx3_ASAP7_75t_L g563 ( .A(n_348), .Y(n_563) );
BUFx2_ASAP7_75t_L g633 ( .A(n_348), .Y(n_633) );
BUFx3_ASAP7_75t_L g684 ( .A(n_348), .Y(n_684) );
BUFx2_ASAP7_75t_SL g733 ( .A(n_348), .Y(n_733) );
INVx2_ASAP7_75t_L g396 ( .A(n_351), .Y(n_396) );
INVx2_ASAP7_75t_SL g394 ( .A(n_352), .Y(n_394) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_375), .Y(n_352) );
NOR3xp33_ASAP7_75t_L g353 ( .A(n_354), .B(n_360), .C(n_368), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_358), .B2(n_359), .Y(n_354) );
OAI22xp5_ASAP7_75t_SL g519 ( .A1(n_356), .A2(n_486), .B1(n_520), .B2(n_521), .Y(n_519) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g588 ( .A(n_357), .Y(n_588) );
OA211x2_ASAP7_75t_L g570 ( .A1(n_359), .A2(n_571), .B(n_572), .C(n_574), .Y(n_570) );
OAI221xp5_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_362), .B1(n_363), .B2(n_365), .C(n_366), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g474 ( .A(n_367), .Y(n_474) );
BUFx4f_ASAP7_75t_L g579 ( .A(n_367), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B1(n_373), .B2(n_374), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_370), .A2(n_490), .B1(n_491), .B2(n_493), .Y(n_489) );
OAI22xp33_ASAP7_75t_L g527 ( .A1(n_370), .A2(n_528), .B1(n_529), .B2(n_531), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_370), .A2(n_374), .B1(n_671), .B2(n_672), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_370), .A2(n_705), .B1(n_817), .B2(n_818), .Y(n_816) );
BUFx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx4_ASAP7_75t_L g599 ( .A(n_371), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_371), .A2(n_625), .B1(n_626), .B2(n_628), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_371), .A2(n_601), .B1(n_786), .B2(n_787), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_384), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_381), .Y(n_376) );
BUFx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx3_ASAP7_75t_L g433 ( .A(n_379), .Y(n_433) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_379), .Y(n_566) );
INVx3_ASAP7_75t_L g683 ( .A(n_379), .Y(n_683) );
BUFx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_389), .Y(n_384) );
BUFx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_391), .Y(n_814) );
BUFx4f_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
BUFx2_ASAP7_75t_L g430 ( .A(n_392), .Y(n_430) );
BUFx2_ASAP7_75t_L g506 ( .A(n_392), .Y(n_506) );
BUFx2_ASAP7_75t_L g537 ( .A(n_392), .Y(n_537) );
BUFx2_ASAP7_75t_L g569 ( .A(n_392), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B1(n_509), .B2(n_676), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_439), .B2(n_440), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g438 ( .A(n_404), .Y(n_438) );
NAND3x1_ASAP7_75t_L g404 ( .A(n_405), .B(n_422), .C(n_431), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_411), .Y(n_405) );
OAI21xp5_ASAP7_75t_SL g406 ( .A1(n_407), .A2(n_408), .B(n_409), .Y(n_406) );
OAI21xp5_ASAP7_75t_SL g444 ( .A1(n_407), .A2(n_445), .B(n_446), .Y(n_444) );
BUFx2_ASAP7_75t_L g793 ( .A(n_410), .Y(n_793) );
BUFx3_ASAP7_75t_L g822 ( .A(n_410), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_415), .Y(n_411) );
BUFx2_ASAP7_75t_SL g448 ( .A(n_414), .Y(n_448) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_414), .Y(n_479) );
BUFx2_ASAP7_75t_SL g577 ( .A(n_414), .Y(n_577) );
BUFx2_ASAP7_75t_L g699 ( .A(n_416), .Y(n_699) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx5_ASAP7_75t_L g573 ( .A(n_417), .Y(n_573) );
INVx2_ASAP7_75t_L g744 ( .A(n_417), .Y(n_744) );
INVx4_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_L g452 ( .A(n_421), .Y(n_452) );
BUFx4f_ASAP7_75t_L g700 ( .A(n_421), .Y(n_700) );
BUFx2_ASAP7_75t_L g720 ( .A(n_421), .Y(n_720) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_427), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx5_ASAP7_75t_SL g459 ( .A(n_426), .Y(n_459) );
INVx1_ASAP7_75t_L g546 ( .A(n_426), .Y(n_546) );
INVx2_ASAP7_75t_L g557 ( .A(n_426), .Y(n_557) );
INVx2_ASAP7_75t_SL g694 ( .A(n_426), .Y(n_694) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_437), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_435), .A2(n_781), .B1(n_782), .B2(n_783), .Y(n_780) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
AO22x2_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_467), .B1(n_468), .B2(n_508), .Y(n_440) );
INVx3_ASAP7_75t_L g508 ( .A(n_441), .Y(n_508) );
XOR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_466), .Y(n_441) );
NAND2x1_ASAP7_75t_SL g442 ( .A(n_443), .B(n_456), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_449), .Y(n_443) );
BUFx4f_ASAP7_75t_SL g707 ( .A(n_447), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .C(n_453), .Y(n_449) );
BUFx2_ASAP7_75t_L g595 ( .A(n_454), .Y(n_595) );
INVx2_ASAP7_75t_L g667 ( .A(n_454), .Y(n_667) );
INVx4_ASAP7_75t_L g821 ( .A(n_454), .Y(n_821) );
NOR2x1_ASAP7_75t_L g456 ( .A(n_457), .B(n_461), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
INVx1_ASAP7_75t_L g646 ( .A(n_459), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
INVx2_ASAP7_75t_L g608 ( .A(n_463), .Y(n_608) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
XOR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_507), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_494), .Y(n_469) );
NOR3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_480), .C(n_489), .Y(n_470) );
OAI221xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B1(n_474), .B2(n_475), .C(n_476), .Y(n_471) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B1(n_485), .B2(n_486), .Y(n_480) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_484), .A2(n_795), .B1(n_796), .B2(n_797), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_486), .A2(n_587), .B1(n_588), .B2(n_589), .Y(n_586) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_492), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_500), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx1_ASAP7_75t_SL g543 ( .A(n_499), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_504), .Y(n_500) );
INVx2_ASAP7_75t_L g777 ( .A(n_502), .Y(n_777) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx3_ASAP7_75t_L g558 ( .A(n_503), .Y(n_558) );
INVx2_ASAP7_75t_L g636 ( .A(n_503), .Y(n_636) );
INVx2_ASAP7_75t_L g739 ( .A(n_503), .Y(n_739) );
INVx1_ASAP7_75t_L g676 ( .A(n_509), .Y(n_676) );
XOR2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_580), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B1(n_552), .B2(n_553), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_532), .Y(n_517) );
NOR3xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_522), .C(n_527), .Y(n_518) );
OAI21xp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B(n_526), .Y(n_522) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_530), .Y(n_529) );
NOR3xp33_ASAP7_75t_L g532 ( .A(n_533), .B(n_538), .C(n_544), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_535), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B1(n_542), .B2(n_543), .Y(n_538) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_547), .B1(n_548), .B2(n_549), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_549), .A2(n_653), .B1(n_696), .B2(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g779 ( .A(n_550), .Y(n_779) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND4xp75_ASAP7_75t_L g554 ( .A(n_555), .B(n_564), .C(n_570), .D(n_578), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_559), .Y(n_555) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx4_ASAP7_75t_L g612 ( .A(n_561), .Y(n_612) );
INVx4_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_568), .Y(n_564) );
INVx1_ASAP7_75t_L g690 ( .A(n_569), .Y(n_690) );
BUFx6f_ASAP7_75t_L g722 ( .A(n_573), .Y(n_722) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .B1(n_640), .B2(n_675), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
XNOR2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_615), .Y(n_582) );
XOR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_614), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_603), .Y(n_584) );
NOR3xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_590), .C(n_596), .Y(n_585) );
OAI21xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B(n_594), .Y(n_590) );
BUFx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI21xp5_ASAP7_75t_SL g621 ( .A1(n_593), .A2(n_622), .B(n_623), .Y(n_621) );
INVx4_ASAP7_75t_L g665 ( .A(n_593), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B1(n_600), .B2(n_601), .Y(n_596) );
INVx3_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g703 ( .A(n_599), .Y(n_703) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g705 ( .A(n_602), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_610), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
XOR2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_639), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_629), .Y(n_616) );
NOR3xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_621), .C(n_624), .Y(n_617) );
INVx2_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_SL g790 ( .A(n_627), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_634), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_638), .Y(n_634) );
INVx1_ASAP7_75t_L g675 ( .A(n_640), .Y(n_675) );
INVx2_ASAP7_75t_L g674 ( .A(n_641), .Y(n_674) );
AND2x2_ASAP7_75t_SL g641 ( .A(n_642), .B(n_659), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_650), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_647), .Y(n_643) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_658), .Y(n_650) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NOR3xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_663), .C(n_670), .Y(n_659) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B1(n_667), .B2(n_668), .C(n_669), .Y(n_663) );
OAI221xp5_ASAP7_75t_L g788 ( .A1(n_664), .A2(n_789), .B1(n_790), .B2(n_791), .C(n_792), .Y(n_788) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
CKINVDCx16_ASAP7_75t_R g753 ( .A(n_677), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_710), .B2(n_751), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g709 ( .A(n_680), .Y(n_709) );
AND4x1_ASAP7_75t_L g680 ( .A(n_681), .B(n_691), .C(n_698), .D(n_706), .Y(n_680) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_689), .B2(n_690), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_687), .A2(n_812), .B1(n_813), .B2(n_814), .Y(n_811) );
BUFx2_ASAP7_75t_R g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B1(n_704), .B2(n_705), .Y(n_701) );
INVx2_ASAP7_75t_SL g751 ( .A(n_710), .Y(n_751) );
XNOR2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_735), .Y(n_710) );
XOR2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_734), .Y(n_711) );
NAND3x1_ASAP7_75t_L g712 ( .A(n_713), .B(n_724), .C(n_729), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_718), .Y(n_713) );
OAI21xp5_ASAP7_75t_SL g714 ( .A1(n_715), .A2(n_716), .B(n_717), .Y(n_714) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_721), .C(n_723), .Y(n_718) );
AND2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_728), .Y(n_724) );
INVx3_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
XOR2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_750), .Y(n_735) );
NAND4xp75_ASAP7_75t_L g736 ( .A(n_737), .B(n_741), .C(n_746), .D(n_749), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_740), .Y(n_737) );
AND2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
NOR2x1_ASAP7_75t_L g755 ( .A(n_756), .B(n_760), .Y(n_755) );
OR2x2_ASAP7_75t_SL g827 ( .A(n_756), .B(n_761), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_759), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_757), .B(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_758), .B(n_801), .Y(n_830) );
CKINVDCx16_ASAP7_75t_R g801 ( .A(n_759), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
OAI222xp33_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_800), .B1(n_802), .B2(n_823), .C1(n_825), .C2(n_828), .Y(n_767) );
INVx1_ASAP7_75t_L g799 ( .A(n_769), .Y(n_799) );
AND2x2_ASAP7_75t_SL g769 ( .A(n_770), .B(n_784), .Y(n_769) );
NOR3xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_775), .C(n_780), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_777), .B1(n_778), .B2(n_779), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_777), .A2(n_779), .B1(n_807), .B2(n_808), .Y(n_806) );
NOR3xp33_ASAP7_75t_SL g784 ( .A(n_785), .B(n_788), .C(n_794), .Y(n_784) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g824 ( .A(n_804), .Y(n_824) );
AND4x1_ASAP7_75t_L g804 ( .A(n_805), .B(n_809), .C(n_815), .D(n_819), .Y(n_804) );
INVx3_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_826), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_829), .Y(n_828) );
endmodule