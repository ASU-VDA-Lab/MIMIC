module real_aes_9014_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_182;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g418 ( .A(n_0), .Y(n_418) );
INVx1_ASAP7_75t_L g497 ( .A(n_1), .Y(n_497) );
INVx1_ASAP7_75t_L g129 ( .A(n_2), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_3), .A2(n_36), .B1(n_154), .B2(n_443), .Y(n_466) );
AOI21xp33_ASAP7_75t_L g161 ( .A1(n_4), .A2(n_145), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_5), .B(n_143), .Y(n_509) );
AND2x6_ASAP7_75t_L g122 ( .A(n_6), .B(n_123), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_7), .A2(n_232), .B(n_233), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_8), .B(n_37), .Y(n_419) );
INVx1_ASAP7_75t_L g167 ( .A(n_9), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_10), .B(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g491 ( .A(n_11), .Y(n_491) );
INVx1_ASAP7_75t_L g114 ( .A(n_12), .Y(n_114) );
INVx1_ASAP7_75t_L g238 ( .A(n_13), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_14), .B(n_135), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_15), .B(n_110), .Y(n_480) );
AO32x2_ASAP7_75t_L g464 ( .A1(n_16), .A2(n_109), .A3(n_143), .B1(n_445), .B2(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_17), .B(n_154), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_18), .B(n_150), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_19), .B(n_110), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_20), .A2(n_48), .B1(n_154), .B2(n_443), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_21), .B(n_145), .Y(n_195) );
OAI222xp33_ASAP7_75t_L g99 ( .A1(n_22), .A2(n_100), .B1(n_699), .B2(n_700), .C1(n_705), .C2(n_710), .Y(n_99) );
INVx1_ASAP7_75t_L g699 ( .A(n_22), .Y(n_699) );
AOI22xp33_ASAP7_75t_SL g444 ( .A1(n_23), .A2(n_73), .B1(n_135), .B2(n_154), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_24), .B(n_154), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_25), .B(n_157), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_26), .A2(n_236), .B(n_237), .C(n_239), .Y(n_235) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_27), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_28), .B(n_140), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_29), .B(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g182 ( .A(n_30), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_31), .B(n_140), .Y(n_436) );
INVx2_ASAP7_75t_L g120 ( .A(n_32), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_33), .B(n_154), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_34), .B(n_140), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_35), .A2(n_122), .B(n_125), .C(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g180 ( .A(n_38), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_39), .B(n_133), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_40), .B(n_154), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_41), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_42), .A2(n_83), .B1(n_202), .B2(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_43), .B(n_154), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_44), .B(n_154), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g183 ( .A(n_45), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_46), .B(n_496), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_47), .B(n_145), .Y(n_226) );
AOI22xp33_ASAP7_75t_SL g484 ( .A1(n_49), .A2(n_59), .B1(n_135), .B2(n_154), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_50), .A2(n_125), .B1(n_135), .B2(n_178), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_51), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_52), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_53), .B(n_154), .Y(n_451) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_54), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_55), .B(n_154), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_56), .A2(n_153), .B(n_165), .C(n_166), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_57), .Y(n_215) );
INVx1_ASAP7_75t_L g163 ( .A(n_58), .Y(n_163) );
INVx1_ASAP7_75t_L g123 ( .A(n_60), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_61), .B(n_154), .Y(n_498) );
INVx1_ASAP7_75t_L g113 ( .A(n_62), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_63), .Y(n_716) );
AO32x2_ASAP7_75t_L g440 ( .A1(n_64), .A2(n_143), .A3(n_218), .B1(n_441), .B2(n_445), .Y(n_440) );
INVx1_ASAP7_75t_L g516 ( .A(n_65), .Y(n_516) );
INVx1_ASAP7_75t_L g431 ( .A(n_66), .Y(n_431) );
A2O1A1Ixp33_ASAP7_75t_SL g149 ( .A1(n_67), .A2(n_150), .B(n_151), .C(n_153), .Y(n_149) );
INVxp67_ASAP7_75t_L g152 ( .A(n_68), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_69), .B(n_135), .Y(n_432) );
INVx1_ASAP7_75t_L g715 ( .A(n_70), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_71), .Y(n_185) );
INVx1_ASAP7_75t_L g208 ( .A(n_72), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_74), .A2(n_122), .B(n_125), .C(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_75), .B(n_443), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_76), .B(n_135), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_77), .B(n_130), .Y(n_198) );
INVx2_ASAP7_75t_L g111 ( .A(n_78), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_79), .B(n_150), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_80), .B(n_135), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g124 ( .A1(n_81), .A2(n_122), .B(n_125), .C(n_128), .Y(n_124) );
OR2x2_ASAP7_75t_L g416 ( .A(n_82), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g698 ( .A(n_82), .Y(n_698) );
OR2x2_ASAP7_75t_L g719 ( .A(n_82), .B(n_709), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_84), .A2(n_97), .B1(n_135), .B2(n_136), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_85), .B(n_140), .Y(n_168) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_86), .A2(n_99), .B1(n_711), .B2(n_720), .C1(n_730), .C2(n_736), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_86), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_86), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_87), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_88), .A2(n_122), .B(n_125), .C(n_221), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_89), .Y(n_228) );
INVx1_ASAP7_75t_L g148 ( .A(n_90), .Y(n_148) );
CKINVDCx16_ASAP7_75t_R g234 ( .A(n_91), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_92), .B(n_130), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_93), .B(n_135), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_94), .B(n_143), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_95), .A2(n_145), .B(n_146), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_96), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OAI22xp5_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_414), .B1(n_420), .B2(n_695), .Y(n_101) );
INVx1_ASAP7_75t_L g703 ( .A(n_102), .Y(n_703) );
BUFx2_ASAP7_75t_L g724 ( .A(n_102), .Y(n_724) );
NAND2x1_ASAP7_75t_L g102 ( .A(n_103), .B(n_330), .Y(n_102) );
NOR5xp2_ASAP7_75t_L g103 ( .A(n_104), .B(n_253), .C(n_285), .D(n_300), .E(n_317), .Y(n_103) );
A2O1A1Ixp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_169), .B(n_190), .C(n_241), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_141), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_106), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_106), .B(n_305), .Y(n_368) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_107), .B(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_107), .B(n_187), .Y(n_254) );
AND2x2_ASAP7_75t_L g295 ( .A(n_107), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_107), .B(n_264), .Y(n_299) );
OR2x2_ASAP7_75t_L g336 ( .A(n_107), .B(n_175), .Y(n_336) );
INVx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g174 ( .A(n_108), .B(n_175), .Y(n_174) );
INVx3_ASAP7_75t_L g244 ( .A(n_108), .Y(n_244) );
OR2x2_ASAP7_75t_L g407 ( .A(n_108), .B(n_247), .Y(n_407) );
AO21x2_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_115), .B(n_137), .Y(n_108) );
AO21x2_ASAP7_75t_L g175 ( .A1(n_109), .A2(n_176), .B(n_184), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_109), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g203 ( .A(n_109), .Y(n_203) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_110), .Y(n_143) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_111), .B(n_112), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OAI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_117), .B(n_124), .Y(n_115) );
OAI22xp33_ASAP7_75t_L g176 ( .A1(n_117), .A2(n_155), .B1(n_177), .B2(n_183), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_117), .A2(n_208), .B(n_209), .Y(n_207) );
NAND2x1p5_ASAP7_75t_L g117 ( .A(n_118), .B(n_122), .Y(n_117) );
AND2x4_ASAP7_75t_L g145 ( .A(n_118), .B(n_122), .Y(n_145) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
INVx1_ASAP7_75t_L g496 ( .A(n_119), .Y(n_496) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g126 ( .A(n_120), .Y(n_126) );
INVx1_ASAP7_75t_L g136 ( .A(n_120), .Y(n_136) );
INVx1_ASAP7_75t_L g127 ( .A(n_121), .Y(n_127) );
INVx3_ASAP7_75t_L g131 ( .A(n_121), .Y(n_131) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_121), .Y(n_133) );
INVx1_ASAP7_75t_L g150 ( .A(n_121), .Y(n_150) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_121), .Y(n_179) );
INVx4_ASAP7_75t_SL g155 ( .A(n_122), .Y(n_155) );
OAI21xp5_ASAP7_75t_L g429 ( .A1(n_122), .A2(n_430), .B(n_433), .Y(n_429) );
BUFx3_ASAP7_75t_L g445 ( .A(n_122), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_122), .A2(n_450), .B(n_454), .Y(n_449) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_122), .A2(n_490), .B(n_494), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_122), .A2(n_503), .B(n_506), .Y(n_502) );
INVx5_ASAP7_75t_L g147 ( .A(n_125), .Y(n_147) );
AND2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
BUFx3_ASAP7_75t_L g202 ( .A(n_126), .Y(n_202) );
INVx1_ASAP7_75t_L g443 ( .A(n_126), .Y(n_443) );
O2A1O1Ixp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_130), .B(n_132), .C(n_134), .Y(n_128) );
O2A1O1Ixp5_ASAP7_75t_SL g430 ( .A1(n_130), .A2(n_153), .B(n_431), .C(n_432), .Y(n_430) );
INVx2_ASAP7_75t_L g467 ( .A(n_130), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_130), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_130), .A2(n_513), .B(n_514), .Y(n_512) );
INVx5_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_131), .B(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_131), .B(n_167), .Y(n_166) );
OAI22xp5_ASAP7_75t_SL g441 ( .A1(n_131), .A2(n_133), .B1(n_442), .B2(n_444), .Y(n_441) );
INVx2_ASAP7_75t_L g165 ( .A(n_133), .Y(n_165) );
INVx4_ASAP7_75t_L g224 ( .A(n_133), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_133), .A2(n_466), .B1(n_467), .B2(n_468), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_133), .A2(n_467), .B1(n_483), .B2(n_484), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_134), .A2(n_491), .B(n_492), .C(n_493), .Y(n_490) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_139), .B(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_139), .B(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g218 ( .A(n_140), .Y(n_218) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_140), .A2(n_231), .B(n_240), .Y(n_230) );
OA21x2_ASAP7_75t_L g428 ( .A1(n_140), .A2(n_429), .B(n_436), .Y(n_428) );
OA21x2_ASAP7_75t_L g448 ( .A1(n_140), .A2(n_449), .B(n_457), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_141), .A2(n_310), .B1(n_311), .B2(n_314), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_141), .B(n_244), .Y(n_393) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_159), .Y(n_141) );
AND2x2_ASAP7_75t_L g189 ( .A(n_142), .B(n_175), .Y(n_189) );
AND2x2_ASAP7_75t_L g246 ( .A(n_142), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g251 ( .A(n_142), .Y(n_251) );
INVx3_ASAP7_75t_L g264 ( .A(n_142), .Y(n_264) );
OR2x2_ASAP7_75t_L g284 ( .A(n_142), .B(n_247), .Y(n_284) );
AND2x2_ASAP7_75t_L g303 ( .A(n_142), .B(n_160), .Y(n_303) );
BUFx2_ASAP7_75t_L g335 ( .A(n_142), .Y(n_335) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_156), .Y(n_142) );
INVx4_ASAP7_75t_L g158 ( .A(n_143), .Y(n_158) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_143), .A2(n_502), .B(n_509), .Y(n_501) );
BUFx2_ASAP7_75t_L g232 ( .A(n_145), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_149), .C(n_155), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g162 ( .A1(n_147), .A2(n_155), .B(n_163), .C(n_164), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_147), .A2(n_155), .B(n_234), .C(n_235), .Y(n_233) );
INVx1_ASAP7_75t_L g453 ( .A(n_150), .Y(n_453) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_154), .Y(n_225) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_157), .A2(n_161), .B(n_168), .Y(n_160) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_SL g204 ( .A(n_158), .B(n_205), .Y(n_204) );
NAND3xp33_ASAP7_75t_L g481 ( .A(n_158), .B(n_445), .C(n_482), .Y(n_481) );
AO21x1_ASAP7_75t_L g571 ( .A1(n_158), .A2(n_482), .B(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g250 ( .A(n_159), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
BUFx2_ASAP7_75t_L g173 ( .A(n_160), .Y(n_173) );
INVx2_ASAP7_75t_L g188 ( .A(n_160), .Y(n_188) );
OR2x2_ASAP7_75t_L g266 ( .A(n_160), .B(n_247), .Y(n_266) );
AND2x2_ASAP7_75t_L g296 ( .A(n_160), .B(n_175), .Y(n_296) );
AND2x2_ASAP7_75t_L g313 ( .A(n_160), .B(n_244), .Y(n_313) );
AND2x2_ASAP7_75t_L g353 ( .A(n_160), .B(n_264), .Y(n_353) );
AND2x2_ASAP7_75t_SL g389 ( .A(n_160), .B(n_189), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_165), .A2(n_455), .B(n_456), .Y(n_454) );
O2A1O1Ixp5_ASAP7_75t_L g515 ( .A1(n_165), .A2(n_495), .B(n_516), .C(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NAND2xp33_ASAP7_75t_SL g170 ( .A(n_171), .B(n_186), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_174), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_172), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
OAI21xp33_ASAP7_75t_L g327 ( .A1(n_173), .A2(n_189), .B(n_328), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_173), .B(n_175), .Y(n_383) );
AND2x2_ASAP7_75t_L g319 ( .A(n_174), .B(n_320), .Y(n_319) );
INVx3_ASAP7_75t_L g247 ( .A(n_175), .Y(n_247) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_175), .Y(n_345) );
OAI22xp5_ASAP7_75t_SL g178 ( .A1(n_179), .A2(n_180), .B1(n_181), .B2(n_182), .Y(n_178) );
INVx2_ASAP7_75t_L g181 ( .A(n_179), .Y(n_181) );
INVx4_ASAP7_75t_L g236 ( .A(n_179), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_186), .B(n_244), .Y(n_412) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_187), .A2(n_355), .B1(n_356), .B2(n_361), .Y(n_354) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
AND2x2_ASAP7_75t_L g245 ( .A(n_188), .B(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g283 ( .A(n_188), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_SL g320 ( .A(n_188), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_189), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g374 ( .A(n_189), .Y(n_374) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_216), .Y(n_191) );
INVx4_ASAP7_75t_L g260 ( .A(n_192), .Y(n_260) );
AND2x2_ASAP7_75t_L g338 ( .A(n_192), .B(n_305), .Y(n_338) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_206), .Y(n_192) );
INVx3_ASAP7_75t_L g257 ( .A(n_193), .Y(n_257) );
AND2x2_ASAP7_75t_L g271 ( .A(n_193), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g275 ( .A(n_193), .Y(n_275) );
INVx2_ASAP7_75t_L g289 ( .A(n_193), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_193), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g346 ( .A(n_193), .B(n_341), .Y(n_346) );
AND2x2_ASAP7_75t_L g411 ( .A(n_193), .B(n_381), .Y(n_411) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_204), .Y(n_193) );
AOI21xp5_ASAP7_75t_SL g194 ( .A1(n_195), .A2(n_196), .B(n_203), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_200), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_200), .A2(n_211), .B(n_212), .Y(n_210) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g239 ( .A(n_202), .Y(n_239) );
INVx1_ASAP7_75t_L g213 ( .A(n_203), .Y(n_213) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_203), .A2(n_489), .B(n_499), .Y(n_488) );
OA21x2_ASAP7_75t_L g510 ( .A1(n_203), .A2(n_511), .B(n_518), .Y(n_510) );
AND2x2_ASAP7_75t_L g252 ( .A(n_206), .B(n_230), .Y(n_252) );
INVx2_ASAP7_75t_L g272 ( .A(n_206), .Y(n_272) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_213), .B(n_214), .Y(n_206) );
INVx1_ASAP7_75t_L g277 ( .A(n_216), .Y(n_277) );
AND2x2_ASAP7_75t_L g323 ( .A(n_216), .B(n_271), .Y(n_323) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_229), .Y(n_216) );
INVx2_ASAP7_75t_L g262 ( .A(n_217), .Y(n_262) );
INVx1_ASAP7_75t_L g270 ( .A(n_217), .Y(n_270) );
AND2x2_ASAP7_75t_L g288 ( .A(n_217), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_217), .B(n_272), .Y(n_326) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_227), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_226), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_225), .Y(n_221) );
AND2x2_ASAP7_75t_L g305 ( .A(n_229), .B(n_262), .Y(n_305) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g258 ( .A(n_230), .Y(n_258) );
AND2x2_ASAP7_75t_L g341 ( .A(n_230), .B(n_272), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_236), .B(n_238), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_236), .A2(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g493 ( .A(n_236), .Y(n_493) );
OAI21xp5_ASAP7_75t_SL g241 ( .A1(n_242), .A2(n_248), .B(n_252), .Y(n_241) );
INVx1_ASAP7_75t_SL g286 ( .A(n_242), .Y(n_286) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_245), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_243), .B(n_250), .Y(n_343) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g292 ( .A(n_244), .B(n_247), .Y(n_292) );
AND2x2_ASAP7_75t_L g321 ( .A(n_244), .B(n_265), .Y(n_321) );
OR2x2_ASAP7_75t_L g324 ( .A(n_244), .B(n_284), .Y(n_324) );
AOI222xp33_ASAP7_75t_L g388 ( .A1(n_245), .A2(n_337), .B1(n_389), .B2(n_390), .C1(n_392), .C2(n_394), .Y(n_388) );
BUFx2_ASAP7_75t_L g302 ( .A(n_247), .Y(n_302) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g291 ( .A(n_250), .B(n_292), .Y(n_291) );
INVx3_ASAP7_75t_SL g308 ( .A(n_250), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_250), .B(n_302), .Y(n_362) );
AND2x2_ASAP7_75t_L g297 ( .A(n_252), .B(n_257), .Y(n_297) );
INVx1_ASAP7_75t_L g316 ( .A(n_252), .Y(n_316) );
OAI221xp5_ASAP7_75t_SL g253 ( .A1(n_254), .A2(n_255), .B1(n_259), .B2(n_263), .C(n_267), .Y(n_253) );
OR2x2_ASAP7_75t_L g325 ( .A(n_255), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
AND2x2_ASAP7_75t_L g310 ( .A(n_257), .B(n_280), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_257), .B(n_270), .Y(n_350) );
AND2x2_ASAP7_75t_L g355 ( .A(n_257), .B(n_305), .Y(n_355) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_257), .Y(n_365) );
NAND2x1_ASAP7_75t_SL g376 ( .A(n_257), .B(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g261 ( .A(n_258), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g281 ( .A(n_258), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_258), .B(n_276), .Y(n_307) );
INVx1_ASAP7_75t_L g373 ( .A(n_258), .Y(n_373) );
INVx1_ASAP7_75t_L g348 ( .A(n_259), .Y(n_348) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx1_ASAP7_75t_L g360 ( .A(n_260), .Y(n_360) );
NOR2xp67_ASAP7_75t_L g372 ( .A(n_260), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g377 ( .A(n_261), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_261), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g280 ( .A(n_262), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_262), .B(n_272), .Y(n_293) );
INVx1_ASAP7_75t_L g359 ( .A(n_262), .Y(n_359) );
INVx1_ASAP7_75t_L g380 ( .A(n_263), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OAI21xp5_ASAP7_75t_SL g267 ( .A1(n_268), .A2(n_273), .B(n_282), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
AND2x2_ASAP7_75t_L g413 ( .A(n_269), .B(n_346), .Y(n_413) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g381 ( .A(n_270), .B(n_341), .Y(n_381) );
AOI32xp33_ASAP7_75t_L g294 ( .A1(n_271), .A2(n_277), .A3(n_295), .B1(n_297), .B2(n_298), .Y(n_294) );
AOI322xp5_ASAP7_75t_L g396 ( .A1(n_271), .A2(n_303), .A3(n_386), .B1(n_397), .B2(n_398), .C1(n_399), .C2(n_401), .Y(n_396) );
INVx2_ASAP7_75t_L g276 ( .A(n_272), .Y(n_276) );
INVx1_ASAP7_75t_L g386 ( .A(n_272), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_277), .B1(n_278), .B2(n_279), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_274), .B(n_280), .Y(n_329) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_275), .B(n_341), .Y(n_391) );
INVx1_ASAP7_75t_L g278 ( .A(n_276), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_276), .B(n_305), .Y(n_395) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_284), .B(n_379), .Y(n_378) );
OAI221xp5_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_287), .B1(n_290), .B2(n_293), .C(n_294), .Y(n_285) );
OR2x2_ASAP7_75t_L g306 ( .A(n_287), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g315 ( .A(n_287), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g340 ( .A(n_288), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g344 ( .A(n_298), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OAI221xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_304), .B1(n_306), .B2(n_308), .C(n_309), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_302), .A2(n_333), .B1(n_337), .B2(n_338), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_303), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g408 ( .A(n_303), .Y(n_408) );
INVx1_ASAP7_75t_L g402 ( .A(n_305), .Y(n_402) );
INVx1_ASAP7_75t_SL g337 ( .A(n_306), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_308), .B(n_336), .Y(n_398) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_313), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g379 ( .A(n_313), .Y(n_379) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
OAI221xp5_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_322), .B1(n_324), .B2(n_325), .C(n_327), .Y(n_317) );
NOR2xp33_ASAP7_75t_SL g318 ( .A(n_319), .B(n_321), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_319), .A2(n_337), .B1(n_383), .B2(n_384), .Y(n_382) );
CKINVDCx14_ASAP7_75t_R g322 ( .A(n_323), .Y(n_322) );
OAI21xp33_ASAP7_75t_L g401 ( .A1(n_324), .A2(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NOR3xp33_ASAP7_75t_SL g330 ( .A(n_331), .B(n_363), .C(n_387), .Y(n_330) );
NAND4xp25_ASAP7_75t_L g331 ( .A(n_332), .B(n_339), .C(n_347), .D(n_354), .Y(n_331) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g410 ( .A(n_335), .Y(n_410) );
INVx3_ASAP7_75t_SL g404 ( .A(n_336), .Y(n_404) );
OR2x2_ASAP7_75t_L g409 ( .A(n_336), .B(n_410), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_342), .B1(n_344), .B2(n_346), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_341), .B(n_359), .Y(n_400) );
INVxp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI21xp5_ASAP7_75t_SL g347 ( .A1(n_348), .A2(n_349), .B(n_351), .Y(n_347) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
INVxp67_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI211xp5_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_366), .B(n_369), .C(n_382), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g397 ( .A(n_368), .Y(n_397) );
AOI222xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_374), .B1(n_375), .B2(n_378), .C1(n_380), .C2(n_381), .Y(n_369) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND4xp25_ASAP7_75t_SL g406 ( .A(n_379), .B(n_407), .C(n_408), .D(n_409), .Y(n_406) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND3xp33_ASAP7_75t_SL g387 ( .A(n_388), .B(n_396), .C(n_405), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_411), .B1(n_412), .B2(n_413), .Y(n_405) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g702 ( .A(n_415), .Y(n_702) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g697 ( .A(n_417), .B(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g709 ( .A(n_417), .Y(n_709) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx1_ASAP7_75t_L g704 ( .A(n_420), .Y(n_704) );
OR2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_616), .Y(n_420) );
NAND3xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_565), .C(n_607), .Y(n_421) );
AOI211xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_474), .B(n_519), .C(n_541), .Y(n_422) );
OAI211xp5_ASAP7_75t_SL g423 ( .A1(n_424), .A2(n_437), .B(n_458), .C(n_469), .Y(n_423) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_425), .B(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g628 ( .A(n_425), .B(n_545), .Y(n_628) );
BUFx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g530 ( .A(n_426), .B(n_461), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_426), .B(n_448), .Y(n_647) );
INVx1_ASAP7_75t_L g665 ( .A(n_426), .Y(n_665) );
AND2x2_ASAP7_75t_L g674 ( .A(n_426), .B(n_562), .Y(n_674) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g557 ( .A(n_427), .B(n_448), .Y(n_557) );
AND2x2_ASAP7_75t_L g615 ( .A(n_427), .B(n_562), .Y(n_615) );
INVx1_ASAP7_75t_L g659 ( .A(n_427), .Y(n_659) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g536 ( .A(n_428), .B(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g544 ( .A(n_428), .Y(n_544) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_428), .Y(n_584) );
INVxp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_446), .Y(n_438) );
AND2x2_ASAP7_75t_L g523 ( .A(n_439), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g556 ( .A(n_439), .Y(n_556) );
OR2x2_ASAP7_75t_L g682 ( .A(n_439), .B(n_683), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_439), .B(n_448), .Y(n_686) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g461 ( .A(n_440), .Y(n_461) );
INVx1_ASAP7_75t_L g472 ( .A(n_440), .Y(n_472) );
AND2x2_ASAP7_75t_L g545 ( .A(n_440), .B(n_463), .Y(n_545) );
AND2x2_ASAP7_75t_L g585 ( .A(n_440), .B(n_464), .Y(n_585) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_445), .A2(n_512), .B(n_515), .Y(n_511) );
INVxp67_ASAP7_75t_L g627 ( .A(n_446), .Y(n_627) );
AND2x4_ASAP7_75t_L g652 ( .A(n_446), .B(n_545), .Y(n_652) );
BUFx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_SL g543 ( .A(n_447), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g462 ( .A(n_448), .B(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g531 ( .A(n_448), .B(n_464), .Y(n_531) );
INVx1_ASAP7_75t_L g537 ( .A(n_448), .Y(n_537) );
INVx2_ASAP7_75t_L g563 ( .A(n_448), .Y(n_563) );
AND2x2_ASAP7_75t_L g579 ( .A(n_448), .B(n_580), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B(n_453), .Y(n_450) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_459), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx2_ASAP7_75t_L g534 ( .A(n_461), .Y(n_534) );
AND2x2_ASAP7_75t_L g642 ( .A(n_461), .B(n_463), .Y(n_642) );
AND2x2_ASAP7_75t_L g559 ( .A(n_462), .B(n_544), .Y(n_559) );
AND2x2_ASAP7_75t_L g658 ( .A(n_462), .B(n_659), .Y(n_658) );
NOR2xp67_ASAP7_75t_L g580 ( .A(n_463), .B(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g683 ( .A(n_463), .B(n_544), .Y(n_683) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx2_ASAP7_75t_L g473 ( .A(n_464), .Y(n_473) );
AND2x2_ASAP7_75t_L g562 ( .A(n_464), .B(n_563), .Y(n_562) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_467), .A2(n_495), .B(n_497), .C(n_498), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_467), .A2(n_507), .B(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
AND2x2_ASAP7_75t_L g608 ( .A(n_471), .B(n_543), .Y(n_608) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_472), .B(n_544), .Y(n_593) );
INVx2_ASAP7_75t_L g592 ( .A(n_473), .Y(n_592) );
OAI222xp33_ASAP7_75t_L g596 ( .A1(n_473), .A2(n_536), .B1(n_597), .B2(n_599), .C1(n_600), .C2(n_603), .Y(n_596) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_485), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g521 ( .A(n_478), .Y(n_521) );
OR2x2_ASAP7_75t_L g632 ( .A(n_478), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx3_ASAP7_75t_L g554 ( .A(n_479), .Y(n_554) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_479), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g611 ( .A(n_479), .B(n_525), .Y(n_611) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g572 ( .A(n_480), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_485), .A2(n_575), .B1(n_614), .B2(n_615), .Y(n_613) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_500), .Y(n_485) );
INVx3_ASAP7_75t_L g547 ( .A(n_486), .Y(n_547) );
OR2x2_ASAP7_75t_L g680 ( .A(n_486), .B(n_556), .Y(n_680) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g553 ( .A(n_487), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g569 ( .A(n_487), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g577 ( .A(n_487), .B(n_525), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_487), .B(n_501), .Y(n_633) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g524 ( .A(n_488), .B(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g528 ( .A(n_488), .B(n_501), .Y(n_528) );
AND2x2_ASAP7_75t_L g604 ( .A(n_488), .B(n_551), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_488), .B(n_510), .Y(n_644) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_500), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g560 ( .A(n_500), .B(n_521), .Y(n_560) );
AND2x2_ASAP7_75t_L g564 ( .A(n_500), .B(n_554), .Y(n_564) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_510), .Y(n_500) );
INVx3_ASAP7_75t_L g525 ( .A(n_501), .Y(n_525) );
AND2x2_ASAP7_75t_L g550 ( .A(n_501), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g685 ( .A(n_501), .B(n_668), .Y(n_685) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_510), .Y(n_539) );
INVx2_ASAP7_75t_L g551 ( .A(n_510), .Y(n_551) );
AND2x2_ASAP7_75t_L g595 ( .A(n_510), .B(n_571), .Y(n_595) );
INVx1_ASAP7_75t_L g638 ( .A(n_510), .Y(n_638) );
OR2x2_ASAP7_75t_L g669 ( .A(n_510), .B(n_571), .Y(n_669) );
AND2x2_ASAP7_75t_L g689 ( .A(n_510), .B(n_525), .Y(n_689) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_522), .B(n_526), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g527 ( .A(n_521), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_521), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g646 ( .A(n_523), .Y(n_646) );
INVx2_ASAP7_75t_SL g540 ( .A(n_524), .Y(n_540) );
AND2x2_ASAP7_75t_L g660 ( .A(n_524), .B(n_554), .Y(n_660) );
INVx2_ASAP7_75t_L g606 ( .A(n_525), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_525), .B(n_638), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_529), .B1(n_532), .B2(n_538), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_528), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g694 ( .A(n_528), .Y(n_694) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g619 ( .A(n_530), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_530), .B(n_562), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_531), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g635 ( .A(n_531), .B(n_584), .Y(n_635) );
INVx2_ASAP7_75t_L g691 ( .A(n_531), .Y(n_691) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
AND2x2_ASAP7_75t_L g561 ( .A(n_534), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_534), .B(n_579), .Y(n_612) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_536), .B(n_556), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g673 ( .A(n_539), .Y(n_673) );
O2A1O1Ixp33_ASAP7_75t_SL g623 ( .A1(n_540), .A2(n_624), .B(n_626), .C(n_629), .Y(n_623) );
OR2x2_ASAP7_75t_L g650 ( .A(n_540), .B(n_554), .Y(n_650) );
OAI221xp5_ASAP7_75t_SL g541 ( .A1(n_542), .A2(n_546), .B1(n_548), .B2(n_555), .C(n_558), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_543), .B(n_545), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_543), .B(n_592), .Y(n_599) );
AND2x2_ASAP7_75t_L g641 ( .A(n_543), .B(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g677 ( .A(n_543), .Y(n_677) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_544), .Y(n_568) );
INVx1_ASAP7_75t_L g581 ( .A(n_544), .Y(n_581) );
NOR2xp67_ASAP7_75t_L g601 ( .A(n_547), .B(n_602), .Y(n_601) );
INVxp67_ASAP7_75t_L g655 ( .A(n_547), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_547), .B(n_595), .Y(n_671) );
INVx2_ASAP7_75t_L g657 ( .A(n_548), .Y(n_657) );
OR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_552), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g598 ( .A(n_550), .B(n_569), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_L g607 ( .A1(n_550), .A2(n_566), .B(n_608), .C(n_609), .Y(n_607) );
AND2x2_ASAP7_75t_L g576 ( .A(n_551), .B(n_571), .Y(n_576) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_555), .B(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
OR2x2_ASAP7_75t_L g624 ( .A(n_556), .B(n_625), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B1(n_561), .B2(n_564), .Y(n_558) );
INVx1_ASAP7_75t_L g678 ( .A(n_560), .Y(n_678) );
INVx1_ASAP7_75t_L g625 ( .A(n_562), .Y(n_625) );
INVx1_ASAP7_75t_L g676 ( .A(n_564), .Y(n_676) );
AOI211xp5_ASAP7_75t_SL g565 ( .A1(n_566), .A2(n_569), .B(n_573), .C(n_596), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g588 ( .A(n_568), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g639 ( .A(n_569), .Y(n_639) );
AND2x2_ASAP7_75t_L g688 ( .A(n_569), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OAI21xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_578), .B(n_586), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx2_ASAP7_75t_L g602 ( .A(n_576), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_576), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g594 ( .A(n_577), .B(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g670 ( .A(n_577), .Y(n_670) );
OAI32xp33_ASAP7_75t_L g681 ( .A1(n_577), .A2(n_629), .A3(n_636), .B1(n_677), .B2(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_SL g578 ( .A(n_579), .B(n_582), .Y(n_578) );
INVx1_ASAP7_75t_SL g649 ( .A(n_579), .Y(n_649) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_SL g589 ( .A(n_585), .Y(n_589) );
OAI21xp33_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_590), .B(n_594), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI22xp33_ASAP7_75t_L g661 ( .A1(n_588), .A2(n_636), .B1(n_662), .B2(n_664), .Y(n_661) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_592), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g629 ( .A(n_595), .Y(n_629) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2x1p5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g622 ( .A(n_606), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_612), .B(n_613), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_615), .A2(n_657), .B1(n_658), .B2(n_660), .C(n_661), .Y(n_656) );
NAND5xp2_ASAP7_75t_L g616 ( .A(n_617), .B(n_640), .C(n_656), .D(n_666), .E(n_684), .Y(n_616) );
AOI211xp5_ASAP7_75t_SL g617 ( .A1(n_618), .A2(n_620), .B(n_623), .C(n_630), .Y(n_617) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g687 ( .A(n_624), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_634), .B2(n_636), .Y(n_630) );
INVx1_ASAP7_75t_SL g663 ( .A(n_633), .Y(n_663) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI322xp33_ASAP7_75t_L g645 ( .A1(n_636), .A2(n_646), .A3(n_647), .B1(n_648), .B2(n_649), .C1(n_650), .C2(n_651), .Y(n_645) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g648 ( .A(n_638), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_638), .B(n_663), .Y(n_662) );
AOI211xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_643), .B(n_645), .C(n_653), .Y(n_640) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_649), .A2(n_676), .B1(n_677), .B2(n_678), .Y(n_675) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g692 ( .A(n_659), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_674), .B1(n_675), .B2(n_679), .C(n_681), .Y(n_666) );
OAI211xp5_ASAP7_75t_SL g667 ( .A1(n_668), .A2(n_670), .B(n_671), .C(n_672), .Y(n_667) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g693 ( .A(n_669), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .B1(n_687), .B2(n_688), .C(n_690), .Y(n_684) );
AOI21xp33_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_692), .B(n_693), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_695), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_701) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NOR2x2_ASAP7_75t_L g708 ( .A(n_698), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
NAND2xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_717), .Y(n_712) );
NOR2xp33_ASAP7_75t_SL g713 ( .A(n_714), .B(n_716), .Y(n_713) );
INVx1_ASAP7_75t_SL g735 ( .A(n_714), .Y(n_735) );
INVx1_ASAP7_75t_L g734 ( .A(n_716), .Y(n_734) );
OA21x2_ASAP7_75t_L g737 ( .A1(n_716), .A2(n_728), .B(n_735), .Y(n_737) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_719), .Y(n_726) );
BUFx2_ASAP7_75t_L g728 ( .A(n_719), .Y(n_728) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_726), .B(n_727), .Y(n_721) );
INVx1_ASAP7_75t_L g725 ( .A(n_724), .Y(n_725) );
NOR2xp33_ASAP7_75t_SL g727 ( .A(n_728), .B(n_729), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_731), .Y(n_730) );
CKINVDCx6p67_ASAP7_75t_R g731 ( .A(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
endmodule