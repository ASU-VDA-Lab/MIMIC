module fake_jpeg_1796_n_176 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_176);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx8_ASAP7_75t_SL g47 ( 
.A(n_34),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_63),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_64),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_44),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_0),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_48),
.B1(n_49),
.B2(n_55),
.Y(n_75)
);

OAI22x1_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_82),
.B1(n_64),
.B2(n_52),
.Y(n_94)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_45),
.C(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_78),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_53),
.B1(n_58),
.B2(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_81),
.B(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_84),
.B(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_81),
.B(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_68),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_90),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_67),
.B1(n_63),
.B2(n_56),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_95),
.B1(n_86),
.B2(n_98),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_80),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_49),
.B(n_1),
.C(n_2),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_3),
.Y(n_100)
);

BUFx6f_ASAP7_75t_SL g92 ( 
.A(n_72),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_73),
.B1(n_58),
.B2(n_53),
.Y(n_110)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

OR2x2_ASAP7_75t_SL g96 ( 
.A(n_78),
.B(n_52),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_97),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_0),
.B(n_1),
.Y(n_99)
);

AOI32xp33_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_9),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_62),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_104),
.B(n_12),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_106),
.B(n_118),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_114),
.B1(n_42),
.B2(n_37),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_64),
.B1(n_77),
.B2(n_46),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_112),
.B1(n_25),
.B2(n_24),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_46),
.B1(n_50),
.B2(n_6),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_50),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_28),
.C(n_27),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_96),
.A2(n_23),
.B1(n_39),
.B2(n_38),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_115),
.A2(n_117),
.B1(n_92),
.B2(n_22),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_86),
.B(n_8),
.Y(n_118)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_125),
.B1(n_126),
.B2(n_131),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_98),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_121),
.B(n_137),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_128),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_129),
.C(n_133),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_35),
.B(n_32),
.C(n_29),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_11),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_132),
.B(n_136),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_138),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_100),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_111),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_14),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_112),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_145),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_116),
.B(n_16),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_152),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_116),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_15),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_146),
.B(n_147),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_18),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_151),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_18),
.B(n_19),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_155),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_130),
.C(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_141),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_159),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_153),
.B1(n_142),
.B2(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_161),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_159),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_160),
.B(n_154),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_162),
.C(n_168),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_162),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_143),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_169),
.B(n_165),
.Y(n_174)
);

AOI221xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_156),
.B1(n_163),
.B2(n_143),
.C(n_148),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_144),
.Y(n_176)
);


endmodule