module fake_jpeg_23172_n_84 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_84);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_84;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx4_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_6),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_22),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_23),
.Y(n_24)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_14),
.B1(n_15),
.B2(n_11),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_15),
.B1(n_18),
.B2(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_12),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_12),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_11),
.B1(n_9),
.B2(n_22),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_31),
.B1(n_25),
.B2(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

AOI32xp33_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_25),
.A3(n_26),
.B1(n_13),
.B2(n_3),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_24),
.C(n_27),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_26),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_42),
.B1(n_10),
.B2(n_37),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_24),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_48),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_49),
.B(n_53),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_38),
.C(n_33),
.Y(n_51)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_48),
.C(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_32),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_56),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_64),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_65),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_16),
.C(n_36),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_21),
.C(n_20),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_25),
.C(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_66),
.B(n_68),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_71),
.Y(n_77)
);

AO221x1_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_45),
.B1(n_28),
.B2(n_2),
.C(n_3),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_16),
.B(n_1),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_72),
.B(n_45),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_59),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_74),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_59),
.Y(n_76)
);

NAND4xp25_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_67),
.C(n_16),
.D(n_28),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_6),
.B1(n_7),
.B2(n_28),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_79),
.A2(n_77),
.B1(n_1),
.B2(n_2),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_81),
.A2(n_80),
.B1(n_78),
.B2(n_4),
.Y(n_82)
);

NAND4xp25_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_73),
.C(n_28),
.D(n_0),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_0),
.Y(n_84)
);


endmodule