module fake_jpeg_2795_n_545 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_545);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_545;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_293;
wire n_38;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_441;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g119 ( 
.A(n_45),
.Y(n_119)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_53),
.Y(n_101)
);

HAxp5_ASAP7_75t_SL g50 ( 
.A(n_32),
.B(n_0),
.CON(n_50),
.SN(n_50)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_50),
.A2(n_0),
.B(n_1),
.Y(n_121)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_27),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_54),
.B(n_61),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_16),
.B(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_63),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_60),
.B(n_67),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_8),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_8),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_62),
.B(n_70),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_0),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_32),
.Y(n_65)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_32),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_15),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_16),
.B(n_8),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_76),
.B(n_85),
.Y(n_146)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_6),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_78),
.B(n_79),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_37),
.B(n_6),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_15),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_29),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_83),
.B(n_90),
.Y(n_139)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_37),
.Y(n_84)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_18),
.B(n_9),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_34),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_96),
.Y(n_130)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_15),
.Y(n_89)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_18),
.B(n_9),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVx2_ASAP7_75t_R g96 ( 
.A(n_42),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_63),
.A2(n_31),
.B1(n_42),
.B2(n_44),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_109),
.A2(n_150),
.B1(n_154),
.B2(n_155),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_81),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_120),
.B(n_135),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_1),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_86),
.A2(n_31),
.B1(n_44),
.B2(n_19),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_91),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_45),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_136),
.Y(n_161)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_45),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_137),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_92),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_138),
.B(n_143),
.Y(n_203)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_48),
.Y(n_141)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_88),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_73),
.Y(n_148)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_94),
.A2(n_24),
.B1(n_43),
.B2(n_26),
.Y(n_150)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_48),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_65),
.A2(n_44),
.B1(n_34),
.B2(n_24),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_79),
.A2(n_30),
.B1(n_41),
.B2(n_40),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_47),
.A2(n_30),
.B1(n_41),
.B2(n_40),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_52),
.Y(n_156)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

AO22x1_ASAP7_75t_SL g159 ( 
.A1(n_121),
.A2(n_50),
.B1(n_84),
.B2(n_95),
.Y(n_159)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_159),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_160),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_155),
.A2(n_33),
.B1(n_64),
.B2(n_74),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_163),
.A2(n_153),
.B1(n_133),
.B2(n_115),
.Y(n_222)
);

NOR2x1_ASAP7_75t_R g165 ( 
.A(n_149),
.B(n_96),
.Y(n_165)
);

OAI21x1_ASAP7_75t_SL g239 ( 
.A1(n_165),
.A2(n_167),
.B(n_189),
.Y(n_239)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_105),
.B(n_77),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_168),
.B(n_169),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_130),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_173),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_43),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_185),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_149),
.Y(n_175)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_176),
.Y(n_215)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_178),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_97),
.B(n_122),
.C(n_151),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_179),
.B(n_202),
.C(n_206),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_140),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_182),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_101),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_184),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_101),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_130),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_187),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_129),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_188),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_125),
.A2(n_93),
.B1(n_55),
.B2(n_80),
.Y(n_189)
);

CKINVDCx12_ASAP7_75t_R g190 ( 
.A(n_104),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_131),
.B(n_26),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_193),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_139),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_26),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_194),
.B(n_199),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_104),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_100),
.B(n_43),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_107),
.B(n_126),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_99),
.B(n_72),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_205),
.A2(n_98),
.B1(n_117),
.B2(n_145),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_134),
.B(n_24),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_123),
.B(n_33),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_113),
.B1(n_132),
.B2(n_110),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_209),
.B(n_195),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_187),
.A2(n_150),
.B1(n_147),
.B2(n_127),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_220),
.B1(n_222),
.B2(n_236),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_147),
.B1(n_127),
.B2(n_142),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_167),
.B(n_128),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_228),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_162),
.A2(n_118),
.B1(n_114),
.B2(n_34),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_204),
.A2(n_158),
.B1(n_102),
.B2(n_69),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_243),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_162),
.A2(n_142),
.B1(n_124),
.B2(n_116),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_164),
.A2(n_124),
.B1(n_116),
.B2(n_158),
.Y(n_237)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_204),
.A2(n_46),
.B1(n_102),
.B2(n_75),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_241),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_249),
.Y(n_276)
);

AND2x6_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_165),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_247),
.B(n_252),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_218),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_242),
.B(n_238),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_251),
.B(n_180),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_174),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_159),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_256),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_159),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_218),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_264),
.Y(n_298)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_230),
.B(n_167),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_261),
.Y(n_300)
);

CKINVDCx10_ASAP7_75t_R g262 ( 
.A(n_211),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_216),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_219),
.B(n_191),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_266),
.B(n_268),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_267),
.A2(n_273),
.B1(n_160),
.B2(n_170),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_219),
.B(n_199),
.Y(n_268)
);

INVx13_ASAP7_75t_L g269 ( 
.A(n_211),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_269),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_239),
.A2(n_164),
.B(n_181),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_270),
.A2(n_225),
.B(n_177),
.Y(n_308)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_212),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_271),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_235),
.B(n_194),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_272),
.B(n_274),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_232),
.B(n_203),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_232),
.B(n_179),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_275),
.B(n_196),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_277),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_234),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_290),
.C(n_304),
.Y(n_314)
);

OAI21xp33_ASAP7_75t_L g282 ( 
.A1(n_270),
.A2(n_221),
.B(n_240),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_261),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_235),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_285),
.B(n_305),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_253),
.A2(n_230),
.B1(n_240),
.B2(n_233),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_288),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_228),
.C(n_175),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_254),
.A2(n_239),
.B(n_189),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_292),
.A2(n_301),
.B(n_308),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_256),
.A2(n_243),
.B1(n_209),
.B2(n_228),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_293),
.A2(n_295),
.B1(n_296),
.B2(n_303),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_256),
.A2(n_228),
.B1(n_213),
.B2(n_226),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_256),
.A2(n_213),
.B1(n_215),
.B2(n_208),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_262),
.Y(n_297)
);

INVx13_ASAP7_75t_L g315 ( 
.A(n_297),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_254),
.A2(n_227),
.B(n_225),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_266),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_248),
.A2(n_166),
.B1(n_215),
.B2(n_200),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_180),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_250),
.B(n_186),
.C(n_201),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_250),
.C(n_263),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_246),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_307),
.B(n_249),
.Y(n_317)
);

AND2x6_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_247),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_309),
.B(n_327),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_310),
.B(n_331),
.Y(n_352)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_313),
.Y(n_344)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_294),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_316),
.B(n_319),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_317),
.Y(n_366)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_276),
.Y(n_318)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_318),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_294),
.B(n_252),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_321),
.B(n_300),
.C(n_261),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_297),
.Y(n_323)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_323),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_253),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_324),
.B(n_326),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_280),
.B(n_290),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_306),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_279),
.B(n_257),
.Y(n_326)
);

OA21x2_ASAP7_75t_L g327 ( 
.A1(n_289),
.A2(n_254),
.B(n_273),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_298),
.Y(n_328)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_328),
.Y(n_349)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_298),
.Y(n_329)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_329),
.Y(n_354)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_330),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_283),
.B(n_272),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_299),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_335),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_284),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_278),
.Y(n_336)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_336),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_308),
.A2(n_255),
.B(n_259),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_337),
.A2(n_338),
.B(n_301),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_289),
.A2(n_307),
.B(n_292),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_291),
.Y(n_339)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_339),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_285),
.B(n_267),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_286),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_295),
.A2(n_248),
.B1(n_268),
.B2(n_247),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_341),
.A2(n_304),
.B1(n_305),
.B2(n_287),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_261),
.Y(n_342)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_342),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_343),
.A2(n_350),
.B1(n_311),
.B2(n_332),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_345),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_311),
.A2(n_288),
.B1(n_296),
.B2(n_293),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_341),
.A2(n_289),
.B1(n_287),
.B2(n_248),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_353),
.A2(n_368),
.B1(n_332),
.B2(n_333),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_338),
.A2(n_300),
.B(n_277),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_362),
.Y(n_380)
);

XNOR2x1_ASAP7_75t_SL g360 ( 
.A(n_313),
.B(n_305),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_360),
.B(n_327),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_370),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_310),
.B(n_286),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_364),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_312),
.C(n_342),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_328),
.A2(n_248),
.B1(n_303),
.B2(n_245),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_317),
.B(n_267),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_374),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_325),
.B(n_265),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_271),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_372),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_314),
.B(n_186),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_318),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_334),
.B(n_216),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_264),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_339),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_377),
.B(n_379),
.Y(n_429)
);

AOI21xp33_ASAP7_75t_L g378 ( 
.A1(n_357),
.A2(n_329),
.B(n_337),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_378),
.A2(n_395),
.B(n_345),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_366),
.B(n_323),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_321),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_381),
.B(n_393),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_383),
.B(n_392),
.C(n_397),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_384),
.A2(n_394),
.B1(n_353),
.B2(n_349),
.Y(n_416)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_344),
.Y(n_385)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_385),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_312),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_399),
.Y(n_412)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_388),
.Y(n_417)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_344),
.Y(n_390)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_390),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_348),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_391),
.B(n_406),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_342),
.C(n_327),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_347),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_346),
.A2(n_320),
.B(n_333),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_396),
.B(n_405),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_336),
.C(n_330),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_309),
.C(n_320),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_400),
.C(n_404),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_360),
.B(n_367),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_281),
.C(n_258),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_347),
.Y(n_401)
);

INVxp33_ASAP7_75t_L g430 ( 
.A(n_401),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_351),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_402),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_373),
.B(n_281),
.C(n_216),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_352),
.B(n_315),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_365),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_365),
.B(n_315),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_361),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_392),
.B(n_346),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_408),
.B(n_422),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_376),
.B(n_359),
.C(n_348),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_411),
.B(n_415),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_413),
.A2(n_183),
.B1(n_171),
.B2(n_210),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_403),
.B(n_361),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_416),
.A2(n_423),
.B1(n_427),
.B2(n_435),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_376),
.B(n_354),
.C(n_349),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_424),
.Y(n_457)
);

BUFx5_ASAP7_75t_L g419 ( 
.A(n_381),
.Y(n_419)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_419),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_421),
.B(n_425),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_382),
.B(n_387),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_389),
.A2(n_354),
.B1(n_368),
.B2(n_356),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_382),
.B(n_358),
.C(n_356),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_398),
.B(n_358),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_386),
.A2(n_244),
.B1(n_245),
.B2(n_260),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_426),
.B(n_177),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_389),
.A2(n_260),
.B1(n_229),
.B2(n_208),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_380),
.B(n_208),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_432),
.B(n_210),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_407),
.A2(n_400),
.B1(n_404),
.B2(n_399),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_397),
.C(n_383),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_439),
.C(n_442),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_409),
.B(n_405),
.C(n_391),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_423),
.A2(n_229),
.B1(n_176),
.B2(n_172),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_441),
.A2(n_449),
.B1(n_459),
.B2(n_197),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_410),
.B(n_212),
.C(n_198),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_435),
.A2(n_188),
.B1(n_269),
.B2(n_183),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_444),
.A2(n_28),
.B1(n_17),
.B2(n_15),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_433),
.B(n_269),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_445),
.B(n_89),
.Y(n_472)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_446),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_410),
.B(n_171),
.C(n_178),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_454),
.C(n_456),
.Y(n_479)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_420),
.Y(n_448)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_448),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_434),
.A2(n_56),
.B1(n_58),
.B2(n_82),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_450),
.B(n_419),
.Y(n_467)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_451),
.Y(n_466)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_430),
.Y(n_453)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_453),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_424),
.B(n_192),
.C(n_161),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_429),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_12),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_425),
.B(n_192),
.C(n_161),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_430),
.Y(n_458)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_458),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_421),
.A2(n_417),
.B1(n_418),
.B2(n_411),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_414),
.Y(n_460)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_460),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_437),
.A2(n_433),
.B(n_408),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_463),
.A2(n_11),
.B1(n_14),
.B2(n_3),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_452),
.A2(n_431),
.B1(n_428),
.B2(n_427),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_465),
.B(n_468),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_467),
.A2(n_470),
.B1(n_475),
.B2(n_444),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_459),
.A2(n_412),
.B1(n_422),
.B2(n_173),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_440),
.B(n_412),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_443),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_471),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_472),
.B(n_28),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_436),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_474),
.B(n_477),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_438),
.B(n_28),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_439),
.A2(n_28),
.B(n_17),
.Y(n_480)
);

OAI211xp5_ASAP7_75t_L g497 ( 
.A1(n_480),
.A2(n_28),
.B(n_17),
.C(n_15),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_457),
.C(n_440),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_481),
.B(n_482),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_462),
.B(n_443),
.C(n_442),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_467),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_483),
.B(n_485),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_484),
.B(n_491),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_474),
.B(n_447),
.C(n_456),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_464),
.B(n_466),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_488),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_489),
.A2(n_494),
.B1(n_28),
.B2(n_17),
.Y(n_509)
);

NOR2xp67_ASAP7_75t_SL g490 ( 
.A(n_463),
.B(n_454),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_490),
.A2(n_497),
.B(n_498),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_469),
.B(n_445),
.C(n_441),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_478),
.B(n_460),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_492),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_473),
.B(n_449),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_495),
.B(n_461),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_496),
.B(n_17),
.Y(n_512)
);

AOI21x1_ASAP7_75t_L g498 ( 
.A1(n_476),
.A2(n_14),
.B(n_11),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_503),
.Y(n_515)
);

NOR3xp33_ASAP7_75t_L g501 ( 
.A(n_486),
.B(n_479),
.C(n_472),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_501),
.B(n_10),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_481),
.B(n_477),
.C(n_479),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_475),
.C(n_15),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_508),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_487),
.B(n_14),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_509),
.B(n_510),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_485),
.A2(n_493),
.B(n_484),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_489),
.A2(n_491),
.B(n_496),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_511),
.B(n_5),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_512),
.B(n_38),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_10),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_514),
.B(n_517),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_502),
.B(n_10),
.Y(n_517)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_518),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_499),
.B(n_14),
.Y(n_519)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_519),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_505),
.B(n_17),
.C(n_20),
.Y(n_521)
);

MAJx2_ASAP7_75t_L g529 ( 
.A(n_521),
.B(n_523),
.C(n_504),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_522),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_20),
.C(n_38),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_503),
.B(n_5),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_524),
.A2(n_500),
.B(n_501),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_507),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_526),
.B(n_20),
.Y(n_536)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_529),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_530),
.B(n_532),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_515),
.B(n_512),
.C(n_20),
.Y(n_532)
);

AOI322xp5_ASAP7_75t_L g534 ( 
.A1(n_528),
.A2(n_520),
.A3(n_519),
.B1(n_516),
.B2(n_20),
.C1(n_38),
.C2(n_9),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_534),
.A2(n_535),
.B(n_533),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_531),
.B(n_1),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_536),
.B(n_527),
.C(n_38),
.Y(n_540)
);

AO21x1_ASAP7_75t_L g542 ( 
.A1(n_539),
.A2(n_540),
.B(n_541),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_538),
.B(n_537),
.C(n_527),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_542),
.B(n_38),
.C(n_1),
.Y(n_543)
);

A2O1A1Ixp33_ASAP7_75t_L g544 ( 
.A1(n_543),
.A2(n_1),
.B(n_2),
.C(n_286),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_544),
.B(n_2),
.Y(n_545)
);


endmodule