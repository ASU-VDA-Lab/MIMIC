module real_aes_10806_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_656;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_87;
wire n_171;
wire n_676;
wire n_658;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
INVxp67_ASAP7_75t_SL g514 ( .A(n_0), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_0), .A2(n_59), .B1(n_635), .B2(n_642), .Y(n_634) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_1), .Y(n_536) );
INVx1_ASAP7_75t_L g547 ( .A(n_1), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_1), .B(n_55), .Y(n_574) );
AND2x2_ASAP7_75t_L g591 ( .A(n_1), .B(n_538), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_2), .B(n_166), .Y(n_173) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_2), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_3), .B(n_144), .Y(n_214) );
INVxp67_ASAP7_75t_L g506 ( .A(n_4), .Y(n_506) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_4), .A2(n_45), .B1(n_623), .B2(n_626), .C(n_629), .Y(n_622) );
INVxp33_ASAP7_75t_L g600 ( .A(n_5), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_5), .A2(n_30), .B1(n_654), .B2(n_656), .Y(n_653) );
OR2x2_ASAP7_75t_L g620 ( .A(n_6), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g633 ( .A(n_6), .Y(n_633) );
BUFx2_ASAP7_75t_L g539 ( .A(n_7), .Y(n_539) );
INVx1_ASAP7_75t_L g544 ( .A(n_7), .Y(n_544) );
OR2x2_ASAP7_75t_L g573 ( .A(n_7), .B(n_574), .Y(n_573) );
BUFx2_ASAP7_75t_L g695 ( .A(n_7), .Y(n_695) );
INVxp33_ASAP7_75t_L g595 ( .A(n_8), .Y(n_595) );
AOI21xp33_ASAP7_75t_L g662 ( .A1(n_8), .A2(n_663), .B(n_665), .Y(n_662) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_9), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_10), .B(n_122), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_11), .B(n_106), .Y(n_243) );
INVx1_ASAP7_75t_L g551 ( .A(n_12), .Y(n_551) );
NAND2x1p5_ASAP7_75t_L g179 ( .A(n_13), .B(n_106), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_14), .B(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g194 ( .A(n_15), .B(n_195), .Y(n_194) );
INVxp33_ASAP7_75t_L g592 ( .A(n_16), .Y(n_592) );
NAND2xp33_ASAP7_75t_SL g659 ( .A(n_16), .B(n_660), .Y(n_659) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_17), .Y(n_89) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_18), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_19), .B(n_126), .Y(n_216) );
INVx1_ASAP7_75t_L g689 ( .A(n_20), .Y(n_689) );
NAND2xp33_ASAP7_75t_L g174 ( .A(n_21), .B(n_175), .Y(n_174) );
NAND2xp33_ASAP7_75t_L g241 ( .A(n_22), .B(n_175), .Y(n_241) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_23), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_24), .Y(n_223) );
OAI221xp5_ASAP7_75t_L g565 ( .A1(n_25), .A2(n_46), .B1(n_566), .B2(n_575), .C(n_579), .Y(n_565) );
INVx1_ASAP7_75t_L g668 ( .A(n_25), .Y(n_668) );
INVx1_ASAP7_75t_L g621 ( .A(n_26), .Y(n_621) );
INVx1_ASAP7_75t_L g632 ( .A(n_26), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_27), .B(n_143), .Y(n_178) );
OAI21x1_ASAP7_75t_L g108 ( .A1(n_28), .A2(n_49), .B(n_109), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_29), .A2(n_116), .B(n_199), .C(n_201), .Y(n_198) );
INVxp33_ASAP7_75t_L g586 ( .A(n_30), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_31), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_32), .B(n_120), .Y(n_137) );
NAND2xp33_ASAP7_75t_L g167 ( .A(n_33), .B(n_161), .Y(n_167) );
AND2x6_ASAP7_75t_L g83 ( .A(n_34), .B(n_84), .Y(n_83) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_34), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_34), .B(n_701), .Y(n_748) );
INVx1_ASAP7_75t_L g555 ( .A(n_35), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_36), .B(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_37), .B(n_200), .Y(n_240) );
NAND2xp33_ASAP7_75t_L g215 ( .A(n_38), .B(n_161), .Y(n_215) );
INVx1_ASAP7_75t_L g84 ( .A(n_39), .Y(n_84) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_39), .Y(n_701) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_40), .Y(n_231) );
INVx1_ASAP7_75t_L g560 ( .A(n_41), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_42), .B(n_161), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_43), .Y(n_135) );
AND2x2_ASAP7_75t_L g203 ( .A(n_44), .B(n_126), .Y(n_203) );
INVxp33_ASAP7_75t_L g527 ( .A(n_45), .Y(n_527) );
INVx1_ASAP7_75t_L g676 ( .A(n_46), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_47), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g513 ( .A(n_48), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_50), .Y(n_177) );
NAND2xp33_ASAP7_75t_L g112 ( .A(n_51), .B(n_92), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_52), .B(n_166), .Y(n_165) );
BUFx10_ASAP7_75t_L g717 ( .A(n_53), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_54), .B(n_91), .Y(n_238) );
INVx2_ASAP7_75t_L g538 ( .A(n_55), .Y(n_538) );
NAND2xp33_ASAP7_75t_L g121 ( .A(n_56), .B(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_57), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_58), .B(n_175), .Y(n_237) );
INVxp33_ASAP7_75t_L g521 ( .A(n_59), .Y(n_521) );
INVx1_ASAP7_75t_L g732 ( .A(n_60), .Y(n_732) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_61), .Y(n_202) );
INVx2_ASAP7_75t_L g109 ( .A(n_62), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_63), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_64), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_65), .B(n_147), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_66), .Y(n_210) );
INVx1_ASAP7_75t_L g193 ( .A(n_67), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_68), .Y(n_225) );
AND2x2_ASAP7_75t_L g233 ( .A(n_69), .B(n_106), .Y(n_233) );
INVx1_ASAP7_75t_L g564 ( .A(n_70), .Y(n_564) );
INVx2_ASAP7_75t_L g512 ( .A(n_71), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g722 ( .A(n_72), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_73), .B(n_126), .Y(n_125) );
BUFx3_ASAP7_75t_L g617 ( .A(n_74), .Y(n_617) );
INVx1_ASAP7_75t_L g645 ( .A(n_74), .Y(n_645) );
BUFx3_ASAP7_75t_L g618 ( .A(n_75), .Y(n_618) );
INVx1_ASAP7_75t_L g625 ( .A(n_75), .Y(n_625) );
XNOR2xp5_ASAP7_75t_L g499 ( .A(n_76), .B(n_500), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_94), .B(n_498), .Y(n_77) );
BUFx2_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
AND2x2_ASAP7_75t_L g79 ( .A(n_80), .B(n_85), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx8_ASAP7_75t_L g124 ( .A(n_82), .Y(n_124) );
NOR2xp67_ASAP7_75t_L g185 ( .A(n_82), .B(n_186), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_82), .A2(n_221), .B(n_227), .Y(n_220) );
INVx8_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
BUFx2_ASAP7_75t_L g168 ( .A(n_83), .Y(n_168) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_86), .Y(n_85) );
AO21x1_ASAP7_75t_L g746 ( .A1(n_86), .A2(n_747), .B(n_748), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g86 ( .A(n_87), .B(n_90), .Y(n_86) );
OAI21x1_ASAP7_75t_L g189 ( .A1(n_87), .A2(n_190), .B(n_194), .Y(n_189) );
BUFx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx3_ASAP7_75t_L g145 ( .A(n_88), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_88), .A2(n_165), .B(n_167), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_88), .Y(n_232) );
BUFx12f_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx5_ASAP7_75t_L g116 ( .A(n_89), .Y(n_116) );
INVx5_ASAP7_75t_L g123 ( .A(n_89), .Y(n_123) );
O2A1O1Ixp33_ASAP7_75t_L g134 ( .A1(n_89), .A2(n_135), .B(n_136), .C(n_137), .Y(n_134) );
HB1xp67_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g136 ( .A(n_91), .Y(n_136) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx2_ASAP7_75t_L g114 ( .A(n_92), .Y(n_114) );
INVx2_ASAP7_75t_L g163 ( .A(n_92), .Y(n_163) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_93), .Y(n_120) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_93), .Y(n_122) );
INVx2_ASAP7_75t_L g144 ( .A(n_93), .Y(n_144) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_93), .Y(n_192) );
INVx1_ASAP7_75t_L g197 ( .A(n_93), .Y(n_197) );
INVx2_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
NAND3x1_ASAP7_75t_L g96 ( .A(n_97), .B(n_361), .C(n_441), .Y(n_96) );
NOR4xp75_ASAP7_75t_L g97 ( .A(n_98), .B(n_282), .C(n_311), .D(n_337), .Y(n_97) );
NAND3x1_ASAP7_75t_L g98 ( .A(n_99), .B(n_244), .C(n_266), .Y(n_98) );
OAI21xp5_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_149), .B(n_180), .Y(n_99) );
INVxp33_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_102), .B(n_128), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_104), .B(n_271), .Y(n_301) );
OR2x2_ASAP7_75t_L g383 ( .A(n_104), .B(n_263), .Y(n_383) );
INVx2_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g258 ( .A(n_105), .Y(n_258) );
INVx1_ASAP7_75t_SL g343 ( .A(n_105), .Y(n_343) );
BUFx2_ASAP7_75t_L g408 ( .A(n_105), .Y(n_408) );
OA21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_110), .B(n_125), .Y(n_105) );
BUFx4f_ASAP7_75t_L g132 ( .A(n_106), .Y(n_132) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_106), .A2(n_110), .B(n_125), .Y(n_151) );
INVx3_ASAP7_75t_L g157 ( .A(n_106), .Y(n_157) );
INVx4_ASAP7_75t_L g187 ( .A(n_106), .Y(n_187) );
OA21x2_ASAP7_75t_L g317 ( .A1(n_106), .A2(n_110), .B(n_125), .Y(n_317) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g148 ( .A(n_107), .Y(n_148) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g127 ( .A(n_108), .Y(n_127) );
OAI21x1_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_117), .B(n_124), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_113), .B(n_115), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_115), .A2(n_173), .B(n_174), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_115), .A2(n_214), .B(n_215), .Y(n_213) );
CKINVDCx6p67_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g226 ( .A(n_116), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_121), .B(n_123), .Y(n_117) );
NOR2xp67_ASAP7_75t_L g224 ( .A(n_119), .B(n_225), .Y(n_224) );
INVx5_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g141 ( .A(n_122), .Y(n_141) );
INVx2_ASAP7_75t_L g166 ( .A(n_122), .Y(n_166) );
INVx2_ASAP7_75t_SL g200 ( .A(n_122), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_122), .B(n_223), .Y(n_222) );
AOI21x1_ASAP7_75t_L g159 ( .A1(n_123), .A2(n_160), .B(n_162), .Y(n_159) );
INVx1_ASAP7_75t_L g242 ( .A(n_123), .Y(n_242) );
OAI21x1_ASAP7_75t_L g133 ( .A1(n_124), .A2(n_134), .B(n_138), .Y(n_133) );
OAI21x1_ASAP7_75t_L g171 ( .A1(n_124), .A2(n_172), .B(n_176), .Y(n_171) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_124), .A2(n_209), .B(n_213), .Y(n_208) );
OAI21x1_ASAP7_75t_L g235 ( .A1(n_124), .A2(n_236), .B(n_239), .Y(n_235) );
BUFx5_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g396 ( .A(n_128), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_SL g360 ( .A(n_129), .B(n_326), .Y(n_360) );
NAND2xp33_ASAP7_75t_R g492 ( .A(n_129), .B(n_326), .Y(n_492) );
BUFx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_130), .B(n_317), .Y(n_323) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g310 ( .A(n_131), .B(n_272), .Y(n_310) );
OR2x2_ASAP7_75t_L g381 ( .A(n_131), .B(n_154), .Y(n_381) );
AND2x2_ASAP7_75t_L g430 ( .A(n_131), .B(n_263), .Y(n_430) );
OAI21x1_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B(n_146), .Y(n_131) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_132), .A2(n_171), .B(n_179), .Y(n_170) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_132), .A2(n_208), .B(n_216), .Y(n_207) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_132), .A2(n_133), .B(n_146), .Y(n_261) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_132), .A2(n_171), .B(n_179), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .B(n_142), .C(n_145), .Y(n_138) );
O2A1O1Ixp5_ASAP7_75t_L g176 ( .A1(n_140), .A2(n_145), .B(n_177), .C(n_178), .Y(n_176) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g161 ( .A(n_144), .Y(n_161) );
INVx2_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
O2A1O1Ixp5_ASAP7_75t_L g209 ( .A1(n_145), .A2(n_210), .B(n_211), .C(n_212), .Y(n_209) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_149), .A2(n_432), .B1(n_437), .B2(n_439), .Y(n_431) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
AOI32xp33_ASAP7_75t_L g425 ( .A1(n_150), .A2(n_309), .A3(n_349), .B1(n_426), .B2(n_427), .Y(n_425) );
OAI322xp33_ASAP7_75t_L g442 ( .A1(n_150), .A2(n_443), .A3(n_444), .B1(n_445), .B2(n_448), .C1(n_451), .C2(n_453), .Y(n_442) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g270 ( .A(n_151), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g495 ( .A(n_151), .Y(n_495) );
INVx2_ASAP7_75t_L g397 ( .A(n_152), .Y(n_397) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_170), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_153), .B(n_263), .Y(n_304) );
INVx2_ASAP7_75t_L g375 ( .A(n_153), .Y(n_375) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g274 ( .A(n_154), .B(n_264), .Y(n_274) );
AND2x2_ASAP7_75t_L g326 ( .A(n_154), .B(n_265), .Y(n_326) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OAI21x1_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_158), .B(n_169), .Y(n_155) );
OAI21x1_ASAP7_75t_L g234 ( .A1(n_156), .A2(n_235), .B(n_243), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_156), .A2(n_158), .B(n_169), .Y(n_272) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_164), .B(n_168), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_161), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g211 ( .A(n_163), .Y(n_211) );
INVx2_ASAP7_75t_L g300 ( .A(n_170), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_175), .B(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g744 ( .A(n_177), .Y(n_744) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_204), .Y(n_180) );
INVx2_ASAP7_75t_L g320 ( .A(n_181), .Y(n_320) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g252 ( .A(n_182), .B(n_219), .Y(n_252) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g289 ( .A(n_183), .B(n_219), .Y(n_289) );
AND2x2_ASAP7_75t_L g292 ( .A(n_183), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g329 ( .A(n_183), .Y(n_329) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g250 ( .A(n_184), .Y(n_250) );
AOI21x1_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_188), .B(n_203), .Y(n_184) );
INVx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_187), .A2(n_220), .B(n_233), .Y(n_219) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_187), .A2(n_220), .B(n_233), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_198), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_193), .Y(n_190) );
NOR2xp33_ASAP7_75t_SL g230 ( .A(n_191), .B(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx3_ASAP7_75t_L g477 ( .A(n_204), .Y(n_477) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_217), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_206), .B(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g254 ( .A(n_206), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_206), .B(n_250), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_206), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_206), .B(n_217), .Y(n_359) );
AND2x2_ASAP7_75t_L g436 ( .A(n_206), .B(n_416), .Y(n_436) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g297 ( .A(n_207), .Y(n_297) );
AND2x2_ASAP7_75t_L g330 ( .A(n_207), .B(n_219), .Y(n_330) );
AND2x2_ASAP7_75t_L g267 ( .A(n_217), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVxp67_ASAP7_75t_SL g246 ( .A(n_218), .Y(n_246) );
OR2x2_ASAP7_75t_L g306 ( .A(n_218), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_234), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_224), .B(n_226), .Y(n_221) );
OAI21xp33_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_230), .B(n_232), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_229), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_229), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_232), .A2(n_237), .B(n_238), .Y(n_236) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_234), .Y(n_255) );
INVx1_ASAP7_75t_L g281 ( .A(n_234), .Y(n_281) );
INVx1_ASAP7_75t_L g296 ( .A(n_234), .Y(n_296) );
AND2x2_ASAP7_75t_L g328 ( .A(n_234), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g401 ( .A(n_234), .B(n_297), .Y(n_401) );
INVx1_ASAP7_75t_L g416 ( .A(n_234), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_242), .Y(n_239) );
OAI21xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_251), .B(n_256), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_249), .B(n_386), .Y(n_440) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g307 ( .A(n_250), .Y(n_307) );
INVxp67_ASAP7_75t_SL g450 ( .A(n_250), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_251), .A2(n_303), .B1(n_305), .B2(n_308), .Y(n_302) );
AND2x4_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g340 ( .A(n_252), .Y(n_340) );
AND2x2_ASAP7_75t_L g426 ( .A(n_252), .B(n_393), .Y(n_426) );
NAND2xp67_ASAP7_75t_L g497 ( .A(n_252), .B(n_401), .Y(n_497) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g470 ( .A(n_254), .Y(n_470) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
OR2x2_ASAP7_75t_L g333 ( .A(n_258), .B(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g457 ( .A(n_258), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_259), .B(n_423), .Y(n_422) );
NAND2x1_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
INVx1_ASAP7_75t_L g276 ( .A(n_260), .Y(n_276) );
AND2x4_ASAP7_75t_SL g374 ( .A(n_260), .B(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g444 ( .A(n_260), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_260), .B(n_300), .Y(n_458) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g347 ( .A(n_261), .Y(n_347) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_261), .Y(n_390) );
INVx1_ASAP7_75t_L g476 ( .A(n_262), .Y(n_476) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g373 ( .A(n_263), .B(n_317), .Y(n_373) );
AND2x2_ASAP7_75t_L g419 ( .A(n_263), .B(n_317), .Y(n_419) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_270), .B1(n_273), .B2(n_277), .Y(n_266) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_268), .Y(n_479) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g278 ( .A(n_269), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g423 ( .A(n_271), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_271), .B(n_355), .Y(n_462) );
BUFx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g334 ( .A(n_274), .Y(n_334) );
AND2x4_ASAP7_75t_L g345 ( .A(n_274), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g406 ( .A(n_274), .B(n_407), .Y(n_406) );
O2A1O1Ixp5_ASAP7_75t_L g475 ( .A1(n_275), .A2(n_333), .B(n_476), .C(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_278), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx2_ASAP7_75t_SL g293 ( .A(n_280), .Y(n_293) );
INVx1_ASAP7_75t_L g352 ( .A(n_280), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_280), .B(n_297), .Y(n_386) );
INVx1_ASAP7_75t_L g288 ( .A(n_281), .Y(n_288) );
OAI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_298), .B(n_302), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2x1_ASAP7_75t_SL g284 ( .A(n_285), .B(n_290), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_287), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g488 ( .A(n_288), .B(n_292), .Y(n_488) );
AND2x2_ASAP7_75t_L g335 ( .A(n_289), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g377 ( .A(n_289), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_289), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_289), .B(n_394), .Y(n_405) );
AND2x2_ASAP7_75t_L g420 ( .A(n_289), .B(n_401), .Y(n_420) );
OAI221xp5_ASAP7_75t_L g454 ( .A1(n_290), .A2(n_306), .B1(n_455), .B2(n_457), .C(n_459), .Y(n_454) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
AND2x4_ASAP7_75t_L g400 ( .A(n_292), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g452 ( .A(n_292), .B(n_394), .Y(n_452) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_293), .Y(n_368) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g336 ( .A(n_295), .Y(n_336) );
INVx1_ASAP7_75t_L g369 ( .A(n_295), .Y(n_369) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
BUFx3_ASAP7_75t_L g394 ( .A(n_297), .Y(n_394) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
AND2x2_ASAP7_75t_L g308 ( .A(n_299), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_300), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_303), .B(n_322), .Y(n_438) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g403 ( .A(n_304), .B(n_390), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_305), .A2(n_402), .B1(n_491), .B2(n_496), .Y(n_490) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g434 ( .A(n_307), .Y(n_434) );
AND2x2_ASAP7_75t_L g446 ( .A(n_309), .B(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_310), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g357 ( .A(n_310), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_331), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_318), .B1(n_321), .B2(n_327), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g474 ( .A(n_315), .Y(n_474) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVxp67_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVxp67_ASAP7_75t_L g410 ( .A(n_322), .Y(n_410) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g428 ( .A(n_324), .Y(n_428) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g485 ( .A(n_326), .B(n_346), .Y(n_485) );
AND2x2_ASAP7_75t_L g489 ( .A(n_326), .B(n_408), .Y(n_489) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx1_ASAP7_75t_L g353 ( .A(n_328), .Y(n_353) );
AND2x2_ASAP7_75t_L g482 ( .A(n_328), .B(n_352), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_335), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI32xp33_ASAP7_75t_L g417 ( .A1(n_335), .A2(n_418), .A3(n_419), .B1(n_420), .B2(n_421), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_341), .B(n_348), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NOR2x1p5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g355 ( .A(n_343), .Y(n_355) );
INVx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g473 ( .A(n_346), .Y(n_473) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_354), .B1(n_358), .B2(n_360), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_351), .Y(n_411) );
INVx1_ASAP7_75t_L g471 ( .A(n_352), .Y(n_471) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NOR3xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_398), .C(n_424), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_363), .B(n_384), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_370), .B1(n_376), .B2(n_378), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_369), .Y(n_365) );
INVxp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g465 ( .A(n_367), .Y(n_465) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
AND2x4_ASAP7_75t_L g460 ( .A(n_372), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g447 ( .A(n_373), .Y(n_447) );
INVx2_ASAP7_75t_L g418 ( .A(n_374), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_374), .B(n_494), .Y(n_493) );
BUFx2_ASAP7_75t_L g413 ( .A(n_375), .Y(n_413) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2x1_ASAP7_75t_SL g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g388 ( .A(n_383), .B(n_389), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .B1(n_391), .B2(n_395), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVxp67_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_390), .Y(n_461) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g494 ( .A(n_394), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_417), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_402), .B1(n_404), .B2(n_406), .C(n_409), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_401), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g464 ( .A(n_401), .Y(n_464) );
INVx2_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NOR4xp25_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .C(n_412), .D(n_414), .Y(n_409) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g443 ( .A(n_415), .B(n_440), .Y(n_443) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g453 ( .A(n_419), .Y(n_453) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_431), .Y(n_424) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NOR3xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_454), .C(n_466), .Y(n_441) );
AND2x2_ASAP7_75t_L g456 ( .A(n_444), .B(n_447), .Y(n_456) );
INVxp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI21xp33_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_462), .B(n_463), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
NAND3xp33_ASAP7_75t_SL g466 ( .A(n_467), .B(n_478), .C(n_490), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_472), .B(n_475), .Y(n_467) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_470), .B(n_471), .Y(n_469) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
O2A1O1Ixp5_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_480), .B(n_483), .C(n_486), .Y(n_478) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2x1p5_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
OAI221xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B1(n_697), .B2(n_704), .C(n_741), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_500), .A2(n_742), .B1(n_744), .B2(n_745), .Y(n_741) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_606), .Y(n_502) );
NOR3xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_565), .C(n_584), .Y(n_503) );
OAI33xp33_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_520), .A3(n_534), .B1(n_540), .B2(n_548), .B3(n_556), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B1(n_514), .B2(n_515), .Y(n_505) );
BUFx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g559 ( .A(n_510), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_513), .Y(n_510) );
INVx1_ASAP7_75t_L g578 ( .A(n_511), .Y(n_578) );
AND2x4_ASAP7_75t_L g603 ( .A(n_511), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x4_ASAP7_75t_L g518 ( .A(n_512), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_512), .B(n_513), .Y(n_526) );
INVx1_ASAP7_75t_L g533 ( .A(n_512), .Y(n_533) );
INVx1_ASAP7_75t_L g583 ( .A(n_512), .Y(n_583) );
AND2x2_ASAP7_75t_L g599 ( .A(n_512), .B(n_513), .Y(n_599) );
INVx2_ASAP7_75t_L g519 ( .A(n_513), .Y(n_519) );
INVx1_ASAP7_75t_L g532 ( .A(n_513), .Y(n_532) );
INVx1_ASAP7_75t_L g571 ( .A(n_513), .Y(n_571) );
INVx1_ASAP7_75t_L g605 ( .A(n_513), .Y(n_605) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx3_ASAP7_75t_L g589 ( .A(n_517), .Y(n_589) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_518), .Y(n_563) );
AND2x4_ASAP7_75t_L g582 ( .A(n_519), .B(n_583), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B1(n_527), .B2(n_528), .Y(n_520) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g550 ( .A(n_524), .Y(n_550) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g692 ( .A(n_525), .B(n_573), .Y(n_692) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
AND2x2_ASAP7_75t_L g554 ( .A(n_532), .B(n_533), .Y(n_554) );
OR2x6_ASAP7_75t_L g534 ( .A(n_535), .B(n_539), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g546 ( .A(n_538), .Y(n_546) );
BUFx2_ASAP7_75t_L g609 ( .A(n_539), .Y(n_609) );
CKINVDCx8_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
INVx5_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OR2x6_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x4_ASAP7_75t_L g590 ( .A(n_544), .B(n_591), .Y(n_590) );
NAND2x1p5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
OAI22xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_551), .B1(n_552), .B2(n_555), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_551), .A2(n_560), .B1(n_678), .B2(n_683), .Y(n_677) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_555), .A2(n_612), .B1(n_622), .B2(n_634), .C(n_646), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_560), .B1(n_561), .B2(n_564), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_564), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2x1_ASAP7_75t_SL g568 ( .A(n_569), .B(n_572), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2x1p5_ASAP7_75t_L g576 ( .A(n_572), .B(n_577), .Y(n_576) );
NAND2x1p5_ASAP7_75t_L g580 ( .A(n_572), .B(n_581), .Y(n_580) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx4f_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
BUFx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x6_ASAP7_75t_L g593 ( .A(n_581), .B(n_590), .Y(n_593) );
BUFx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_594), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B1(n_592), .B2(n_593), .Y(n_585) );
BUFx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x4_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
AND2x4_ASAP7_75t_L g596 ( .A(n_590), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g601 ( .A(n_590), .B(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_600), .B2(n_601), .Y(n_594) );
INVx2_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
INVx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_610), .B1(n_689), .B2(n_690), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND4xp25_ASAP7_75t_L g610 ( .A(n_611), .B(n_652), .C(n_677), .D(n_685), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_615), .B(n_619), .Y(n_614) );
INVx2_ASAP7_75t_SL g661 ( .A(n_615), .Y(n_661) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_616), .Y(n_628) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
AND2x4_ASAP7_75t_L g624 ( .A(n_617), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g640 ( .A(n_617), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_618), .Y(n_641) );
AND2x4_ASAP7_75t_L g644 ( .A(n_618), .B(n_645), .Y(n_644) );
AND2x4_ASAP7_75t_L g683 ( .A(n_619), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g679 ( .A(n_620), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g687 ( .A(n_620), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g650 ( .A(n_621), .Y(n_650) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_SL g655 ( .A(n_624), .Y(n_655) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_624), .Y(n_684) );
INVx1_ASAP7_75t_L g682 ( .A(n_625), .Y(n_682) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x4_ASAP7_75t_L g646 ( .A(n_627), .B(n_647), .Y(n_646) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx3_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
BUFx3_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_SL g712 ( .A(n_631), .Y(n_712) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
AND2x4_ASAP7_75t_L g667 ( .A(n_632), .B(n_651), .Y(n_667) );
INVx2_ASAP7_75t_L g651 ( .A(n_633), .Y(n_651) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g664 ( .A(n_638), .Y(n_664) );
INVx6_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g696 ( .A(n_639), .B(n_649), .Y(n_696) );
AND2x4_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g675 ( .A(n_640), .Y(n_675) );
INVx1_ASAP7_75t_L g672 ( .A(n_641), .Y(n_672) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_644), .Y(n_658) );
INVx2_ASAP7_75t_L g688 ( .A(n_644), .Y(n_688) );
INVx1_ASAP7_75t_L g681 ( .A(n_645), .Y(n_681) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x4_ASAP7_75t_L g669 ( .A(n_649), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g673 ( .A(n_649), .B(n_674), .Y(n_673) );
AND2x4_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
AOI322xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_659), .A3(n_662), .B1(n_668), .B2(n_669), .C1(n_673), .C2(n_676), .Y(n_652) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
BUFx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx2_ASAP7_75t_SL g719 ( .A(n_669), .Y(n_719) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g715 ( .A(n_671), .Y(n_715) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
BUFx3_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx6_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx4_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx5_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x4_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x4_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
BUFx3_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
CKINVDCx5p33_ASAP7_75t_R g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_701), .B(n_703), .Y(n_708) );
INVx1_ASAP7_75t_SL g747 ( .A(n_701), .Y(n_747) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_720), .B1(n_736), .B2(n_740), .Y(n_704) );
BUFx12f_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
CKINVDCx20_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
BUFx6f_ASAP7_75t_L g743 ( .A(n_707), .Y(n_743) );
OR2x6_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
OR2x4_ASAP7_75t_L g739 ( .A(n_708), .B(n_710), .Y(n_739) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI31xp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_713), .A3(n_716), .B(n_718), .Y(n_710) );
BUFx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx6_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_720), .A2(n_739), .B1(n_740), .B2(n_743), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_726), .B1(n_734), .B2(n_735), .Y(n_720) );
CKINVDCx16_ASAP7_75t_R g734 ( .A(n_721), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_721) );
INVx1_ASAP7_75t_L g724 ( .A(n_722), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_723), .Y(n_725) );
INVx1_ASAP7_75t_L g735 ( .A(n_726), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
CKINVDCx14_ASAP7_75t_R g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx8_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
BUFx2_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
endmodule