module fake_jpeg_21764_n_73 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_6),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_4),
.B(n_7),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_18),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_12),
.B1(n_11),
.B2(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_21),
.B(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_15),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_19),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_29),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_34),
.B(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_32),
.Y(n_35)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_17),
.B1(n_24),
.B2(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2x1_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_32),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_29),
.A2(n_8),
.B1(n_14),
.B2(n_9),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_30),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_18),
.C(n_20),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_50),
.C(n_39),
.Y(n_52)
);

NOR4xp25_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_10),
.C(n_9),
.D(n_20),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_35),
.C(n_43),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_16),
.C(n_11),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_56),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_54),
.B(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_40),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_57),
.A2(n_59),
.B(n_60),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_42),
.B1(n_35),
.B2(n_38),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_52),
.B1(n_11),
.B2(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_16),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_0),
.C(n_1),
.Y(n_65)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_63),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_65),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_1),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_SL g70 ( 
.A1(n_67),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_61),
.B1(n_67),
.B2(n_3),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_69),
.A2(n_70),
.B(n_4),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_5),
.C(n_6),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_5),
.C(n_7),
.Y(n_73)
);


endmodule