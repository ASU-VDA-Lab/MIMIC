module fake_jpeg_23832_n_43 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_0),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_5),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_1),
.B(n_4),
.Y(n_15)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_2),
.C(n_3),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_18),
.C(n_23),
.Y(n_26)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_19),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_3),
.B(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_14),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_15),
.Y(n_20)
);

HAxp5_ASAP7_75t_SL g29 ( 
.A(n_20),
.B(n_21),
.CON(n_29),
.SN(n_29)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_8),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_7),
.B(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_24),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_16),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_28),
.Y(n_38)
);

AND2x4_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_13),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_26),
.B(n_32),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_33),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_12),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_37),
.A2(n_38),
.B(n_28),
.Y(n_39)
);

NAND4xp25_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_28),
.C(n_37),
.D(n_29),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_40),
.B1(n_29),
.B2(n_34),
.Y(n_42)
);

BUFx24_ASAP7_75t_SL g43 ( 
.A(n_42),
.Y(n_43)
);


endmodule