module fake_jpeg_26625_n_173 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVxp33_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_33),
.Y(n_38)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_23),
.B(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_25),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_29),
.C(n_35),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_14),
.C(n_20),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_17),
.B1(n_28),
.B2(n_33),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_45),
.B1(n_34),
.B2(n_33),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_46),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_31),
.A2(n_28),
.B1(n_14),
.B2(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_16),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_32),
.Y(n_53)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_60),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_31),
.B1(n_37),
.B2(n_28),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_16),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_19),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_61),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_26),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_63),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_72),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_47),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_30),
.B1(n_34),
.B2(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_48),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_82),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_36),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_70),
.B(n_22),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_87),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_63),
.A2(n_27),
.B(n_20),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_27),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_41),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_36),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_24),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_100),
.Y(n_118)
);

OA21x2_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_71),
.B(n_68),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_101),
.B(n_106),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_59),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_102),
.B(n_103),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_24),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_77),
.Y(n_104)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_22),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_109),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_71),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

AOI22x1_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_36),
.B1(n_30),
.B2(n_43),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_91),
.B1(n_80),
.B2(n_62),
.Y(n_115)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_114),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_85),
.A3(n_94),
.B1(n_89),
.B2(n_78),
.C1(n_111),
.C2(n_73),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_113),
.B1(n_121),
.B2(n_119),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_78),
.C(n_81),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_121),
.C(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_78),
.Y(n_119)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_85),
.C(n_75),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_125),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_83),
.C(n_92),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_75),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_30),
.Y(n_139)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_106),
.B(n_80),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_133),
.B(n_134),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_139),
.C(n_117),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_115),
.A2(n_98),
.B1(n_101),
.B2(n_91),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_132),
.B(n_140),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_95),
.B(n_98),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_52),
.B1(n_90),
.B2(n_65),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_100),
.Y(n_143)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_138),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_2),
.B(n_3),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_135),
.C(n_25),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

AOI321xp33_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_127),
.A3(n_112),
.B1(n_123),
.B2(n_124),
.C(n_116),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_146),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_41),
.C(n_60),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_13),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_149),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_15),
.C(n_25),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_140),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_150),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_148),
.A2(n_141),
.B(n_145),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_152),
.A2(n_153),
.B(n_2),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_148),
.A2(n_138),
.B1(n_128),
.B2(n_132),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_2),
.C(n_3),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_151),
.A2(n_11),
.B1(n_9),
.B2(n_15),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_158),
.B(n_159),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_11),
.B(n_9),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_163),
.C(n_156),
.Y(n_164)
);

AOI211xp5_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_162),
.B(n_6),
.C(n_7),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_154),
.A2(n_4),
.B(n_5),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_5),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_164),
.B(n_165),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_157),
.C(n_6),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_6),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_168),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_172),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);


endmodule