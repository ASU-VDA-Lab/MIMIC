module fake_ibex_911_n_4401 (n_151, n_85, n_599, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_421, n_738, n_475, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_768, n_338, n_173, n_696, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_762, n_410, n_308, n_675, n_463, n_624, n_706, n_411, n_135, n_520, n_684, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_744, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_728, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_752, n_668, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_232, n_380, n_749, n_281, n_559, n_425, n_4401);

input n_151;
input n_85;
input n_599;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_421;
input n_738;
input n_475;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_768;
input n_338;
input n_173;
input n_696;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_684;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_744;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_752;
input n_668;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4401;

wire n_1084;
wire n_4368;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_845;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4204;
wire n_4364;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_773;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3272;
wire n_3255;
wire n_3674;
wire n_4249;
wire n_1652;
wire n_969;
wire n_1954;
wire n_1859;
wire n_2183;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_4372;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_4353;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_4343;
wire n_1722;
wire n_4371;
wire n_3931;
wire n_911;
wire n_2023;
wire n_781;
wire n_2720;
wire n_3870;
wire n_4179;
wire n_802;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_4360;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_1782;
wire n_963;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_4399;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_4378;
wire n_850;
wire n_4169;
wire n_3175;
wire n_3729;
wire n_4239;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4172;
wire n_1730;
wire n_4277;
wire n_1307;
wire n_875;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_3982;
wire n_2605;
wire n_2343;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_4285;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3896;
wire n_3753;
wire n_3533;
wire n_2192;
wire n_1766;
wire n_3566;
wire n_3184;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_824;
wire n_4304;
wire n_4348;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4160;
wire n_4382;
wire n_787;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_3969;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_4311;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_852;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3884;
wire n_3949;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2436;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_1841;
wire n_1070;
wire n_2472;
wire n_4389;
wire n_777;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3699;
wire n_1955;
wire n_3668;
wire n_4312;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_3973;
wire n_1313;
wire n_4214;
wire n_4223;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_4295;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_3858;
wire n_772;
wire n_4182;
wire n_810;
wire n_1401;
wire n_3764;
wire n_4173;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_4259;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_4188;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_784;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_1326;
wire n_971;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_4393;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_4283;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_4392;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_4352;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_4258;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_4290;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_4252;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2625;
wire n_2444;
wire n_1742;
wire n_2350;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3887;
wire n_3963;
wire n_3800;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4103;
wire n_3583;
wire n_2019;
wire n_4126;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_4400;
wire n_2499;
wire n_3370;
wire n_4359;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_4331;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_819;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_4098;
wire n_3471;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_4156;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_4355;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_4308;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_3054;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_4293;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_4253;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4122;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_4374;
wire n_1140;
wire n_1985;
wire n_4375;
wire n_4205;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_2573;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_2423;
wire n_4230;
wire n_859;
wire n_3849;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_4333;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_4330;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_3813;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_4033;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_3364;
wire n_1236;
wire n_4384;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4323;
wire n_4184;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_4325;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_4337;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_4292;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_4362;
wire n_3568;
wire n_944;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_3331;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_2999;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_4347;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_4307;
wire n_3526;
wire n_2102;
wire n_4356;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_4151;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_2991;
wire n_847;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_4365;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_4215;
wire n_4315;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3797;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3584;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_4379;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_882;
wire n_4157;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_814;
wire n_3829;
wire n_1864;
wire n_943;
wire n_4317;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_4297;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_803;
wire n_2570;
wire n_4051;
wire n_4321;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1599;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_3070;
wire n_2842;
wire n_3646;
wire n_2635;
wire n_3477;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_817;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_4255;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_4361;
wire n_3974;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_3495;
wire n_863;
wire n_2185;
wire n_4141;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2979;
wire n_2376;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_4291;
wire n_3419;
wire n_3629;
wire n_807;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_4117;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_3735;
wire n_4154;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_4318;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_4385;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4195;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_3925;
wire n_4089;
wire n_4176;
wire n_1683;
wire n_1185;
wire n_4256;
wire n_3575;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_4278;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_4322;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_1004;
wire n_947;
wire n_4276;
wire n_831;
wire n_3929;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2684;
wire n_2875;
wire n_3284;
wire n_2524;
wire n_3835;
wire n_1437;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_3927;
wire n_2422;
wire n_4185;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_4381;
wire n_1917;
wire n_4314;
wire n_1444;
wire n_4133;
wire n_920;
wire n_4316;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_4306;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_991;
wire n_1331;
wire n_1223;
wire n_961;
wire n_2127;
wire n_3747;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_4388;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_4138;
wire n_4121;
wire n_3552;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_4142;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4118;
wire n_4183;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_4284;
wire n_1458;
wire n_1694;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3673;
wire n_3476;
wire n_4066;
wire n_3990;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1850;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_4123;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2683;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_4305;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_4339;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_3878;
wire n_4016;
wire n_798;
wire n_2849;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_4286;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_785;
wire n_2180;
wire n_1952;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_4289;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3912;
wire n_3778;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1348;
wire n_1289;
wire n_838;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_4099;
wire n_4377;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_4264;
wire n_789;
wire n_1942;
wire n_4326;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2698;
wire n_2274;
wire n_1617;
wire n_1839;
wire n_3899;
wire n_4149;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_3930;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_4319;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_4383;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_3745;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_4287;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_4300;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_4022;
wire n_4212;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_4320;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_4357;
wire n_3096;
wire n_3333;
wire n_839;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_4366;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_1238;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_4139;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_4288;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_4340;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2447;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_3784;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_775;
wire n_3273;
wire n_4367;
wire n_950;
wire n_2700;
wire n_3139;
wire n_1222;
wire n_4282;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3928;
wire n_3619;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_4334;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_4338;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_833;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_1513;
wire n_3740;
wire n_4397;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_4344;
wire n_2366;
wire n_4229;
wire n_4294;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_4351;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4111;
wire n_4162;
wire n_4200;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_4341;
wire n_4328;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_792;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_3059;
wire n_2567;
wire n_3085;
wire n_1242;
wire n_2867;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_4189;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_4390;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_794;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_4058;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4148;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3576;
wire n_3109;
wire n_1961;
wire n_3491;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_4265;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2864;
wire n_2406;
wire n_1632;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4017;
wire n_1547;
wire n_946;
wire n_1542;
wire n_1362;
wire n_1586;
wire n_3497;
wire n_4178;
wire n_4324;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4313;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3586;
wire n_956;
wire n_3561;
wire n_790;
wire n_4125;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_2574;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_4242;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_4279;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_4235;
wire n_1438;
wire n_3972;
wire n_3774;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_4350;
wire n_4380;
wire n_1361;
wire n_1187;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_3102;
wire n_2872;
wire n_3173;
wire n_4281;
wire n_4345;
wire n_2411;
wire n_4332;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_4210;
wire n_4049;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_3305;
wire n_1572;
wire n_1635;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_4310;
wire n_3786;
wire n_4061;
wire n_1329;
wire n_2637;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3655;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_3050;
wire n_2666;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_4363;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_4196;
wire n_4335;
wire n_2371;
wire n_914;
wire n_3992;
wire n_4147;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4301;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3547;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4267;
wire n_4386;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_2296;
wire n_4342;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_4302;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_1488;
wire n_849;
wire n_980;
wire n_3067;
wire n_3380;
wire n_2227;
wire n_2652;
wire n_2928;
wire n_1074;
wire n_3225;
wire n_3557;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3823;
wire n_3369;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_4266;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_3124;
wire n_999;
wire n_2634;
wire n_3286;
wire n_2982;
wire n_1092;
wire n_4038;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_783;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_4274;
wire n_1062;
wire n_4395;
wire n_1230;
wire n_1516;
wire n_1027;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2303;
wire n_2618;
wire n_2357;
wire n_2653;
wire n_2855;
wire n_3938;
wire n_4354;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_4296;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_4088;
wire n_2136;
wire n_4309;
wire n_4027;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_3056;
wire n_2560;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3189;
wire n_3052;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_4275;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_1762;
wire n_940;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_2168;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_4108;
wire n_2057;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_799;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4226;
wire n_1551;
wire n_3793;
wire n_4153;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_4329;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_4327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_4396;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_809;
wire n_3691;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_4280;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_4394;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1678;
wire n_1091;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_970;
wire n_3654;
wire n_3980;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_4387;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_1655;
wire n_984;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

INVx1_ASAP7_75t_L g772 ( 
.A(n_150),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_523),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_279),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_21),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_182),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_455),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_567),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_115),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_514),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_627),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_747),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_635),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_487),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_539),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_26),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_69),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_258),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_452),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_35),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_40),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_770),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_490),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_759),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_76),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_323),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_764),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_117),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_507),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_162),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_339),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_643),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_762),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_757),
.Y(n_804)
);

BUFx10_ASAP7_75t_L g805 ( 
.A(n_607),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_229),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_506),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_557),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_324),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_72),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_180),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_103),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_3),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_354),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_639),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_278),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_112),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_406),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_249),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_193),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_644),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_312),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_356),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_113),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_125),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_218),
.Y(n_826)
);

BUFx2_ASAP7_75t_SL g827 ( 
.A(n_765),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_614),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_444),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_94),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_497),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_273),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_598),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_508),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_620),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_624),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_676),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_625),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_494),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_599),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_139),
.Y(n_841)
);

INVx1_ASAP7_75t_SL g842 ( 
.A(n_258),
.Y(n_842)
);

INVxp33_ASAP7_75t_L g843 ( 
.A(n_139),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_715),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_451),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_4),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_760),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_555),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_136),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_769),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_657),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_30),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_459),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_538),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_612),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_312),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_318),
.Y(n_857)
);

BUFx5_ASAP7_75t_L g858 ( 
.A(n_690),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_130),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_341),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_265),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_445),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_339),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_281),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_332),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_754),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_392),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_584),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_120),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_2),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_571),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_481),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_559),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_354),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_86),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_372),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_591),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_192),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_512),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_579),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_143),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_250),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_252),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_50),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_684),
.Y(n_885)
);

INVxp67_ASAP7_75t_SL g886 ( 
.A(n_393),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_588),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_87),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_449),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_761),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_131),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_120),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_405),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_61),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_300),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_38),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_424),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_431),
.Y(n_898)
);

BUFx5_ASAP7_75t_L g899 ( 
.A(n_119),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_533),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_609),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_679),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_372),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_528),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_477),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_771),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_78),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_457),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_187),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_534),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_188),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_269),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_500),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_728),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_402),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_529),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_610),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_336),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_768),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_182),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_206),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_93),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_675),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_659),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_418),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_577),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_41),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_556),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_436),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_704),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_541),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_425),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_230),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_463),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_406),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_230),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_102),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_567),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_383),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_269),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_64),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_551),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_362),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_695),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_133),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_429),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_702),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_362),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_683),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_276),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_663),
.Y(n_951)
);

CKINVDCx16_ASAP7_75t_R g952 ( 
.A(n_727),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_475),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_75),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_517),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_242),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_418),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_464),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_597),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_241),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_593),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_552),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_197),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_84),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_474),
.Y(n_965)
);

BUFx10_ASAP7_75t_L g966 ( 
.A(n_190),
.Y(n_966)
);

INVx1_ASAP7_75t_SL g967 ( 
.A(n_758),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_748),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_729),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_611),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_56),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_206),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_300),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_151),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_159),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_426),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_78),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_52),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_39),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_545),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_435),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_735),
.Y(n_982)
);

BUFx8_ASAP7_75t_SL g983 ( 
.A(n_83),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_24),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_678),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_604),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_199),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_530),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_132),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_129),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_631),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_147),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_609),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_487),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_367),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_751),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_227),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_737),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_361),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_298),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_490),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_396),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_701),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_613),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_504),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_58),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_717),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_608),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_183),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_286),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_574),
.Y(n_1011)
);

BUFx8_ASAP7_75t_SL g1012 ( 
.A(n_99),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_596),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_109),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_335),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_543),
.Y(n_1016)
);

INVxp67_ASAP7_75t_SL g1017 ( 
.A(n_31),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_3),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_221),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_562),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_506),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_385),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_590),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_423),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_750),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_352),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_582),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_671),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_474),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_63),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_734),
.Y(n_1031)
);

BUFx10_ASAP7_75t_L g1032 ( 
.A(n_180),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_463),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_236),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_450),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_152),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_548),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_43),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_40),
.Y(n_1039)
);

BUFx2_ASAP7_75t_SL g1040 ( 
.A(n_603),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_585),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_450),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_421),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_219),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_722),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_57),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_135),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_746),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_16),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_98),
.Y(n_1050)
);

BUFx10_ASAP7_75t_L g1051 ( 
.A(n_274),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_376),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_133),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_674),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_0),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_316),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_192),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_480),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_592),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_288),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_677),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_59),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_97),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_12),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_744),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_654),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_328),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_263),
.Y(n_1068)
);

CKINVDCx16_ASAP7_75t_R g1069 ( 
.A(n_703),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_594),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_503),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_64),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_31),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_217),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_749),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_187),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_493),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_19),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_478),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_603),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_546),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_561),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_311),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_209),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_574),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_67),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_5),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_403),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_164),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_200),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_525),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_386),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_745),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_556),
.Y(n_1094)
);

INVx1_ASAP7_75t_SL g1095 ( 
.A(n_248),
.Y(n_1095)
);

BUFx5_ASAP7_75t_L g1096 ( 
.A(n_587),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_128),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_742),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_711),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_126),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_234),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_688),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_87),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_600),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_342),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_1),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_69),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_766),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_433),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_393),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_467),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_265),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_619),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_740),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_503),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_448),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_218),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_39),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_378),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_65),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_752),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_159),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_595),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_132),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_589),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_601),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_136),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_66),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_113),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_241),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_368),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_6),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_341),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_334),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_298),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_435),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_405),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_100),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_656),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_73),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_616),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_755),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_681),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_161),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_305),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_549),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_27),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_606),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_63),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_579),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_489),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_17),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_482),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_718),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_251),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_586),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_636),
.Y(n_1157)
);

INVx1_ASAP7_75t_SL g1158 ( 
.A(n_444),
.Y(n_1158)
);

CKINVDCx16_ASAP7_75t_R g1159 ( 
.A(n_246),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_598),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_472),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_54),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_248),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_705),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_163),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_363),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_22),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_16),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_653),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_322),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_455),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_338),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_183),
.Y(n_1173)
);

BUFx10_ASAP7_75t_L g1174 ( 
.A(n_138),
.Y(n_1174)
);

BUFx2_ASAP7_75t_SL g1175 ( 
.A(n_168),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_285),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_375),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_712),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_402),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_403),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_648),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_541),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_437),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_0),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_146),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_58),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_173),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_293),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_23),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_89),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_443),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_615),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_767),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_27),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_523),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_315),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_232),
.Y(n_1197)
);

BUFx8_ASAP7_75t_SL g1198 ( 
.A(n_124),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_186),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_54),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_439),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_231),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_141),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_739),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_140),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_652),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_114),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_559),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_617),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_615),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_427),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_198),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_515),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_173),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_348),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_743),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_137),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_263),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_586),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_349),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_100),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_756),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_605),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_480),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_274),
.Y(n_1225)
);

CKINVDCx16_ASAP7_75t_R g1226 ( 
.A(n_89),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_90),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_583),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_483),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_763),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_467),
.Y(n_1231)
);

BUFx10_ASAP7_75t_L g1232 ( 
.A(n_532),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_417),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_502),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_630),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_371),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_342),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_565),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_419),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_546),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_680),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_651),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_473),
.Y(n_1243)
);

CKINVDCx16_ASAP7_75t_R g1244 ( 
.A(n_753),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_602),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_325),
.Y(n_1246)
);

INVxp67_ASAP7_75t_SL g1247 ( 
.A(n_940),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_940),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_786),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_940),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_843),
.Y(n_1251)
);

CKINVDCx16_ASAP7_75t_R g1252 ( 
.A(n_1159),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_1226),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_793),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_983),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_969),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1181),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_859),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_859),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1204),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_873),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_873),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_936),
.Y(n_1263)
);

INVxp67_ASAP7_75t_SL g1264 ( 
.A(n_843),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_936),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_952),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1231),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1231),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_793),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1240),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1240),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1069),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_776),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1244),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_776),
.Y(n_1275)
);

CKINVDCx14_ASAP7_75t_R g1276 ( 
.A(n_837),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_988),
.Y(n_1277)
);

INVxp33_ASAP7_75t_SL g1278 ( 
.A(n_1115),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_795),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_983),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_791),
.Y(n_1281)
);

INVxp33_ASAP7_75t_L g1282 ( 
.A(n_1020),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_791),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1012),
.Y(n_1284)
);

INVxp33_ASAP7_75t_L g1285 ( 
.A(n_1125),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1012),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_801),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_801),
.Y(n_1288)
);

INVxp67_ASAP7_75t_SL g1289 ( 
.A(n_1171),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_806),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_806),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_795),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_810),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1198),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_813),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_896),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_810),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_816),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_816),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1198),
.Y(n_1300)
);

CKINVDCx16_ASAP7_75t_R g1301 ( 
.A(n_805),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_785),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_956),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_956),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_837),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_986),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_986),
.Y(n_1307)
);

INVx2_ASAP7_75t_SL g1308 ( 
.A(n_805),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1007),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1000),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1000),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1007),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1030),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1030),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1057),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1061),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1057),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1061),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1075),
.Y(n_1319)
);

INVxp67_ASAP7_75t_L g1320 ( 
.A(n_1049),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1063),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_813),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_1063),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1075),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1132),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1132),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1189),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1189),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1197),
.Y(n_1329)
);

INVxp33_ASAP7_75t_SL g1330 ( 
.A(n_773),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1197),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1217),
.Y(n_1332)
);

CKINVDCx16_ASAP7_75t_R g1333 ( 
.A(n_805),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_1217),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_899),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1204),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_823),
.Y(n_1337)
);

INVxp67_ASAP7_75t_SL g1338 ( 
.A(n_899),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1157),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_899),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_899),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_899),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_899),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_899),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1096),
.Y(n_1345)
);

INVxp33_ASAP7_75t_SL g1346 ( 
.A(n_774),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1157),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1096),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_775),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_823),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_832),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1096),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1096),
.Y(n_1353)
);

CKINVDCx16_ASAP7_75t_R g1354 ( 
.A(n_966),
.Y(n_1354)
);

INVxp33_ASAP7_75t_SL g1355 ( 
.A(n_779),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_1092),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_780),
.Y(n_1357)
);

INVxp67_ASAP7_75t_SL g1358 ( 
.A(n_1096),
.Y(n_1358)
);

INVxp33_ASAP7_75t_SL g1359 ( 
.A(n_784),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_832),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_840),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1096),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1096),
.Y(n_1363)
);

INVx4_ASAP7_75t_R g1364 ( 
.A(n_802),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1109),
.Y(n_1365)
);

INVxp33_ASAP7_75t_SL g1366 ( 
.A(n_789),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_796),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1130),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_858),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_798),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_809),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1149),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1160),
.Y(n_1373)
);

CKINVDCx16_ASAP7_75t_R g1374 ( 
.A(n_966),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_772),
.Y(n_1375)
);

INVxp33_ASAP7_75t_SL g1376 ( 
.A(n_811),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_812),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_814),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_840),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_777),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_778),
.Y(n_1381)
);

INVxp33_ASAP7_75t_SL g1382 ( 
.A(n_817),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_788),
.Y(n_1383)
);

CKINVDCx16_ASAP7_75t_R g1384 ( 
.A(n_966),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_790),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_1351),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1248),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1251),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1251),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1357),
.Y(n_1390)
);

AND2x6_ASAP7_75t_L g1391 ( 
.A(n_1250),
.B(n_944),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1276),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1260),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1264),
.B(n_799),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1247),
.B(n_1256),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_1351),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1257),
.B(n_923),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1335),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1365),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1335),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1348),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1368),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1260),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1372),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1373),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1361),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1357),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1349),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1348),
.Y(n_1409)
);

INVx4_ASAP7_75t_L g1410 ( 
.A(n_1308),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1323),
.B(n_947),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1340),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1258),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1370),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1341),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1342),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1361),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1276),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1254),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1259),
.Y(n_1420)
);

INVx6_ASAP7_75t_L g1421 ( 
.A(n_1301),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1261),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1262),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1263),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1265),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1334),
.B(n_1230),
.Y(n_1426)
);

BUFx8_ASAP7_75t_L g1427 ( 
.A(n_1249),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1369),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1267),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1296),
.B(n_800),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1268),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1305),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1270),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1320),
.B(n_924),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1343),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1356),
.B(n_1239),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1344),
.Y(n_1437)
);

INVxp33_ASAP7_75t_L g1438 ( 
.A(n_1367),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1309),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1260),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1282),
.B(n_782),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1271),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1260),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1338),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1358),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1282),
.B(n_1243),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1345),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1312),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1352),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1369),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1316),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1333),
.B(n_1354),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1285),
.B(n_803),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1353),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1362),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1336),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1336),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1318),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_1330),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1336),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1336),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1363),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1273),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1275),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1281),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1285),
.B(n_1032),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1283),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1319),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1324),
.Y(n_1469)
);

OA21x2_ASAP7_75t_L g1470 ( 
.A1(n_1375),
.A2(n_991),
.B(n_847),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1269),
.A2(n_861),
.B1(n_863),
.B2(n_841),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1289),
.B(n_807),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1287),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1371),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1367),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1377),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1288),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1290),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1380),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1291),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1293),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1297),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1298),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1299),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1303),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1381),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1302),
.B(n_808),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1339),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1304),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1347),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1277),
.B(n_1032),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1374),
.B(n_1032),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1302),
.B(n_1245),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1383),
.B(n_819),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1278),
.B(n_818),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1384),
.B(n_1355),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1252),
.B(n_1051),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1385),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1306),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1266),
.A2(n_824),
.B1(n_826),
.B2(n_822),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1307),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1310),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1311),
.B(n_1313),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1280),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1378),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1279),
.A2(n_861),
.B1(n_863),
.B2(n_841),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1314),
.B(n_1234),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1315),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1317),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1321),
.Y(n_1510)
);

CKINVDCx20_ASAP7_75t_R g1511 ( 
.A(n_1292),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1325),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1272),
.B(n_1051),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1326),
.B(n_820),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1327),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1284),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1328),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1329),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1346),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1331),
.Y(n_1520)
);

INVx5_ASAP7_75t_L g1521 ( 
.A(n_1364),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1332),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1274),
.B(n_1051),
.Y(n_1523)
);

CKINVDCx11_ASAP7_75t_R g1524 ( 
.A(n_1295),
.Y(n_1524)
);

INVx4_ASAP7_75t_L g1525 ( 
.A(n_1286),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1382),
.B(n_804),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1255),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1294),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1253),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1300),
.B(n_825),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1359),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1366),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1376),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1322),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_1337),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1350),
.A2(n_828),
.B1(n_831),
.B2(n_829),
.Y(n_1536)
);

INVx6_ASAP7_75t_L g1537 ( 
.A(n_1360),
.Y(n_1537)
);

AND2x6_ASAP7_75t_L g1538 ( 
.A(n_1379),
.B(n_944),
.Y(n_1538)
);

CKINVDCx16_ASAP7_75t_R g1539 ( 
.A(n_1301),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1264),
.B(n_830),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1264),
.B(n_1227),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1248),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1296),
.B(n_821),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1278),
.A2(n_834),
.B1(n_848),
.B2(n_845),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1276),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1248),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1365),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1365),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1365),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1276),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1264),
.B(n_846),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1264),
.B(n_849),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1260),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1260),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1264),
.B(n_854),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1365),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1260),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1365),
.Y(n_1558)
);

INVx4_ASAP7_75t_L g1559 ( 
.A(n_1308),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1248),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1369),
.A2(n_991),
.B(n_847),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1260),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1365),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1365),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1365),
.Y(n_1565)
);

CKINVDCx16_ASAP7_75t_R g1566 ( 
.A(n_1301),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1260),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1264),
.B(n_855),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1251),
.B(n_1174),
.Y(n_1569)
);

OA21x2_ASAP7_75t_L g1570 ( 
.A1(n_1369),
.A2(n_1113),
.B(n_1108),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1251),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1365),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1248),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1365),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1260),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1251),
.Y(n_1576)
);

AOI22x1_ASAP7_75t_SL g1577 ( 
.A1(n_1351),
.A2(n_878),
.B1(n_884),
.B2(n_882),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1276),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1365),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1365),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1264),
.B(n_856),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1248),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1365),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_1276),
.Y(n_1584)
);

NAND2xp33_ASAP7_75t_L g1585 ( 
.A(n_1251),
.B(n_858),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1296),
.B(n_835),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1251),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1251),
.A2(n_860),
.B1(n_862),
.B2(n_857),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1251),
.B(n_1174),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1251),
.Y(n_1590)
);

NOR3xp33_ASAP7_75t_L g1591 ( 
.A(n_1252),
.B(n_1017),
.C(n_886),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1251),
.B(n_1174),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1248),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1365),
.Y(n_1594)
);

INVx5_ASAP7_75t_L g1595 ( 
.A(n_1260),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1335),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1251),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_R g1598 ( 
.A(n_1280),
.B(n_781),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1335),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1335),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1248),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1251),
.B(n_787),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1335),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1248),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1365),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1248),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1404),
.Y(n_1607)
);

AOI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1447),
.A2(n_906),
.B(n_866),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1463),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1404),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1444),
.B(n_949),
.C(n_919),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1445),
.B(n_968),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1463),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1463),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1487),
.A2(n_869),
.B1(n_870),
.B2(n_867),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1494),
.B(n_783),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1547),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1389),
.B(n_1232),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1388),
.B(n_839),
.Y(n_1619)
);

BUFx3_ASAP7_75t_L g1620 ( 
.A(n_1421),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1487),
.A2(n_883),
.B1(n_909),
.B2(n_872),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1510),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1547),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1548),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1571),
.B(n_1232),
.Y(n_1625)
);

INVxp33_ASAP7_75t_L g1626 ( 
.A(n_1576),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1510),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1510),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1548),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1394),
.A2(n_911),
.B1(n_915),
.B2(n_910),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1410),
.B(n_967),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1597),
.B(n_982),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_L g1633 ( 
.A(n_1585),
.B(n_1025),
.C(n_998),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1605),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1394),
.A2(n_920),
.B1(n_925),
.B2(n_917),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1479),
.B(n_1045),
.Y(n_1636)
);

AND2x6_ASAP7_75t_L g1637 ( 
.A(n_1492),
.B(n_1031),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1587),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1494),
.B(n_792),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1410),
.B(n_985),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1520),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1520),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1524),
.Y(n_1643)
);

AND2x6_ASAP7_75t_L g1644 ( 
.A(n_1540),
.B(n_1031),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1559),
.B(n_927),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1602),
.B(n_1590),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_1569),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1605),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1541),
.B(n_794),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1399),
.Y(n_1650)
);

BUFx3_ASAP7_75t_L g1651 ( 
.A(n_1421),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1520),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1464),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1486),
.B(n_1048),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1540),
.B(n_797),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1402),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1465),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1427),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1405),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1467),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1438),
.B(n_1232),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1498),
.B(n_1054),
.Y(n_1662)
);

INVxp67_ASAP7_75t_SL g1663 ( 
.A(n_1390),
.Y(n_1663)
);

BUFx10_ASAP7_75t_L g1664 ( 
.A(n_1530),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1501),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1549),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1556),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1473),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1501),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1558),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1551),
.A2(n_934),
.B1(n_935),
.B2(n_931),
.Y(n_1671)
);

NOR2x1p5_ASAP7_75t_L g1672 ( 
.A(n_1525),
.B(n_864),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1477),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1563),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1551),
.B(n_815),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1478),
.Y(n_1676)
);

INVx4_ASAP7_75t_L g1677 ( 
.A(n_1521),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1564),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1561),
.Y(n_1679)
);

OR2x6_ASAP7_75t_L g1680 ( 
.A(n_1519),
.B(n_1040),
.Y(n_1680)
);

NAND2xp33_ASAP7_75t_L g1681 ( 
.A(n_1391),
.B(n_858),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1472),
.B(n_836),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1472),
.B(n_838),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1565),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1441),
.A2(n_942),
.B1(n_943),
.B2(n_939),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1559),
.B(n_1216),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1481),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1552),
.B(n_844),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1572),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1483),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1484),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1555),
.B(n_1568),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1489),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1514),
.A2(n_946),
.B1(n_954),
.B2(n_945),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1499),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1502),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1453),
.B(n_1102),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1581),
.B(n_850),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1514),
.B(n_851),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1574),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1589),
.B(n_1121),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1512),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1518),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1470),
.A2(n_981),
.B1(n_993),
.B2(n_974),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1592),
.Y(n_1705)
);

BUFx6f_ASAP7_75t_L g1706 ( 
.A(n_1470),
.Y(n_1706)
);

INVx5_ASAP7_75t_L g1707 ( 
.A(n_1391),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1579),
.Y(n_1708)
);

AOI21x1_ASAP7_75t_L g1709 ( 
.A1(n_1449),
.A2(n_1154),
.B(n_1139),
.Y(n_1709)
);

BUFx16f_ASAP7_75t_R g1710 ( 
.A(n_1427),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1580),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1583),
.Y(n_1712)
);

BUFx4f_ASAP7_75t_L g1713 ( 
.A(n_1538),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1395),
.B(n_885),
.Y(n_1714)
);

INVx4_ASAP7_75t_SL g1715 ( 
.A(n_1538),
.Y(n_1715)
);

INVx11_ASAP7_75t_L g1716 ( 
.A(n_1538),
.Y(n_1716)
);

INVxp67_ASAP7_75t_SL g1717 ( 
.A(n_1407),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1594),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1515),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1515),
.Y(n_1720)
);

CKINVDCx16_ASAP7_75t_R g1721 ( 
.A(n_1539),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1526),
.B(n_890),
.Y(n_1722)
);

AND2x6_ASAP7_75t_L g1723 ( 
.A(n_1497),
.B(n_1242),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1503),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1517),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1493),
.B(n_1164),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_R g1727 ( 
.A(n_1504),
.B(n_1229),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1517),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1466),
.B(n_1169),
.Y(n_1729)
);

NAND3xp33_ASAP7_75t_L g1730 ( 
.A(n_1455),
.B(n_1178),
.C(n_995),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1387),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1542),
.Y(n_1732)
);

NOR2x1p5_ASAP7_75t_L g1733 ( 
.A(n_1525),
.B(n_865),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1436),
.B(n_902),
.Y(n_1734)
);

BUFx2_ASAP7_75t_L g1735 ( 
.A(n_1408),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1430),
.B(n_914),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1475),
.Y(n_1737)
);

NAND3xp33_ASAP7_75t_L g1738 ( 
.A(n_1570),
.B(n_997),
.C(n_994),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1480),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1480),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1430),
.B(n_930),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1482),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1546),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1596),
.B(n_951),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1482),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1560),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1573),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1491),
.B(n_1446),
.Y(n_1748)
);

NOR3xp33_ASAP7_75t_L g1749 ( 
.A(n_1471),
.B(n_1506),
.C(n_1536),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1582),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1459),
.Y(n_1751)
);

BUFx6f_ASAP7_75t_L g1752 ( 
.A(n_1570),
.Y(n_1752)
);

INVxp67_ASAP7_75t_L g1753 ( 
.A(n_1414),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1566),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1596),
.B(n_996),
.Y(n_1755)
);

INVxp33_ASAP7_75t_L g1756 ( 
.A(n_1534),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1531),
.B(n_1003),
.Y(n_1757)
);

INVx3_ASAP7_75t_L g1758 ( 
.A(n_1485),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1411),
.B(n_1028),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1397),
.B(n_1065),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1485),
.Y(n_1761)
);

INVxp67_ASAP7_75t_SL g1762 ( 
.A(n_1599),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1593),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1474),
.B(n_871),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1521),
.B(n_1002),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1426),
.B(n_1066),
.Y(n_1766)
);

INVx11_ASAP7_75t_L g1767 ( 
.A(n_1538),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1601),
.Y(n_1768)
);

INVxp33_ASAP7_75t_L g1769 ( 
.A(n_1495),
.Y(n_1769)
);

NAND3xp33_ASAP7_75t_L g1770 ( 
.A(n_1599),
.B(n_1005),
.C(n_1004),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1476),
.B(n_842),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1532),
.B(n_1533),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1604),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1508),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1513),
.B(n_1093),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1523),
.B(n_1098),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1509),
.Y(n_1777)
);

AOI21x1_ASAP7_75t_L g1778 ( 
.A1(n_1600),
.A2(n_1113),
.B(n_1108),
.Y(n_1778)
);

CKINVDCx6p67_ASAP7_75t_R g1779 ( 
.A(n_1521),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1522),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1606),
.Y(n_1781)
);

INVx2_ASAP7_75t_SL g1782 ( 
.A(n_1505),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1588),
.B(n_1099),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1428),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1428),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1450),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1413),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1507),
.B(n_1114),
.Y(n_1788)
);

NOR2x1p5_ASAP7_75t_L g1789 ( 
.A(n_1516),
.B(n_874),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1434),
.B(n_1142),
.Y(n_1790)
);

INVx2_ASAP7_75t_SL g1791 ( 
.A(n_1527),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1450),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1591),
.A2(n_1014),
.B1(n_1023),
.B2(n_1006),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1543),
.B(n_1143),
.Y(n_1794)
);

INVx8_ASAP7_75t_L g1795 ( 
.A(n_1391),
.Y(n_1795)
);

INVx2_ASAP7_75t_SL g1796 ( 
.A(n_1530),
.Y(n_1796)
);

BUFx10_ASAP7_75t_L g1797 ( 
.A(n_1392),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1528),
.B(n_1029),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1420),
.Y(n_1799)
);

INVx4_ASAP7_75t_L g1800 ( 
.A(n_1391),
.Y(n_1800)
);

INVx3_ASAP7_75t_L g1801 ( 
.A(n_1422),
.Y(n_1801)
);

INVx2_ASAP7_75t_SL g1802 ( 
.A(n_1452),
.Y(n_1802)
);

INVx3_ASAP7_75t_L g1803 ( 
.A(n_1423),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1424),
.Y(n_1804)
);

BUFx6f_ASAP7_75t_L g1805 ( 
.A(n_1425),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1429),
.Y(n_1806)
);

NAND2xp33_ASAP7_75t_R g1807 ( 
.A(n_1432),
.B(n_875),
.Y(n_1807)
);

INVx5_ASAP7_75t_L g1808 ( 
.A(n_1393),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1431),
.Y(n_1809)
);

AO22x2_ASAP7_75t_L g1810 ( 
.A1(n_1577),
.A2(n_1175),
.B1(n_882),
.B2(n_884),
.Y(n_1810)
);

BUFx2_ASAP7_75t_L g1811 ( 
.A(n_1598),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1433),
.Y(n_1812)
);

INVx4_ASAP7_75t_L g1813 ( 
.A(n_1398),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1442),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1600),
.B(n_1193),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1603),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1603),
.A2(n_1034),
.B1(n_1037),
.B2(n_1033),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1400),
.Y(n_1818)
);

BUFx3_ASAP7_75t_L g1819 ( 
.A(n_1529),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1586),
.Y(n_1820)
);

A2O1A1Ixp33_ASAP7_75t_L g1821 ( 
.A1(n_1412),
.A2(n_1041),
.B(n_1042),
.C(n_1039),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1544),
.A2(n_1052),
.B1(n_1053),
.B2(n_1043),
.Y(n_1822)
);

BUFx6f_ASAP7_75t_L g1823 ( 
.A(n_1393),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1415),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1416),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1435),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_1419),
.Y(n_1827)
);

OAI21xp33_ASAP7_75t_SL g1828 ( 
.A1(n_1437),
.A2(n_1060),
.B(n_1055),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1454),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1401),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1462),
.Y(n_1831)
);

INVx3_ASAP7_75t_L g1832 ( 
.A(n_1409),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1595),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1595),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1500),
.Y(n_1835)
);

BUFx6f_ASAP7_75t_L g1836 ( 
.A(n_1393),
.Y(n_1836)
);

BUFx10_ASAP7_75t_L g1837 ( 
.A(n_1418),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1595),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1496),
.B(n_1206),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1403),
.Y(n_1840)
);

BUFx8_ASAP7_75t_SL g1841 ( 
.A(n_1511),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1403),
.B(n_1209),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1403),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1440),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1440),
.B(n_1222),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1440),
.Y(n_1846)
);

CKINVDCx6p67_ASAP7_75t_R g1847 ( 
.A(n_1535),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1443),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1545),
.B(n_1235),
.Y(n_1849)
);

INVx1_ASAP7_75t_SL g1850 ( 
.A(n_1537),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1443),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1443),
.Y(n_1852)
);

NOR2x1p5_ASAP7_75t_L g1853 ( 
.A(n_1550),
.B(n_876),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1456),
.B(n_858),
.Y(n_1854)
);

INVx3_ASAP7_75t_L g1855 ( 
.A(n_1456),
.Y(n_1855)
);

BUFx4f_ASAP7_75t_L g1856 ( 
.A(n_1535),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1456),
.B(n_858),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1457),
.Y(n_1858)
);

BUFx6f_ASAP7_75t_L g1859 ( 
.A(n_1457),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_SL g1860 ( 
.A1(n_1577),
.A2(n_878),
.B1(n_913),
.B2(n_900),
.Y(n_1860)
);

BUFx2_ASAP7_75t_L g1861 ( 
.A(n_1439),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1578),
.B(n_833),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1457),
.Y(n_1863)
);

INVxp33_ASAP7_75t_L g1864 ( 
.A(n_1535),
.Y(n_1864)
);

INVx2_ASAP7_75t_SL g1865 ( 
.A(n_1537),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1460),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1584),
.B(n_833),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1460),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1460),
.Y(n_1869)
);

INVx4_ASAP7_75t_L g1870 ( 
.A(n_1448),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1461),
.Y(n_1871)
);

INVx2_ASAP7_75t_SL g1872 ( 
.A(n_1451),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1461),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1461),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1553),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1553),
.Y(n_1876)
);

AND3x2_ASAP7_75t_L g1877 ( 
.A(n_1386),
.B(n_913),
.C(n_900),
.Y(n_1877)
);

AOI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1458),
.A2(n_1067),
.B1(n_1068),
.B2(n_1064),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1553),
.Y(n_1879)
);

BUFx2_ASAP7_75t_L g1880 ( 
.A(n_1468),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1554),
.Y(n_1881)
);

AOI21x1_ASAP7_75t_L g1882 ( 
.A1(n_1554),
.A2(n_1241),
.B(n_1085),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_SL g1883 ( 
.A(n_1469),
.B(n_833),
.Y(n_1883)
);

BUFx3_ASAP7_75t_L g1884 ( 
.A(n_1488),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1554),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1557),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1557),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1490),
.B(n_877),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_SL g1889 ( 
.A1(n_1396),
.A2(n_916),
.B1(n_1027),
.B2(n_1022),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1557),
.B(n_833),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1406),
.Y(n_1891)
);

HB1xp67_ASAP7_75t_L g1892 ( 
.A(n_1417),
.Y(n_1892)
);

BUFx4f_ASAP7_75t_L g1893 ( 
.A(n_1562),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1562),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1575),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1562),
.B(n_1077),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1567),
.B(n_852),
.Y(n_1897)
);

AND3x2_ASAP7_75t_L g1898 ( 
.A(n_1567),
.B(n_1022),
.C(n_916),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1567),
.Y(n_1899)
);

INVx4_ASAP7_75t_L g1900 ( 
.A(n_1575),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1575),
.B(n_879),
.Y(n_1901)
);

INVx2_ASAP7_75t_SL g1902 ( 
.A(n_1388),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1404),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1389),
.B(n_880),
.Y(n_1904)
);

AOI22x1_ASAP7_75t_L g1905 ( 
.A1(n_1480),
.A2(n_1241),
.B1(n_827),
.B2(n_1204),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1769),
.B(n_868),
.Y(n_1906)
);

INVx2_ASAP7_75t_SL g1907 ( 
.A(n_1751),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1724),
.B(n_881),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1650),
.Y(n_1909)
);

OAI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1762),
.A2(n_1046),
.B1(n_1100),
.B2(n_1027),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1656),
.Y(n_1911)
);

NAND2x1p5_ASAP7_75t_L g1912 ( 
.A(n_1751),
.B(n_853),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1758),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_L g1914 ( 
.A(n_1620),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1758),
.A2(n_1100),
.B1(n_1105),
.B2(n_1046),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1659),
.Y(n_1916)
);

HB1xp67_ASAP7_75t_L g1917 ( 
.A(n_1638),
.Y(n_1917)
);

BUFx6f_ASAP7_75t_L g1918 ( 
.A(n_1651),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1805),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1666),
.Y(n_1920)
);

CKINVDCx8_ASAP7_75t_R g1921 ( 
.A(n_1643),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1646),
.B(n_1105),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1902),
.B(n_1086),
.Y(n_1923)
);

INVx2_ASAP7_75t_SL g1924 ( 
.A(n_1664),
.Y(n_1924)
);

BUFx2_ASAP7_75t_L g1925 ( 
.A(n_1735),
.Y(n_1925)
);

INVx3_ASAP7_75t_L g1926 ( 
.A(n_1870),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1820),
.B(n_1667),
.Y(n_1927)
);

BUFx2_ASAP7_75t_L g1928 ( 
.A(n_1819),
.Y(n_1928)
);

BUFx4f_ASAP7_75t_L g1929 ( 
.A(n_1710),
.Y(n_1929)
);

INVxp67_ASAP7_75t_L g1930 ( 
.A(n_1737),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1805),
.Y(n_1931)
);

INVx6_ASAP7_75t_L g1932 ( 
.A(n_1797),
.Y(n_1932)
);

AOI22x1_ASAP7_75t_L g1933 ( 
.A1(n_1679),
.A2(n_1204),
.B1(n_1107),
.B2(n_1110),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1805),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1670),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1626),
.B(n_1135),
.Y(n_1936)
);

CKINVDCx6p67_ASAP7_75t_R g1937 ( 
.A(n_1721),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1674),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1678),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1772),
.B(n_1647),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1705),
.B(n_1135),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1896),
.Y(n_1942)
);

OR2x2_ASAP7_75t_SL g1943 ( 
.A(n_1721),
.B(n_1163),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1684),
.Y(n_1944)
);

AND3x1_ASAP7_75t_L g1945 ( 
.A(n_1749),
.B(n_1188),
.C(n_1163),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1689),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1700),
.Y(n_1947)
);

BUFx6f_ASAP7_75t_L g1948 ( 
.A(n_1893),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1663),
.B(n_1188),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1739),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1896),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1665),
.Y(n_1952)
);

OAI22xp5_ASAP7_75t_SL g1953 ( 
.A1(n_1860),
.A2(n_1210),
.B1(n_1212),
.B2(n_1191),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1870),
.Y(n_1954)
);

BUFx2_ASAP7_75t_L g1955 ( 
.A(n_1727),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1717),
.B(n_1753),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1665),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1708),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_1841),
.Y(n_1959)
);

NAND2x1_ASAP7_75t_L g1960 ( 
.A(n_1800),
.B(n_852),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1711),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1782),
.B(n_1191),
.Y(n_1962)
);

AO22x2_ASAP7_75t_L g1963 ( 
.A1(n_1710),
.A2(n_1212),
.B1(n_1229),
.B2(n_1210),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1904),
.B(n_1238),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1669),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1712),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1800),
.B(n_887),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1718),
.Y(n_1968)
);

AND2x2_ASAP7_75t_SL g1969 ( 
.A(n_1861),
.B(n_1238),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1658),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1669),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1787),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1816),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1748),
.B(n_889),
.Y(n_1974)
);

AND2x4_ASAP7_75t_L g1975 ( 
.A(n_1672),
.B(n_1091),
.Y(n_1975)
);

INVxp67_ASAP7_75t_L g1976 ( 
.A(n_1619),
.Y(n_1976)
);

INVx4_ASAP7_75t_L g1977 ( 
.A(n_1795),
.Y(n_1977)
);

BUFx6f_ASAP7_75t_L g1978 ( 
.A(n_1893),
.Y(n_1978)
);

INVx3_ASAP7_75t_L g1979 ( 
.A(n_1779),
.Y(n_1979)
);

AND2x6_ASAP7_75t_L g1980 ( 
.A(n_1801),
.B(n_1117),
.Y(n_1980)
);

AO21x2_ASAP7_75t_L g1981 ( 
.A1(n_1738),
.A2(n_1778),
.B(n_1709),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1677),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1764),
.B(n_1233),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1799),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1645),
.B(n_888),
.Y(n_1985)
);

INVx2_ASAP7_75t_SL g1986 ( 
.A(n_1664),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1661),
.B(n_958),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1801),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1803),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1733),
.B(n_1118),
.Y(n_1990)
);

NAND3x1_ASAP7_75t_L g1991 ( 
.A(n_1822),
.B(n_1128),
.C(n_1120),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1803),
.Y(n_1992)
);

CKINVDCx20_ASAP7_75t_R g1993 ( 
.A(n_1880),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1804),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1771),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1806),
.Y(n_1996)
);

BUFx2_ASAP7_75t_L g1997 ( 
.A(n_1898),
.Y(n_1997)
);

INVx4_ASAP7_75t_L g1998 ( 
.A(n_1795),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1740),
.Y(n_1999)
);

BUFx3_ASAP7_75t_L g2000 ( 
.A(n_1847),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1765),
.B(n_1131),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1809),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1765),
.B(n_1791),
.Y(n_2003)
);

CKINVDCx20_ASAP7_75t_R g2004 ( 
.A(n_1827),
.Y(n_2004)
);

NAND2x1p5_ASAP7_75t_L g2005 ( 
.A(n_1811),
.B(n_964),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1645),
.B(n_891),
.Y(n_2006)
);

OR2x2_ASAP7_75t_L g2007 ( 
.A(n_1889),
.B(n_1056),
.Y(n_2007)
);

BUFx3_ASAP7_75t_L g2008 ( 
.A(n_1856),
.Y(n_2008)
);

A2O1A1Ixp33_ASAP7_75t_L g2009 ( 
.A1(n_1742),
.A2(n_1745),
.B(n_1761),
.C(n_1611),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1798),
.B(n_1134),
.Y(n_2010)
);

INVx2_ASAP7_75t_SL g2011 ( 
.A(n_1856),
.Y(n_2011)
);

AOI22xp5_ASAP7_75t_L g2012 ( 
.A1(n_1723),
.A2(n_892),
.B1(n_894),
.B2(n_893),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1813),
.Y(n_2013)
);

INVx2_ASAP7_75t_SL g2014 ( 
.A(n_1680),
.Y(n_2014)
);

CKINVDCx14_ASAP7_75t_R g2015 ( 
.A(n_1891),
.Y(n_2015)
);

INVx1_ASAP7_75t_SL g2016 ( 
.A(n_1850),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1813),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1613),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1613),
.Y(n_2019)
);

AND2x4_ASAP7_75t_L g2020 ( 
.A(n_1798),
.B(n_1136),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1618),
.B(n_1078),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1613),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1812),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_L g2024 ( 
.A(n_1802),
.B(n_898),
.Y(n_2024)
);

AOI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1723),
.A2(n_895),
.B1(n_903),
.B2(n_901),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1814),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1774),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1777),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_SL g2029 ( 
.A(n_1884),
.B(n_1872),
.Y(n_2029)
);

BUFx4f_ASAP7_75t_L g2030 ( 
.A(n_1680),
.Y(n_2030)
);

BUFx6f_ASAP7_75t_L g2031 ( 
.A(n_1706),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1715),
.B(n_1145),
.Y(n_2032)
);

AND2x6_ASAP7_75t_L g2033 ( 
.A(n_1795),
.B(n_1148),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1780),
.Y(n_2034)
);

INVx1_ASAP7_75t_SL g2035 ( 
.A(n_1850),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1731),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1732),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1607),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1743),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1746),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1747),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1750),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1715),
.B(n_1150),
.Y(n_2043)
);

NOR2xp33_ASAP7_75t_L g2044 ( 
.A(n_1835),
.B(n_904),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1763),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1610),
.Y(n_2046)
);

AND2x4_ASAP7_75t_L g2047 ( 
.A(n_1677),
.B(n_1151),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_1796),
.B(n_907),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1625),
.B(n_1083),
.Y(n_2049)
);

AND2x4_ASAP7_75t_L g2050 ( 
.A(n_1680),
.B(n_1162),
.Y(n_2050)
);

INVx1_ASAP7_75t_SL g2051 ( 
.A(n_1877),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1768),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_L g2053 ( 
.A(n_1706),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1714),
.B(n_908),
.Y(n_2054)
);

HB1xp67_ASAP7_75t_L g2055 ( 
.A(n_1807),
.Y(n_2055)
);

A2O1A1Ixp33_ASAP7_75t_L g2056 ( 
.A1(n_1611),
.A2(n_1173),
.B(n_1176),
.C(n_1168),
.Y(n_2056)
);

AO22x2_ASAP7_75t_L g2057 ( 
.A1(n_1810),
.A2(n_1146),
.B1(n_1158),
.B2(n_1095),
.Y(n_2057)
);

BUFx3_ASAP7_75t_L g2058 ( 
.A(n_1754),
.Y(n_2058)
);

CKINVDCx16_ASAP7_75t_R g2059 ( 
.A(n_1797),
.Y(n_2059)
);

INVx3_ASAP7_75t_L g2060 ( 
.A(n_1837),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1773),
.Y(n_2061)
);

INVx3_ASAP7_75t_L g2062 ( 
.A(n_1837),
.Y(n_2062)
);

AO22x2_ASAP7_75t_L g2063 ( 
.A1(n_1810),
.A2(n_1172),
.B1(n_1179),
.B2(n_1177),
.Y(n_2063)
);

INVx3_ASAP7_75t_L g2064 ( 
.A(n_1719),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1615),
.B(n_912),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1706),
.Y(n_2066)
);

AND2x4_ASAP7_75t_L g2067 ( 
.A(n_1616),
.B(n_1182),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1729),
.B(n_918),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1824),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_1639),
.B(n_1201),
.Y(n_2070)
);

AO22x2_ASAP7_75t_L g2071 ( 
.A1(n_1738),
.A2(n_1214),
.B1(n_1221),
.B2(n_1211),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_1752),
.Y(n_2072)
);

AND2x4_ASAP7_75t_L g2073 ( 
.A(n_1775),
.B(n_1223),
.Y(n_2073)
);

BUFx6f_ASAP7_75t_L g2074 ( 
.A(n_1752),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1781),
.Y(n_2075)
);

AOI22xp5_ASAP7_75t_L g2076 ( 
.A1(n_1723),
.A2(n_922),
.B1(n_926),
.B2(n_921),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1653),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1729),
.B(n_928),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1825),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_L g2080 ( 
.A(n_1756),
.B(n_929),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1826),
.Y(n_2081)
);

NAND2x1p5_ASAP7_75t_L g2082 ( 
.A(n_1865),
.B(n_1224),
.Y(n_2082)
);

INVx3_ASAP7_75t_L g2083 ( 
.A(n_1720),
.Y(n_2083)
);

NOR2xp33_ASAP7_75t_L g2084 ( 
.A(n_1682),
.B(n_932),
.Y(n_2084)
);

AND2x4_ASAP7_75t_L g2085 ( 
.A(n_1776),
.B(n_1225),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1657),
.Y(n_2086)
);

AND2x4_ASAP7_75t_L g2087 ( 
.A(n_1699),
.B(n_1236),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1632),
.B(n_933),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_1723),
.A2(n_938),
.B1(n_941),
.B2(n_937),
.Y(n_2089)
);

INVx2_ASAP7_75t_SL g2090 ( 
.A(n_1637),
.Y(n_2090)
);

INVxp67_ASAP7_75t_L g2091 ( 
.A(n_1644),
.Y(n_2091)
);

BUFx4f_ASAP7_75t_L g2092 ( 
.A(n_1637),
.Y(n_2092)
);

OR2x2_ASAP7_75t_SL g2093 ( 
.A(n_1892),
.B(n_1888),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1660),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_SL g2095 ( 
.A(n_1707),
.B(n_948),
.Y(n_2095)
);

AND2x4_ASAP7_75t_L g2096 ( 
.A(n_1655),
.B(n_1237),
.Y(n_2096)
);

INVx3_ASAP7_75t_L g2097 ( 
.A(n_1725),
.Y(n_2097)
);

BUFx2_ASAP7_75t_L g2098 ( 
.A(n_1644),
.Y(n_2098)
);

AND2x4_ASAP7_75t_L g2099 ( 
.A(n_1675),
.B(n_1246),
.Y(n_2099)
);

BUFx6f_ASAP7_75t_L g2100 ( 
.A(n_1752),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1668),
.Y(n_2101)
);

OAI221xp5_ASAP7_75t_L g2102 ( 
.A1(n_1822),
.A2(n_953),
.B1(n_957),
.B2(n_955),
.C(n_950),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1713),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1673),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1676),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_1683),
.B(n_852),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_1615),
.B(n_959),
.Y(n_2107)
);

HB1xp67_ASAP7_75t_L g2108 ( 
.A(n_1644),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1632),
.B(n_960),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1617),
.Y(n_2110)
);

INVx1_ASAP7_75t_SL g2111 ( 
.A(n_1644),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1687),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_1621),
.B(n_961),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1623),
.Y(n_2114)
);

BUFx2_ASAP7_75t_L g2115 ( 
.A(n_1828),
.Y(n_2115)
);

INVx1_ASAP7_75t_SL g2116 ( 
.A(n_1901),
.Y(n_2116)
);

NOR2xp33_ASAP7_75t_L g2117 ( 
.A(n_1736),
.B(n_962),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1624),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1629),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1701),
.B(n_963),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_1621),
.B(n_965),
.Y(n_2121)
);

AOI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_1635),
.A2(n_971),
.B1(n_972),
.B2(n_970),
.Y(n_2122)
);

BUFx6f_ASAP7_75t_L g2123 ( 
.A(n_1713),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1690),
.Y(n_2124)
);

INVx4_ASAP7_75t_SL g2125 ( 
.A(n_1637),
.Y(n_2125)
);

BUFx3_ASAP7_75t_L g2126 ( 
.A(n_1833),
.Y(n_2126)
);

AND2x6_ASAP7_75t_L g2127 ( 
.A(n_1634),
.B(n_852),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1691),
.Y(n_2128)
);

INVx5_ASAP7_75t_L g2129 ( 
.A(n_1637),
.Y(n_2129)
);

AND3x4_ASAP7_75t_L g2130 ( 
.A(n_1789),
.B(n_975),
.C(n_973),
.Y(n_2130)
);

AND2x6_ASAP7_75t_L g2131 ( 
.A(n_1648),
.B(n_897),
.Y(n_2131)
);

INVx3_ASAP7_75t_L g2132 ( 
.A(n_1728),
.Y(n_2132)
);

AND2x6_ASAP7_75t_L g2133 ( 
.A(n_1903),
.B(n_897),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1701),
.B(n_976),
.Y(n_2134)
);

INVxp67_ASAP7_75t_L g2135 ( 
.A(n_1736),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_1707),
.B(n_977),
.Y(n_2136)
);

AND2x4_ASAP7_75t_L g2137 ( 
.A(n_1853),
.B(n_897),
.Y(n_2137)
);

INVx4_ASAP7_75t_L g2138 ( 
.A(n_1707),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1693),
.Y(n_2139)
);

BUFx6f_ASAP7_75t_L g2140 ( 
.A(n_1679),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1695),
.Y(n_2141)
);

AND2x4_ASAP7_75t_L g2142 ( 
.A(n_1692),
.B(n_897),
.Y(n_2142)
);

INVxp67_ASAP7_75t_L g2143 ( 
.A(n_1741),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_1635),
.B(n_978),
.Y(n_2144)
);

OAI22xp5_ASAP7_75t_SL g2145 ( 
.A1(n_1793),
.A2(n_979),
.B1(n_984),
.B2(n_980),
.Y(n_2145)
);

AO22x2_ASAP7_75t_L g2146 ( 
.A1(n_1783),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1696),
.Y(n_2147)
);

NOR2xp33_ASAP7_75t_L g2148 ( 
.A(n_1741),
.B(n_987),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1702),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1630),
.B(n_1671),
.Y(n_2150)
);

BUFx2_ASAP7_75t_L g2151 ( 
.A(n_1828),
.Y(n_2151)
);

OAI21xp33_ASAP7_75t_L g2152 ( 
.A1(n_1878),
.A2(n_1215),
.B(n_1213),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1703),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1726),
.B(n_989),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1832),
.Y(n_2155)
);

INVx4_ASAP7_75t_L g2156 ( 
.A(n_1716),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1829),
.Y(n_2157)
);

AND2x4_ASAP7_75t_L g2158 ( 
.A(n_1883),
.B(n_905),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1831),
.Y(n_2159)
);

XNOR2xp5_ASAP7_75t_L g2160 ( 
.A(n_1878),
.B(n_990),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1612),
.Y(n_2161)
);

AND2x4_ASAP7_75t_L g2162 ( 
.A(n_1839),
.B(n_905),
.Y(n_2162)
);

AO22x2_ASAP7_75t_L g2163 ( 
.A1(n_1726),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1832),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1612),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1636),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1636),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_1685),
.B(n_992),
.Y(n_2168)
);

NAND2x1p5_ASAP7_75t_L g2169 ( 
.A(n_1833),
.B(n_905),
.Y(n_2169)
);

BUFx2_ASAP7_75t_L g2170 ( 
.A(n_1744),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1654),
.Y(n_2171)
);

BUFx6f_ASAP7_75t_L g2172 ( 
.A(n_1679),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_1685),
.B(n_999),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1654),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1662),
.Y(n_2175)
);

INVx2_ASAP7_75t_SL g2176 ( 
.A(n_1862),
.Y(n_2176)
);

INVx3_ASAP7_75t_L g2177 ( 
.A(n_1767),
.Y(n_2177)
);

NAND2x1p5_ASAP7_75t_L g2178 ( 
.A(n_1867),
.B(n_905),
.Y(n_2178)
);

AOI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_1757),
.A2(n_1001),
.B1(n_1009),
.B2(n_1008),
.Y(n_2179)
);

INVx2_ASAP7_75t_SL g2180 ( 
.A(n_1788),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1662),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1784),
.Y(n_2182)
);

AOI22x1_ASAP7_75t_L g2183 ( 
.A1(n_1609),
.A2(n_1141),
.B1(n_1161),
.B2(n_1019),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1785),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1786),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1792),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_SL g2187 ( 
.A(n_1631),
.B(n_1010),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1818),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1830),
.Y(n_2189)
);

AO22x2_ASAP7_75t_L g2190 ( 
.A1(n_1697),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_2190)
);

A2O1A1Ixp33_ASAP7_75t_L g2191 ( 
.A1(n_1704),
.A2(n_1011),
.B(n_1015),
.C(n_1013),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1770),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1770),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1730),
.Y(n_2194)
);

AO22x2_ASAP7_75t_L g2195 ( 
.A1(n_1697),
.A2(n_1730),
.B1(n_1633),
.B2(n_1744),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1821),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1755),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1614),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1759),
.B(n_1016),
.Y(n_2199)
);

NOR2xp33_ASAP7_75t_L g2200 ( 
.A(n_1849),
.B(n_1018),
.Y(n_2200)
);

BUFx6f_ASAP7_75t_L g2201 ( 
.A(n_1808),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1755),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1622),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_1627),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1628),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_1766),
.B(n_1021),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1815),
.Y(n_2207)
);

OAI22xp5_ASAP7_75t_L g2208 ( 
.A1(n_1694),
.A2(n_1024),
.B1(n_1035),
.B2(n_1026),
.Y(n_2208)
);

AOI22xp5_ASAP7_75t_L g2209 ( 
.A1(n_1640),
.A2(n_1038),
.B1(n_1044),
.B2(n_1036),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1815),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1641),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1698),
.B(n_1047),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1642),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_SL g2214 ( 
.A(n_1649),
.B(n_1050),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_1722),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1686),
.B(n_1058),
.Y(n_2216)
);

AOI22xp5_ASAP7_75t_L g2217 ( 
.A1(n_1734),
.A2(n_1062),
.B1(n_1070),
.B2(n_1059),
.Y(n_2217)
);

INVx4_ASAP7_75t_L g2218 ( 
.A(n_1808),
.Y(n_2218)
);

HB1xp67_ASAP7_75t_L g2219 ( 
.A(n_1864),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1608),
.Y(n_2220)
);

NOR2xp33_ASAP7_75t_L g2221 ( 
.A(n_1760),
.B(n_1071),
.Y(n_2221)
);

INVx4_ASAP7_75t_SL g2222 ( 
.A(n_1823),
.Y(n_2222)
);

INVxp67_ASAP7_75t_L g2223 ( 
.A(n_1688),
.Y(n_2223)
);

INVx4_ASAP7_75t_L g2224 ( 
.A(n_1808),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1652),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_1854),
.Y(n_2226)
);

AND2x4_ASAP7_75t_L g2227 ( 
.A(n_1790),
.B(n_1019),
.Y(n_2227)
);

INVxp67_ASAP7_75t_L g2228 ( 
.A(n_1794),
.Y(n_2228)
);

AND2x4_ASAP7_75t_L g2229 ( 
.A(n_1817),
.B(n_1019),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_1633),
.B(n_1072),
.Y(n_2230)
);

BUFx6f_ASAP7_75t_L g2231 ( 
.A(n_1834),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1681),
.B(n_1073),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_1854),
.Y(n_2233)
);

AOI22xp5_ASAP7_75t_L g2234 ( 
.A1(n_1842),
.A2(n_1076),
.B1(n_1079),
.B2(n_1074),
.Y(n_2234)
);

INVxp33_ASAP7_75t_L g2235 ( 
.A(n_1905),
.Y(n_2235)
);

INVx3_ASAP7_75t_L g2236 ( 
.A(n_1838),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1842),
.Y(n_2237)
);

OAI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_1845),
.A2(n_1080),
.B1(n_1082),
.B2(n_1081),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1857),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_1845),
.B(n_1084),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1857),
.Y(n_2241)
);

INVx3_ASAP7_75t_L g2242 ( 
.A(n_1900),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_1900),
.B(n_1087),
.Y(n_2243)
);

BUFx6f_ASAP7_75t_L g2244 ( 
.A(n_1882),
.Y(n_2244)
);

INVx8_ASAP7_75t_L g2245 ( 
.A(n_1855),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1890),
.Y(n_2246)
);

BUFx6f_ASAP7_75t_L g2247 ( 
.A(n_1823),
.Y(n_2247)
);

BUFx2_ASAP7_75t_L g2248 ( 
.A(n_1823),
.Y(n_2248)
);

BUFx3_ASAP7_75t_L g2249 ( 
.A(n_1855),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_L g2250 ( 
.A(n_1843),
.B(n_1088),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_1836),
.B(n_1089),
.Y(n_2251)
);

AND2x4_ASAP7_75t_L g2252 ( 
.A(n_1897),
.B(n_1019),
.Y(n_2252)
);

BUFx4f_ASAP7_75t_L g2253 ( 
.A(n_1844),
.Y(n_2253)
);

A2O1A1Ixp33_ASAP7_75t_L g2254 ( 
.A1(n_2197),
.A2(n_1161),
.B(n_1190),
.C(n_1141),
.Y(n_2254)
);

BUFx2_ASAP7_75t_L g2255 ( 
.A(n_1925),
.Y(n_2255)
);

AOI22xp33_ASAP7_75t_L g2256 ( 
.A1(n_1949),
.A2(n_1090),
.B1(n_1097),
.B2(n_1094),
.Y(n_2256)
);

INVx2_ASAP7_75t_SL g2257 ( 
.A(n_1932),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2161),
.B(n_1101),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_1907),
.B(n_1103),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2165),
.B(n_1104),
.Y(n_2260)
);

HB1xp67_ASAP7_75t_L g2261 ( 
.A(n_1925),
.Y(n_2261)
);

HB1xp67_ASAP7_75t_L g2262 ( 
.A(n_1917),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1909),
.Y(n_2263)
);

A2O1A1Ixp33_ASAP7_75t_L g2264 ( 
.A1(n_2202),
.A2(n_1161),
.B(n_1190),
.C(n_1141),
.Y(n_2264)
);

INVx2_ASAP7_75t_SL g2265 ( 
.A(n_1932),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1911),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1916),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1920),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_1930),
.B(n_1106),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_SL g2270 ( 
.A(n_1977),
.B(n_1111),
.Y(n_2270)
);

AOI22xp33_ASAP7_75t_L g2271 ( 
.A1(n_1995),
.A2(n_1112),
.B1(n_1119),
.B2(n_1116),
.Y(n_2271)
);

AOI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_2229),
.A2(n_1122),
.B1(n_1124),
.B2(n_1123),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1935),
.Y(n_2273)
);

AOI22xp33_ASAP7_75t_L g2274 ( 
.A1(n_2168),
.A2(n_1126),
.B1(n_1129),
.B2(n_1127),
.Y(n_2274)
);

BUFx3_ASAP7_75t_L g2275 ( 
.A(n_1928),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1938),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2166),
.B(n_1133),
.Y(n_2277)
);

BUFx2_ASAP7_75t_L g2278 ( 
.A(n_1928),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2167),
.B(n_1137),
.Y(n_2279)
);

BUFx6f_ASAP7_75t_L g2280 ( 
.A(n_2247),
.Y(n_2280)
);

OR2x2_ASAP7_75t_SL g2281 ( 
.A(n_2059),
.B(n_1141),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1939),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2173),
.B(n_1138),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2171),
.B(n_1140),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2174),
.B(n_1144),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2175),
.B(n_1147),
.Y(n_2286)
);

NOR2xp33_ASAP7_75t_L g2287 ( 
.A(n_1906),
.B(n_1152),
.Y(n_2287)
);

INVx5_ASAP7_75t_L g2288 ( 
.A(n_2033),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_1912),
.B(n_1153),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_2030),
.B(n_1155),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2181),
.B(n_1156),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2150),
.B(n_1165),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1944),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1927),
.B(n_1166),
.Y(n_2294)
);

INVx2_ASAP7_75t_SL g2295 ( 
.A(n_1929),
.Y(n_2295)
);

BUFx6f_ASAP7_75t_L g2296 ( 
.A(n_2247),
.Y(n_2296)
);

BUFx2_ASAP7_75t_L g2297 ( 
.A(n_1993),
.Y(n_2297)
);

AND2x4_ASAP7_75t_L g2298 ( 
.A(n_2125),
.B(n_1161),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_SL g2299 ( 
.A(n_2016),
.B(n_1167),
.Y(n_2299)
);

OR2x2_ASAP7_75t_L g2300 ( 
.A(n_1910),
.B(n_1170),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_1946),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1947),
.Y(n_2302)
);

AND2x6_ASAP7_75t_SL g2303 ( 
.A(n_1936),
.B(n_1180),
.Y(n_2303)
);

INVx5_ASAP7_75t_L g2304 ( 
.A(n_2033),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_1976),
.B(n_1183),
.Y(n_2305)
);

BUFx4f_ASAP7_75t_SL g2306 ( 
.A(n_1937),
.Y(n_2306)
);

AOI22xp33_ASAP7_75t_L g2307 ( 
.A1(n_2065),
.A2(n_1184),
.B1(n_1186),
.B2(n_1185),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_2035),
.B(n_1187),
.Y(n_2308)
);

INVx2_ASAP7_75t_SL g2309 ( 
.A(n_2000),
.Y(n_2309)
);

BUFx3_ASAP7_75t_L g2310 ( 
.A(n_1914),
.Y(n_2310)
);

BUFx6f_ASAP7_75t_L g2311 ( 
.A(n_2072),
.Y(n_2311)
);

CKINVDCx5p33_ASAP7_75t_R g2312 ( 
.A(n_1959),
.Y(n_2312)
);

INVx3_ASAP7_75t_L g2313 ( 
.A(n_1977),
.Y(n_2313)
);

BUFx3_ASAP7_75t_L g2314 ( 
.A(n_1914),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2170),
.B(n_1192),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_2125),
.B(n_1190),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2170),
.B(n_1194),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1958),
.Y(n_2318)
);

BUFx3_ASAP7_75t_L g2319 ( 
.A(n_1918),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_2029),
.B(n_1195),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1961),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_SL g2322 ( 
.A(n_1956),
.B(n_1196),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_L g2323 ( 
.A(n_2135),
.B(n_1199),
.Y(n_2323)
);

BUFx2_ASAP7_75t_L g2324 ( 
.A(n_1980),
.Y(n_2324)
);

BUFx3_ASAP7_75t_L g2325 ( 
.A(n_1918),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_1966),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2143),
.B(n_1200),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_SL g2328 ( 
.A(n_2187),
.B(n_1202),
.Y(n_2328)
);

AND2x4_ASAP7_75t_L g2329 ( 
.A(n_2014),
.B(n_1190),
.Y(n_2329)
);

HB1xp67_ASAP7_75t_L g2330 ( 
.A(n_1915),
.Y(n_2330)
);

AOI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_2229),
.A2(n_1203),
.B1(n_1207),
.B2(n_1205),
.Y(n_2331)
);

NOR2xp33_ASAP7_75t_L g2332 ( 
.A(n_1962),
.B(n_1208),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1968),
.Y(n_2333)
);

AND3x1_ASAP7_75t_L g2334 ( 
.A(n_2055),
.B(n_1219),
.C(n_1218),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_SL g2335 ( 
.A(n_2228),
.B(n_1220),
.Y(n_2335)
);

AND2x4_ASAP7_75t_L g2336 ( 
.A(n_1926),
.B(n_8),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_1972),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1984),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2069),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2207),
.B(n_1228),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2069),
.Y(n_2341)
);

BUFx3_ASAP7_75t_L g2342 ( 
.A(n_1921),
.Y(n_2342)
);

OAI21xp33_ASAP7_75t_L g2343 ( 
.A1(n_1940),
.A2(n_1852),
.B(n_1851),
.Y(n_2343)
);

INVx3_ASAP7_75t_L g2344 ( 
.A(n_1998),
.Y(n_2344)
);

BUFx6f_ASAP7_75t_L g2345 ( 
.A(n_2072),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_1999),
.Y(n_2346)
);

AND2x6_ASAP7_75t_L g2347 ( 
.A(n_2111),
.B(n_1836),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_1950),
.Y(n_2348)
);

AND2x6_ASAP7_75t_L g2349 ( 
.A(n_2103),
.B(n_1836),
.Y(n_2349)
);

AND3x2_ASAP7_75t_SL g2350 ( 
.A(n_1963),
.B(n_9),
.C(n_10),
.Y(n_2350)
);

HB1xp67_ASAP7_75t_L g2351 ( 
.A(n_1922),
.Y(n_2351)
);

AND2x4_ASAP7_75t_L g2352 ( 
.A(n_1954),
.B(n_10),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2210),
.B(n_11),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2107),
.B(n_11),
.Y(n_2354)
);

BUFx3_ASAP7_75t_L g2355 ( 
.A(n_2004),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2113),
.B(n_2121),
.Y(n_2356)
);

AOI22xp33_ASAP7_75t_L g2357 ( 
.A1(n_2144),
.A2(n_858),
.B1(n_1871),
.B2(n_1863),
.Y(n_2357)
);

AOI22xp5_ASAP7_75t_L g2358 ( 
.A1(n_2115),
.A2(n_858),
.B1(n_1881),
.B2(n_1879),
.Y(n_2358)
);

NOR2xp33_ASAP7_75t_L g2359 ( 
.A(n_1964),
.B(n_12),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_1924),
.B(n_1859),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2079),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_1950),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2079),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_1986),
.B(n_1859),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2081),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_1980),
.B(n_13),
.Y(n_2366)
);

OAI221xp5_ASAP7_75t_L g2367 ( 
.A1(n_2160),
.A2(n_1894),
.B1(n_1848),
.B2(n_1858),
.C(n_1846),
.Y(n_2367)
);

NAND2xp33_ASAP7_75t_L g2368 ( 
.A(n_1980),
.B(n_1859),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_1973),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2081),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1994),
.Y(n_2371)
);

INVxp67_ASAP7_75t_L g2372 ( 
.A(n_1997),
.Y(n_2372)
);

NOR2x1p5_ASAP7_75t_L g2373 ( 
.A(n_2060),
.B(n_13),
.Y(n_2373)
);

INVx1_ASAP7_75t_SL g2374 ( 
.A(n_2219),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_1996),
.Y(n_2375)
);

NOR2xp67_ASAP7_75t_L g2376 ( 
.A(n_2129),
.B(n_618),
.Y(n_2376)
);

INVx3_ASAP7_75t_L g2377 ( 
.A(n_1998),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2002),
.Y(n_2378)
);

AOI22xp5_ASAP7_75t_L g2379 ( 
.A1(n_2115),
.A2(n_1866),
.B1(n_1868),
.B2(n_1840),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_2129),
.B(n_1869),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2023),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2026),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2151),
.B(n_14),
.Y(n_2383)
);

AOI22xp33_ASAP7_75t_L g2384 ( 
.A1(n_1969),
.A2(n_1874),
.B1(n_1875),
.B2(n_1873),
.Y(n_2384)
);

INVx4_ASAP7_75t_L g2385 ( 
.A(n_2033),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2027),
.Y(n_2386)
);

OAI22xp5_ASAP7_75t_SL g2387 ( 
.A1(n_1943),
.A2(n_17),
.B1(n_14),
.B2(n_15),
.Y(n_2387)
);

AND2x6_ASAP7_75t_SL g2388 ( 
.A(n_1963),
.B(n_15),
.Y(n_2388)
);

AND2x6_ASAP7_75t_L g2389 ( 
.A(n_2103),
.B(n_1876),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2151),
.B(n_18),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2028),
.Y(n_2391)
);

BUFx3_ASAP7_75t_L g2392 ( 
.A(n_2058),
.Y(n_2392)
);

OR2x2_ASAP7_75t_SL g2393 ( 
.A(n_2007),
.B(n_18),
.Y(n_2393)
);

AND2x2_ASAP7_75t_L g2394 ( 
.A(n_2160),
.B(n_19),
.Y(n_2394)
);

OAI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2092),
.A2(n_1899),
.B1(n_1886),
.B2(n_1887),
.Y(n_2395)
);

A2O1A1Ixp33_ASAP7_75t_L g2396 ( 
.A1(n_2044),
.A2(n_1895),
.B(n_1885),
.C(n_22),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2034),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2196),
.B(n_20),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2038),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2154),
.B(n_2240),
.Y(n_2400)
);

BUFx6f_ASAP7_75t_L g2401 ( 
.A(n_2074),
.Y(n_2401)
);

INVx2_ASAP7_75t_SL g2402 ( 
.A(n_2062),
.Y(n_2402)
);

BUFx4f_ASAP7_75t_SL g2403 ( 
.A(n_1979),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2046),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2110),
.Y(n_2405)
);

AOI22xp5_ASAP7_75t_L g2406 ( 
.A1(n_1945),
.A2(n_23),
.B1(n_20),
.B2(n_21),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2010),
.B(n_24),
.Y(n_2407)
);

AOI22xp5_ASAP7_75t_L g2408 ( 
.A1(n_1991),
.A2(n_28),
.B1(n_25),
.B2(n_26),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_1983),
.B(n_25),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2010),
.B(n_28),
.Y(n_2410)
);

BUFx3_ASAP7_75t_L g2411 ( 
.A(n_1970),
.Y(n_2411)
);

INVx4_ASAP7_75t_L g2412 ( 
.A(n_2201),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2036),
.Y(n_2413)
);

AND2x4_ASAP7_75t_L g2414 ( 
.A(n_2003),
.B(n_29),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2114),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2037),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2118),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2020),
.B(n_29),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2039),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2040),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_SL g2421 ( 
.A(n_2129),
.B(n_30),
.Y(n_2421)
);

NAND3xp33_ASAP7_75t_SL g2422 ( 
.A(n_2051),
.B(n_32),
.C(n_33),
.Y(n_2422)
);

INVx3_ASAP7_75t_L g2423 ( 
.A(n_2218),
.Y(n_2423)
);

OAI22xp5_ASAP7_75t_SL g2424 ( 
.A1(n_1953),
.A2(n_2093),
.B1(n_2130),
.B2(n_2005),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2041),
.Y(n_2425)
);

HB1xp67_ASAP7_75t_L g2426 ( 
.A(n_1997),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2020),
.B(n_32),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2119),
.Y(n_2428)
);

NOR2xp33_ASAP7_75t_L g2429 ( 
.A(n_1941),
.B(n_33),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2042),
.Y(n_2430)
);

AND2x4_ASAP7_75t_L g2431 ( 
.A(n_2003),
.B(n_34),
.Y(n_2431)
);

AND2x4_ASAP7_75t_L g2432 ( 
.A(n_2156),
.B(n_34),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_1908),
.B(n_35),
.Y(n_2433)
);

INVx2_ASAP7_75t_SL g2434 ( 
.A(n_2008),
.Y(n_2434)
);

OAI22xp33_ASAP7_75t_L g2435 ( 
.A1(n_1955),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_2015),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2045),
.Y(n_2437)
);

HB1xp67_ASAP7_75t_L g2438 ( 
.A(n_2082),
.Y(n_2438)
);

INVx4_ASAP7_75t_L g2439 ( 
.A(n_2201),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2052),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2061),
.Y(n_2441)
);

NOR2xp33_ASAP7_75t_L g2442 ( 
.A(n_2021),
.B(n_36),
.Y(n_2442)
);

INVx3_ASAP7_75t_L g2443 ( 
.A(n_2218),
.Y(n_2443)
);

AOI22xp33_ASAP7_75t_L g2444 ( 
.A1(n_2102),
.A2(n_42),
.B1(n_37),
.B2(n_41),
.Y(n_2444)
);

NOR2xp33_ASAP7_75t_L g2445 ( 
.A(n_2116),
.B(n_42),
.Y(n_2445)
);

BUFx2_ASAP7_75t_L g2446 ( 
.A(n_1955),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2068),
.B(n_43),
.Y(n_2447)
);

O2A1O1Ixp5_ASAP7_75t_L g2448 ( 
.A1(n_2235),
.A2(n_1960),
.B(n_2227),
.C(n_2220),
.Y(n_2448)
);

NOR3xp33_ASAP7_75t_SL g2449 ( 
.A(n_2215),
.B(n_44),
.C(n_45),
.Y(n_2449)
);

CKINVDCx5p33_ASAP7_75t_R g2450 ( 
.A(n_2137),
.Y(n_2450)
);

NOR2xp33_ASAP7_75t_L g2451 ( 
.A(n_1987),
.B(n_44),
.Y(n_2451)
);

AOI22xp33_ASAP7_75t_L g2452 ( 
.A1(n_2145),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2078),
.B(n_46),
.Y(n_2453)
);

INVx1_ASAP7_75t_SL g2454 ( 
.A(n_2243),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2157),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_SL g2456 ( 
.A(n_2012),
.B(n_47),
.Y(n_2456)
);

NOR2xp67_ASAP7_75t_L g2457 ( 
.A(n_2138),
.B(n_621),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2188),
.Y(n_2458)
);

INVxp67_ASAP7_75t_L g2459 ( 
.A(n_2050),
.Y(n_2459)
);

NOR2x2_ASAP7_75t_L g2460 ( 
.A(n_2057),
.B(n_48),
.Y(n_2460)
);

INVx3_ASAP7_75t_L g2461 ( 
.A(n_2224),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2159),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2075),
.Y(n_2463)
);

OAI22xp5_ASAP7_75t_SL g2464 ( 
.A1(n_2050),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_2464)
);

INVxp67_ASAP7_75t_L g2465 ( 
.A(n_2049),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2120),
.B(n_2134),
.Y(n_2466)
);

NAND2x1p5_ASAP7_75t_L g2467 ( 
.A(n_1948),
.B(n_51),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2077),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2086),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2189),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_SL g2471 ( 
.A(n_2025),
.B(n_49),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_SL g2472 ( 
.A(n_2076),
.B(n_51),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2094),
.Y(n_2473)
);

INVx5_ASAP7_75t_L g2474 ( 
.A(n_1948),
.Y(n_2474)
);

INVx3_ASAP7_75t_L g2475 ( 
.A(n_2224),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2142),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2101),
.Y(n_2477)
);

AND2x4_ASAP7_75t_L g2478 ( 
.A(n_2156),
.B(n_52),
.Y(n_2478)
);

INVx5_ASAP7_75t_L g2479 ( 
.A(n_1978),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2104),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2105),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2112),
.Y(n_2482)
);

NOR2xp33_ASAP7_75t_L g2483 ( 
.A(n_2223),
.B(n_53),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2124),
.Y(n_2484)
);

AOI22xp5_ASAP7_75t_L g2485 ( 
.A1(n_2163),
.A2(n_56),
.B1(n_53),
.B2(n_55),
.Y(n_2485)
);

INVx2_ASAP7_75t_SL g2486 ( 
.A(n_2137),
.Y(n_2486)
);

BUFx3_ASAP7_75t_L g2487 ( 
.A(n_1978),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2142),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_SL g2489 ( 
.A(n_2089),
.B(n_55),
.Y(n_2489)
);

CKINVDCx11_ASAP7_75t_R g2490 ( 
.A(n_1975),
.Y(n_2490)
);

AND2x4_ASAP7_75t_L g2491 ( 
.A(n_2180),
.B(n_57),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_SL g2492 ( 
.A(n_2098),
.B(n_59),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2128),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2139),
.Y(n_2494)
);

BUFx6f_ASAP7_75t_SL g2495 ( 
.A(n_1975),
.Y(n_2495)
);

AOI22xp33_ASAP7_75t_L g2496 ( 
.A1(n_2152),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2141),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_1942),
.Y(n_2498)
);

NAND2x1p5_ASAP7_75t_L g2499 ( 
.A(n_2011),
.B(n_62),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_1951),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2147),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_SL g2502 ( 
.A(n_2098),
.B(n_60),
.Y(n_2502)
);

HB1xp67_ASAP7_75t_L g2503 ( 
.A(n_2251),
.Y(n_2503)
);

AND2x4_ASAP7_75t_L g2504 ( 
.A(n_2106),
.B(n_65),
.Y(n_2504)
);

BUFx3_ASAP7_75t_L g2505 ( 
.A(n_2231),
.Y(n_2505)
);

HB1xp67_ASAP7_75t_L g2506 ( 
.A(n_1923),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2149),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2153),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_L g2509 ( 
.A(n_2117),
.B(n_66),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2047),
.Y(n_2510)
);

NAND2x1p5_ASAP7_75t_L g2511 ( 
.A(n_2253),
.B(n_68),
.Y(n_2511)
);

AOI22xp33_ASAP7_75t_L g2512 ( 
.A1(n_2001),
.A2(n_70),
.B1(n_67),
.B2(n_68),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2186),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_1923),
.B(n_70),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2088),
.B(n_71),
.Y(n_2515)
);

AOI21xp5_ASAP7_75t_L g2516 ( 
.A1(n_2009),
.A2(n_623),
.B(n_622),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2109),
.B(n_71),
.Y(n_2517)
);

AND2x2_ASAP7_75t_L g2518 ( 
.A(n_2122),
.B(n_72),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2047),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2148),
.B(n_73),
.Y(n_2520)
);

NOR3xp33_ASAP7_75t_SL g2521 ( 
.A(n_2084),
.B(n_74),
.C(n_75),
.Y(n_2521)
);

BUFx2_ASAP7_75t_R g2522 ( 
.A(n_1985),
.Y(n_2522)
);

CKINVDCx6p67_ASAP7_75t_R g2523 ( 
.A(n_1990),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2182),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2096),
.B(n_74),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2184),
.Y(n_2526)
);

BUFx6f_ASAP7_75t_L g2527 ( 
.A(n_2074),
.Y(n_2527)
);

INVx6_ASAP7_75t_L g2528 ( 
.A(n_2231),
.Y(n_2528)
);

INVx5_ASAP7_75t_L g2529 ( 
.A(n_2127),
.Y(n_2529)
);

INVx3_ASAP7_75t_L g2530 ( 
.A(n_2138),
.Y(n_2530)
);

NOR2xp33_ASAP7_75t_R g2531 ( 
.A(n_2177),
.B(n_76),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_SL g2532 ( 
.A(n_2006),
.B(n_77),
.Y(n_2532)
);

CKINVDCx5p33_ASAP7_75t_R g2533 ( 
.A(n_1990),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2237),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2185),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2227),
.Y(n_2536)
);

CKINVDCx5p33_ASAP7_75t_R g2537 ( 
.A(n_2208),
.Y(n_2537)
);

AOI22xp33_ASAP7_75t_L g2538 ( 
.A1(n_2001),
.A2(n_80),
.B1(n_77),
.B2(n_79),
.Y(n_2538)
);

AOI22xp5_ASAP7_75t_L g2539 ( 
.A1(n_2163),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2190),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2190),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2096),
.B(n_2099),
.Y(n_2542)
);

BUFx3_ASAP7_75t_L g2543 ( 
.A(n_2126),
.Y(n_2543)
);

HB1xp67_ASAP7_75t_L g2544 ( 
.A(n_2013),
.Y(n_2544)
);

INVx2_ASAP7_75t_SL g2545 ( 
.A(n_2106),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_SL g2546 ( 
.A(n_2080),
.B(n_81),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2099),
.Y(n_2547)
);

NOR2x2_ASAP7_75t_L g2548 ( 
.A(n_2057),
.B(n_82),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2067),
.B(n_82),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2063),
.B(n_83),
.Y(n_2550)
);

BUFx8_ASAP7_75t_L g2551 ( 
.A(n_2162),
.Y(n_2551)
);

INVxp67_ASAP7_75t_L g2552 ( 
.A(n_2048),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_SL g2553 ( 
.A(n_2234),
.B(n_84),
.Y(n_2553)
);

BUFx8_ASAP7_75t_L g2554 ( 
.A(n_2162),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2226),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_SL g2556 ( 
.A(n_2238),
.B(n_85),
.Y(n_2556)
);

NOR2x1p5_ASAP7_75t_L g2557 ( 
.A(n_1982),
.B(n_85),
.Y(n_2557)
);

INVx2_ASAP7_75t_SL g2558 ( 
.A(n_2032),
.Y(n_2558)
);

OR2x6_ASAP7_75t_L g2559 ( 
.A(n_2090),
.B(n_86),
.Y(n_2559)
);

BUFx6f_ASAP7_75t_L g2560 ( 
.A(n_2100),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_2073),
.Y(n_2561)
);

OR2x6_ASAP7_75t_L g2562 ( 
.A(n_2063),
.B(n_88),
.Y(n_2562)
);

INVx4_ASAP7_75t_L g2563 ( 
.A(n_2245),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2067),
.B(n_88),
.Y(n_2564)
);

BUFx8_ASAP7_75t_L g2565 ( 
.A(n_2032),
.Y(n_2565)
);

NOR2xp33_ASAP7_75t_R g2566 ( 
.A(n_2245),
.B(n_90),
.Y(n_2566)
);

AOI21xp5_ASAP7_75t_L g2567 ( 
.A1(n_2220),
.A2(n_628),
.B(n_626),
.Y(n_2567)
);

BUFx6f_ASAP7_75t_L g2568 ( 
.A(n_2100),
.Y(n_2568)
);

INVx1_ASAP7_75t_SL g2569 ( 
.A(n_2043),
.Y(n_2569)
);

INVxp67_ASAP7_75t_L g2570 ( 
.A(n_1974),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2070),
.B(n_91),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2233),
.Y(n_2572)
);

NOR2xp67_ASAP7_75t_L g2573 ( 
.A(n_2091),
.B(n_629),
.Y(n_2573)
);

BUFx8_ASAP7_75t_L g2574 ( 
.A(n_2043),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2070),
.Y(n_2575)
);

INVx5_ASAP7_75t_L g2576 ( 
.A(n_2127),
.Y(n_2576)
);

INVx8_ASAP7_75t_L g2577 ( 
.A(n_2127),
.Y(n_2577)
);

NOR2xp33_ASAP7_75t_L g2578 ( 
.A(n_2200),
.B(n_2024),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2087),
.B(n_91),
.Y(n_2579)
);

INVx2_ASAP7_75t_SL g2580 ( 
.A(n_2087),
.Y(n_2580)
);

AND2x4_ASAP7_75t_L g2581 ( 
.A(n_2073),
.B(n_92),
.Y(n_2581)
);

NOR2xp33_ASAP7_75t_L g2582 ( 
.A(n_2085),
.B(n_92),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2239),
.Y(n_2583)
);

AND2x6_ASAP7_75t_L g2584 ( 
.A(n_2123),
.B(n_1988),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_2085),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2241),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2191),
.B(n_93),
.Y(n_2587)
);

NOR2xp33_ASAP7_75t_L g2588 ( 
.A(n_2214),
.B(n_94),
.Y(n_2588)
);

AND2x4_ASAP7_75t_L g2589 ( 
.A(n_2108),
.B(n_95),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2146),
.Y(n_2590)
);

BUFx3_ASAP7_75t_L g2591 ( 
.A(n_2236),
.Y(n_2591)
);

OAI22xp33_ASAP7_75t_L g2592 ( 
.A1(n_2209),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_2592)
);

NOR3xp33_ASAP7_75t_SL g2593 ( 
.A(n_2221),
.B(n_96),
.C(n_98),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2146),
.Y(n_2594)
);

INVx3_ASAP7_75t_L g2595 ( 
.A(n_2123),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_SL g2596 ( 
.A(n_1913),
.B(n_99),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2155),
.Y(n_2597)
);

NOR2x1p5_ASAP7_75t_L g2598 ( 
.A(n_2216),
.B(n_101),
.Y(n_2598)
);

NOR2x2_ASAP7_75t_L g2599 ( 
.A(n_2017),
.B(n_101),
.Y(n_2599)
);

AND2x4_ASAP7_75t_L g2600 ( 
.A(n_1967),
.B(n_102),
.Y(n_2600)
);

INVx3_ASAP7_75t_L g2601 ( 
.A(n_2242),
.Y(n_2601)
);

AND3x2_ASAP7_75t_SL g2602 ( 
.A(n_2164),
.B(n_103),
.C(n_104),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_1992),
.Y(n_2603)
);

BUFx8_ASAP7_75t_L g2604 ( 
.A(n_2158),
.Y(n_2604)
);

BUFx3_ASAP7_75t_L g2605 ( 
.A(n_2169),
.Y(n_2605)
);

INVx2_ASAP7_75t_SL g2606 ( 
.A(n_2176),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2199),
.B(n_104),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_1989),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2206),
.B(n_105),
.Y(n_2609)
);

AOI22xp5_ASAP7_75t_L g2610 ( 
.A1(n_2194),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_1952),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2054),
.B(n_106),
.Y(n_2612)
);

NOR2xp33_ASAP7_75t_L g2613 ( 
.A(n_2217),
.B(n_107),
.Y(n_2613)
);

OR2x2_ASAP7_75t_L g2614 ( 
.A(n_2179),
.B(n_108),
.Y(n_2614)
);

AOI22xp5_ASAP7_75t_L g2615 ( 
.A1(n_2195),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_2615)
);

INVx2_ASAP7_75t_SL g2616 ( 
.A(n_2158),
.Y(n_2616)
);

HB1xp67_ASAP7_75t_L g2617 ( 
.A(n_2222),
.Y(n_2617)
);

O2A1O1Ixp33_ASAP7_75t_L g2618 ( 
.A1(n_2056),
.A2(n_112),
.B(n_110),
.C(n_111),
.Y(n_2618)
);

OAI22xp5_ASAP7_75t_SL g2619 ( 
.A1(n_2212),
.A2(n_115),
.B1(n_111),
.B2(n_114),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2192),
.B(n_2193),
.Y(n_2620)
);

OR2x2_ASAP7_75t_SL g2621 ( 
.A(n_2230),
.B(n_116),
.Y(n_2621)
);

INVx3_ASAP7_75t_L g2622 ( 
.A(n_2249),
.Y(n_2622)
);

BUFx2_ASAP7_75t_L g2623 ( 
.A(n_2131),
.Y(n_2623)
);

BUFx2_ASAP7_75t_L g2624 ( 
.A(n_2131),
.Y(n_2624)
);

INVxp67_ASAP7_75t_L g2625 ( 
.A(n_2250),
.Y(n_2625)
);

INVx3_ASAP7_75t_L g2626 ( 
.A(n_2031),
.Y(n_2626)
);

AOI22xp33_ASAP7_75t_L g2627 ( 
.A1(n_2195),
.A2(n_2071),
.B1(n_1965),
.B2(n_1971),
.Y(n_2627)
);

BUFx6f_ASAP7_75t_L g2628 ( 
.A(n_2031),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2064),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2083),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_1957),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2097),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2132),
.Y(n_2633)
);

NOR2xp33_ASAP7_75t_L g2634 ( 
.A(n_2232),
.B(n_116),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2071),
.B(n_117),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2095),
.Y(n_2636)
);

INVx4_ASAP7_75t_L g2637 ( 
.A(n_2222),
.Y(n_2637)
);

BUFx8_ASAP7_75t_L g2638 ( 
.A(n_2131),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2136),
.Y(n_2639)
);

AOI22xp33_ASAP7_75t_L g2640 ( 
.A1(n_1981),
.A2(n_121),
.B1(n_118),
.B2(n_119),
.Y(n_2640)
);

O2A1O1Ixp5_ASAP7_75t_L g2641 ( 
.A1(n_1960),
.A2(n_633),
.B(n_634),
.C(n_632),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2178),
.Y(n_2642)
);

OR2x6_ASAP7_75t_L g2643 ( 
.A(n_2053),
.B(n_118),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2198),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2203),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2204),
.Y(n_2646)
);

AOI22xp33_ASAP7_75t_L g2647 ( 
.A1(n_1919),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_2647)
);

OAI21xp33_ASAP7_75t_L g2648 ( 
.A1(n_1933),
.A2(n_122),
.B(n_123),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2205),
.Y(n_2649)
);

HB1xp67_ASAP7_75t_L g2650 ( 
.A(n_2248),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_1931),
.B(n_124),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_SL g2652 ( 
.A(n_2053),
.B(n_125),
.Y(n_2652)
);

AOI21x1_ASAP7_75t_L g2653 ( 
.A1(n_2248),
.A2(n_638),
.B(n_637),
.Y(n_2653)
);

INVxp67_ASAP7_75t_L g2654 ( 
.A(n_2133),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_1934),
.B(n_126),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2211),
.Y(n_2656)
);

INVx5_ASAP7_75t_L g2657 ( 
.A(n_2133),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2213),
.Y(n_2658)
);

INVx5_ASAP7_75t_L g2659 ( 
.A(n_2133),
.Y(n_2659)
);

INVx2_ASAP7_75t_SL g2660 ( 
.A(n_2252),
.Y(n_2660)
);

BUFx6f_ASAP7_75t_L g2661 ( 
.A(n_2066),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2066),
.B(n_127),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2225),
.B(n_127),
.Y(n_2663)
);

AND3x2_ASAP7_75t_SL g2664 ( 
.A(n_2018),
.B(n_128),
.C(n_129),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2019),
.B(n_130),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2022),
.B(n_131),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2246),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2252),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_SL g2669 ( 
.A(n_2140),
.B(n_134),
.Y(n_2669)
);

NAND2xp33_ASAP7_75t_L g2670 ( 
.A(n_2140),
.B(n_640),
.Y(n_2670)
);

NOR2xp33_ASAP7_75t_L g2671 ( 
.A(n_2244),
.B(n_2172),
.Y(n_2671)
);

BUFx3_ASAP7_75t_L g2672 ( 
.A(n_2172),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_1933),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2244),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_SL g2675 ( 
.A(n_2183),
.B(n_134),
.Y(n_2675)
);

AND2x2_ASAP7_75t_L g2676 ( 
.A(n_2183),
.B(n_135),
.Y(n_2676)
);

INVx3_ASAP7_75t_L g2677 ( 
.A(n_1977),
.Y(n_2677)
);

NAND2x1p5_ASAP7_75t_L g2678 ( 
.A(n_1929),
.B(n_138),
.Y(n_2678)
);

OAI22xp5_ASAP7_75t_SL g2679 ( 
.A1(n_1943),
.A2(n_141),
.B1(n_137),
.B2(n_140),
.Y(n_2679)
);

BUFx6f_ASAP7_75t_L g2680 ( 
.A(n_2247),
.Y(n_2680)
);

NOR2xp33_ASAP7_75t_L g2681 ( 
.A(n_1906),
.B(n_142),
.Y(n_2681)
);

INVxp67_ASAP7_75t_L g2682 ( 
.A(n_1907),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_1909),
.Y(n_2683)
);

BUFx3_ASAP7_75t_L g2684 ( 
.A(n_1932),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2161),
.B(n_142),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2161),
.B(n_143),
.Y(n_2686)
);

INVx4_ASAP7_75t_L g2687 ( 
.A(n_1929),
.Y(n_2687)
);

AOI22xp33_ASAP7_75t_L g2688 ( 
.A1(n_1949),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_2688)
);

BUFx6f_ASAP7_75t_L g2689 ( 
.A(n_2247),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_1909),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2161),
.B(n_144),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_1907),
.B(n_145),
.Y(n_2692)
);

NOR3xp33_ASAP7_75t_SL g2693 ( 
.A(n_1959),
.B(n_147),
.C(n_148),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_1909),
.Y(n_2694)
);

AOI22xp5_ASAP7_75t_L g2695 ( 
.A1(n_2229),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2161),
.B(n_149),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2161),
.B(n_151),
.Y(n_2697)
);

NOR2xp33_ASAP7_75t_L g2698 ( 
.A(n_1906),
.B(n_152),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_1909),
.Y(n_2699)
);

NOR2xp33_ASAP7_75t_R g2700 ( 
.A(n_1993),
.B(n_153),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_1909),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_1909),
.Y(n_2702)
);

AND2x4_ASAP7_75t_L g2703 ( 
.A(n_1907),
.B(n_153),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_1909),
.Y(n_2704)
);

CKINVDCx5p33_ASAP7_75t_R g2705 ( 
.A(n_1959),
.Y(n_2705)
);

AND2x4_ASAP7_75t_L g2706 ( 
.A(n_1907),
.B(n_154),
.Y(n_2706)
);

A2O1A1Ixp33_ASAP7_75t_L g2707 ( 
.A1(n_2197),
.A2(n_156),
.B(n_154),
.C(n_155),
.Y(n_2707)
);

BUFx8_ASAP7_75t_L g2708 ( 
.A(n_1928),
.Y(n_2708)
);

INVx5_ASAP7_75t_L g2709 ( 
.A(n_2033),
.Y(n_2709)
);

INVx4_ASAP7_75t_L g2710 ( 
.A(n_1929),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_1909),
.Y(n_2711)
);

INVx3_ASAP7_75t_L g2712 ( 
.A(n_1977),
.Y(n_2712)
);

INVx5_ASAP7_75t_L g2713 ( 
.A(n_2033),
.Y(n_2713)
);

INVx3_ASAP7_75t_SL g2714 ( 
.A(n_1959),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_1909),
.Y(n_2715)
);

INVx2_ASAP7_75t_SL g2716 ( 
.A(n_1932),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2161),
.B(n_155),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2161),
.B(n_156),
.Y(n_2718)
);

AOI22xp5_ASAP7_75t_L g2719 ( 
.A1(n_2229),
.A2(n_160),
.B1(n_157),
.B2(n_158),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_1909),
.Y(n_2720)
);

NOR3xp33_ASAP7_75t_SL g2721 ( 
.A(n_1959),
.B(n_157),
.C(n_158),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_1909),
.Y(n_2722)
);

AOI21xp5_ASAP7_75t_L g2723 ( 
.A1(n_1927),
.A2(n_642),
.B(n_641),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2356),
.B(n_160),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2263),
.Y(n_2725)
);

INVx4_ASAP7_75t_L g2726 ( 
.A(n_2288),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2339),
.Y(n_2727)
);

AOI22xp5_ASAP7_75t_L g2728 ( 
.A1(n_2561),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_2728)
);

A2O1A1Ixp33_ASAP7_75t_L g2729 ( 
.A1(n_2509),
.A2(n_2578),
.B(n_2466),
.C(n_2634),
.Y(n_2729)
);

BUFx3_ASAP7_75t_L g2730 ( 
.A(n_2708),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2330),
.B(n_164),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2341),
.Y(n_2732)
);

NOR2xp33_ASAP7_75t_L g2733 ( 
.A(n_2585),
.B(n_165),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2361),
.Y(n_2734)
);

AND2x2_ASAP7_75t_L g2735 ( 
.A(n_2283),
.B(n_165),
.Y(n_2735)
);

AOI22xp33_ASAP7_75t_L g2736 ( 
.A1(n_2424),
.A2(n_2351),
.B1(n_2679),
.B2(n_2387),
.Y(n_2736)
);

BUFx2_ASAP7_75t_L g2737 ( 
.A(n_2708),
.Y(n_2737)
);

CKINVDCx5p33_ASAP7_75t_R g2738 ( 
.A(n_2312),
.Y(n_2738)
);

NOR2xp33_ASAP7_75t_L g2739 ( 
.A(n_2570),
.B(n_166),
.Y(n_2739)
);

AND2x4_ASAP7_75t_L g2740 ( 
.A(n_2385),
.B(n_166),
.Y(n_2740)
);

INVx4_ASAP7_75t_L g2741 ( 
.A(n_2288),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2394),
.B(n_2465),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2534),
.B(n_167),
.Y(n_2743)
);

INVx4_ASAP7_75t_L g2744 ( 
.A(n_2288),
.Y(n_2744)
);

CKINVDCx5p33_ASAP7_75t_R g2745 ( 
.A(n_2705),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2400),
.B(n_167),
.Y(n_2746)
);

AOI21xp5_ASAP7_75t_L g2747 ( 
.A1(n_2620),
.A2(n_646),
.B(n_645),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2267),
.Y(n_2748)
);

INVx3_ASAP7_75t_L g2749 ( 
.A(n_2637),
.Y(n_2749)
);

CKINVDCx5p33_ASAP7_75t_R g2750 ( 
.A(n_2306),
.Y(n_2750)
);

BUFx2_ASAP7_75t_L g2751 ( 
.A(n_2297),
.Y(n_2751)
);

BUFx6f_ASAP7_75t_L g2752 ( 
.A(n_2311),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2273),
.Y(n_2753)
);

INVxp67_ASAP7_75t_SL g2754 ( 
.A(n_2551),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2272),
.B(n_168),
.Y(n_2755)
);

HB1xp67_ASAP7_75t_L g2756 ( 
.A(n_2255),
.Y(n_2756)
);

INVx6_ASAP7_75t_L g2757 ( 
.A(n_2563),
.Y(n_2757)
);

INVx1_ASAP7_75t_SL g2758 ( 
.A(n_2438),
.Y(n_2758)
);

AND2x2_ASAP7_75t_L g2759 ( 
.A(n_2581),
.B(n_169),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2276),
.Y(n_2760)
);

AND2x4_ASAP7_75t_SL g2761 ( 
.A(n_2385),
.B(n_169),
.Y(n_2761)
);

BUFx8_ASAP7_75t_L g2762 ( 
.A(n_2495),
.Y(n_2762)
);

INVx1_ASAP7_75t_SL g2763 ( 
.A(n_2275),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2272),
.B(n_2331),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2301),
.Y(n_2765)
);

BUFx6f_ASAP7_75t_L g2766 ( 
.A(n_2311),
.Y(n_2766)
);

OR2x2_ASAP7_75t_L g2767 ( 
.A(n_2300),
.B(n_170),
.Y(n_2767)
);

INVx1_ASAP7_75t_SL g2768 ( 
.A(n_2262),
.Y(n_2768)
);

BUFx2_ASAP7_75t_L g2769 ( 
.A(n_2551),
.Y(n_2769)
);

AOI22xp5_ASAP7_75t_L g2770 ( 
.A1(n_2424),
.A2(n_2331),
.B1(n_2323),
.B2(n_2537),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2326),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2581),
.B(n_170),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2542),
.B(n_171),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2266),
.B(n_171),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2268),
.B(n_2282),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2701),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2711),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2722),
.Y(n_2778)
);

HB1xp67_ASAP7_75t_L g2779 ( 
.A(n_2261),
.Y(n_2779)
);

NOR2x1_ASAP7_75t_L g2780 ( 
.A(n_2687),
.B(n_172),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2293),
.B(n_172),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2348),
.Y(n_2782)
);

BUFx2_ASAP7_75t_L g2783 ( 
.A(n_2554),
.Y(n_2783)
);

INVx3_ASAP7_75t_L g2784 ( 
.A(n_2637),
.Y(n_2784)
);

AND2x4_ASAP7_75t_L g2785 ( 
.A(n_2304),
.B(n_174),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2302),
.B(n_174),
.Y(n_2786)
);

BUFx6f_ASAP7_75t_L g2787 ( 
.A(n_2311),
.Y(n_2787)
);

OR2x2_ASAP7_75t_L g2788 ( 
.A(n_2523),
.B(n_175),
.Y(n_2788)
);

OAI22xp5_ASAP7_75t_L g2789 ( 
.A1(n_2695),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2362),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2318),
.B(n_2321),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2555),
.Y(n_2792)
);

INVx1_ASAP7_75t_SL g2793 ( 
.A(n_2490),
.Y(n_2793)
);

INVx3_ASAP7_75t_L g2794 ( 
.A(n_2313),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2572),
.Y(n_2795)
);

AND2x2_ASAP7_75t_L g2796 ( 
.A(n_2506),
.B(n_176),
.Y(n_2796)
);

OAI21xp5_ASAP7_75t_L g2797 ( 
.A1(n_2292),
.A2(n_177),
.B(n_178),
.Y(n_2797)
);

OAI22xp5_ASAP7_75t_L g2798 ( 
.A1(n_2695),
.A2(n_2719),
.B1(n_2367),
.B2(n_2324),
.Y(n_2798)
);

BUFx3_ASAP7_75t_L g2799 ( 
.A(n_2684),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2333),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2337),
.B(n_178),
.Y(n_2801)
);

NOR2xp33_ASAP7_75t_L g2802 ( 
.A(n_2552),
.B(n_2459),
.Y(n_2802)
);

NOR2xp33_ASAP7_75t_R g2803 ( 
.A(n_2436),
.B(n_179),
.Y(n_2803)
);

NOR2xp33_ASAP7_75t_R g2804 ( 
.A(n_2270),
.B(n_179),
.Y(n_2804)
);

AND2x4_ASAP7_75t_L g2805 ( 
.A(n_2304),
.B(n_181),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2583),
.Y(n_2806)
);

HB1xp67_ASAP7_75t_L g2807 ( 
.A(n_2278),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2586),
.Y(n_2808)
);

NAND2x1p5_ASAP7_75t_L g2809 ( 
.A(n_2304),
.B(n_181),
.Y(n_2809)
);

NOR2xp33_ASAP7_75t_L g2810 ( 
.A(n_2533),
.B(n_184),
.Y(n_2810)
);

CKINVDCx20_ASAP7_75t_R g2811 ( 
.A(n_2700),
.Y(n_2811)
);

CKINVDCx11_ASAP7_75t_R g2812 ( 
.A(n_2714),
.Y(n_2812)
);

HB1xp67_ASAP7_75t_L g2813 ( 
.A(n_2643),
.Y(n_2813)
);

OR2x2_ASAP7_75t_L g2814 ( 
.A(n_2454),
.B(n_184),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2375),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2338),
.B(n_185),
.Y(n_2816)
);

NOR2xp67_ASAP7_75t_SL g2817 ( 
.A(n_2709),
.B(n_2713),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2683),
.Y(n_2818)
);

NOR2xp33_ASAP7_75t_L g2819 ( 
.A(n_2625),
.B(n_185),
.Y(n_2819)
);

OAI22xp5_ASAP7_75t_SL g2820 ( 
.A1(n_2281),
.A2(n_2387),
.B1(n_2679),
.B2(n_2393),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2363),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2365),
.Y(n_2822)
);

NAND3xp33_ASAP7_75t_SL g2823 ( 
.A(n_2406),
.B(n_186),
.C(n_188),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2690),
.B(n_189),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2694),
.B(n_189),
.Y(n_2825)
);

NOR2xp33_ASAP7_75t_L g2826 ( 
.A(n_2580),
.B(n_2522),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2378),
.Y(n_2827)
);

AND2x4_ASAP7_75t_L g2828 ( 
.A(n_2709),
.B(n_190),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2370),
.Y(n_2829)
);

HB1xp67_ASAP7_75t_L g2830 ( 
.A(n_2643),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2699),
.Y(n_2831)
);

AND2x2_ASAP7_75t_SL g2832 ( 
.A(n_2589),
.B(n_191),
.Y(n_2832)
);

NAND2xp33_ASAP7_75t_SL g2833 ( 
.A(n_2566),
.B(n_191),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2702),
.B(n_193),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2704),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2715),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2382),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2720),
.B(n_194),
.Y(n_2838)
);

INVx3_ASAP7_75t_SL g2839 ( 
.A(n_2599),
.Y(n_2839)
);

INVx3_ASAP7_75t_L g2840 ( 
.A(n_2313),
.Y(n_2840)
);

BUFx2_ASAP7_75t_L g2841 ( 
.A(n_2554),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2547),
.B(n_194),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2409),
.B(n_195),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2413),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2416),
.Y(n_2845)
);

AOI221xp5_ASAP7_75t_L g2846 ( 
.A1(n_2359),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.C(n_198),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2575),
.B(n_196),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2419),
.B(n_199),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2420),
.B(n_200),
.Y(n_2849)
);

AND2x4_ASAP7_75t_L g2850 ( 
.A(n_2709),
.B(n_201),
.Y(n_2850)
);

INVx4_ASAP7_75t_L g2851 ( 
.A(n_2713),
.Y(n_2851)
);

BUFx8_ASAP7_75t_L g2852 ( 
.A(n_2495),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2425),
.B(n_201),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2386),
.Y(n_2854)
);

AND3x1_ASAP7_75t_L g2855 ( 
.A(n_2693),
.B(n_202),
.C(n_203),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2430),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2437),
.B(n_202),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2399),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2440),
.B(n_203),
.Y(n_2859)
);

AND2x4_ASAP7_75t_L g2860 ( 
.A(n_2713),
.B(n_2563),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2441),
.B(n_204),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2455),
.Y(n_2862)
);

OR2x6_ASAP7_75t_L g2863 ( 
.A(n_2687),
.B(n_204),
.Y(n_2863)
);

OAI22xp5_ASAP7_75t_L g2864 ( 
.A1(n_2719),
.A2(n_208),
.B1(n_205),
.B2(n_207),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2462),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2354),
.B(n_205),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2404),
.Y(n_2867)
);

HB1xp67_ASAP7_75t_L g2868 ( 
.A(n_2643),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2405),
.Y(n_2869)
);

BUFx2_ASAP7_75t_L g2870 ( 
.A(n_2355),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2371),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2451),
.B(n_207),
.Y(n_2872)
);

INVxp67_ASAP7_75t_L g2873 ( 
.A(n_2259),
.Y(n_2873)
);

BUFx6f_ASAP7_75t_L g2874 ( 
.A(n_2345),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2415),
.Y(n_2875)
);

AOI22xp5_ASAP7_75t_L g2876 ( 
.A1(n_2270),
.A2(n_2305),
.B1(n_2332),
.B2(n_2613),
.Y(n_2876)
);

INVx2_ASAP7_75t_SL g2877 ( 
.A(n_2474),
.Y(n_2877)
);

AOI22xp5_ASAP7_75t_L g2878 ( 
.A1(n_2414),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2381),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2442),
.B(n_210),
.Y(n_2880)
);

INVx2_ASAP7_75t_SL g2881 ( 
.A(n_2474),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_SL g2882 ( 
.A(n_2450),
.B(n_211),
.Y(n_2882)
);

OR2x2_ASAP7_75t_SL g2883 ( 
.A(n_2422),
.B(n_211),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2518),
.B(n_2503),
.Y(n_2884)
);

INVxp67_ASAP7_75t_SL g2885 ( 
.A(n_2604),
.Y(n_2885)
);

OR2x2_ASAP7_75t_L g2886 ( 
.A(n_2374),
.B(n_212),
.Y(n_2886)
);

INVx2_ASAP7_75t_SL g2887 ( 
.A(n_2474),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2391),
.B(n_212),
.Y(n_2888)
);

BUFx2_ASAP7_75t_L g2889 ( 
.A(n_2604),
.Y(n_2889)
);

INVx3_ASAP7_75t_L g2890 ( 
.A(n_2344),
.Y(n_2890)
);

HB1xp67_ASAP7_75t_L g2891 ( 
.A(n_2504),
.Y(n_2891)
);

AOI21xp5_ASAP7_75t_L g2892 ( 
.A1(n_2673),
.A2(n_649),
.B(n_647),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2397),
.B(n_213),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2463),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2468),
.Y(n_2895)
);

NOR2xp33_ASAP7_75t_L g2896 ( 
.A(n_2287),
.B(n_213),
.Y(n_2896)
);

INVx2_ASAP7_75t_SL g2897 ( 
.A(n_2479),
.Y(n_2897)
);

BUFx6f_ASAP7_75t_L g2898 ( 
.A(n_2345),
.Y(n_2898)
);

BUFx3_ASAP7_75t_L g2899 ( 
.A(n_2392),
.Y(n_2899)
);

NOR2xp33_ASAP7_75t_L g2900 ( 
.A(n_2372),
.B(n_214),
.Y(n_2900)
);

INVx3_ASAP7_75t_SL g2901 ( 
.A(n_2710),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2417),
.Y(n_2902)
);

BUFx6f_ASAP7_75t_L g2903 ( 
.A(n_2345),
.Y(n_2903)
);

BUFx3_ASAP7_75t_L g2904 ( 
.A(n_2342),
.Y(n_2904)
);

NOR2xp33_ASAP7_75t_L g2905 ( 
.A(n_2335),
.B(n_214),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2429),
.B(n_215),
.Y(n_2906)
);

BUFx6f_ASAP7_75t_L g2907 ( 
.A(n_2401),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2510),
.B(n_215),
.Y(n_2908)
);

AND2x2_ASAP7_75t_L g2909 ( 
.A(n_2562),
.B(n_216),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2469),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2428),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2519),
.B(n_2294),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2346),
.Y(n_2913)
);

INVx3_ASAP7_75t_L g2914 ( 
.A(n_2344),
.Y(n_2914)
);

BUFx3_ASAP7_75t_L g2915 ( 
.A(n_2310),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2473),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2384),
.B(n_216),
.Y(n_2917)
);

INVx4_ASAP7_75t_L g2918 ( 
.A(n_2479),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2369),
.Y(n_2919)
);

A2O1A1Ixp33_ASAP7_75t_L g2920 ( 
.A1(n_2681),
.A2(n_220),
.B(n_217),
.C(n_219),
.Y(n_2920)
);

BUFx3_ASAP7_75t_L g2921 ( 
.A(n_2314),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2477),
.Y(n_2922)
);

NAND2xp33_ASAP7_75t_L g2923 ( 
.A(n_2349),
.B(n_2577),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2480),
.B(n_220),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2481),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2482),
.Y(n_2926)
);

AO22x1_ASAP7_75t_L g2927 ( 
.A1(n_2638),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2484),
.B(n_222),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2493),
.Y(n_2929)
);

BUFx5_ASAP7_75t_L g2930 ( 
.A(n_2349),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_2303),
.B(n_223),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2494),
.Y(n_2932)
);

AOI22xp5_ASAP7_75t_L g2933 ( 
.A1(n_2414),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_2933)
);

INVx2_ASAP7_75t_SL g2934 ( 
.A(n_2479),
.Y(n_2934)
);

BUFx6f_ASAP7_75t_L g2935 ( 
.A(n_2401),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2497),
.Y(n_2936)
);

AOI22xp5_ASAP7_75t_L g2937 ( 
.A1(n_2431),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_2937)
);

BUFx3_ASAP7_75t_L g2938 ( 
.A(n_2319),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2501),
.B(n_227),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2507),
.Y(n_2940)
);

A2O1A1Ixp33_ASAP7_75t_L g2941 ( 
.A1(n_2698),
.A2(n_2594),
.B(n_2590),
.C(n_2396),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2508),
.B(n_228),
.Y(n_2942)
);

OAI22xp5_ASAP7_75t_L g2943 ( 
.A1(n_2485),
.A2(n_231),
.B1(n_228),
.B2(n_229),
.Y(n_2943)
);

AO221x1_ASAP7_75t_L g2944 ( 
.A1(n_2464),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.C(n_235),
.Y(n_2944)
);

BUFx6f_ASAP7_75t_L g2945 ( 
.A(n_2401),
.Y(n_2945)
);

AOI22xp33_ASAP7_75t_L g2946 ( 
.A1(n_2562),
.A2(n_236),
.B1(n_233),
.B2(n_235),
.Y(n_2946)
);

NOR2x1_ASAP7_75t_L g2947 ( 
.A(n_2710),
.B(n_237),
.Y(n_2947)
);

INVx4_ASAP7_75t_L g2948 ( 
.A(n_2577),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2540),
.Y(n_2949)
);

HB1xp67_ASAP7_75t_L g2950 ( 
.A(n_2504),
.Y(n_2950)
);

CKINVDCx11_ASAP7_75t_R g2951 ( 
.A(n_2411),
.Y(n_2951)
);

O2A1O1Ixp33_ASAP7_75t_L g2952 ( 
.A1(n_2514),
.A2(n_2520),
.B(n_2532),
.C(n_2553),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_L g2953 ( 
.A(n_2258),
.B(n_237),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2260),
.B(n_2277),
.Y(n_2954)
);

INVx3_ASAP7_75t_L g2955 ( 
.A(n_2377),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2279),
.B(n_238),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2541),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2524),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2526),
.Y(n_2959)
);

AOI22xp5_ASAP7_75t_L g2960 ( 
.A1(n_2431),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_2960)
);

INVx2_ASAP7_75t_SL g2961 ( 
.A(n_2565),
.Y(n_2961)
);

O2A1O1Ixp33_ASAP7_75t_L g2962 ( 
.A1(n_2607),
.A2(n_242),
.B(n_239),
.C(n_240),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2535),
.Y(n_2963)
);

BUFx6f_ASAP7_75t_L g2964 ( 
.A(n_2527),
.Y(n_2964)
);

AND3x1_ASAP7_75t_SL g2965 ( 
.A(n_2373),
.B(n_243),
.C(n_244),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2284),
.B(n_243),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2703),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2285),
.B(n_244),
.Y(n_2968)
);

AND2x4_ASAP7_75t_L g2969 ( 
.A(n_2377),
.B(n_245),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2286),
.B(n_2291),
.Y(n_2970)
);

AOI22xp33_ASAP7_75t_L g2971 ( 
.A1(n_2562),
.A2(n_247),
.B1(n_245),
.B2(n_246),
.Y(n_2971)
);

AOI22xp5_ASAP7_75t_L g2972 ( 
.A1(n_2582),
.A2(n_250),
.B1(n_247),
.B2(n_249),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_SL g2973 ( 
.A(n_2336),
.B(n_251),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2703),
.Y(n_2974)
);

BUFx3_ASAP7_75t_L g2975 ( 
.A(n_2325),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2706),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_SL g2977 ( 
.A(n_2336),
.B(n_252),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2458),
.Y(n_2978)
);

INVx2_ASAP7_75t_SL g2979 ( 
.A(n_2565),
.Y(n_2979)
);

BUFx4f_ASAP7_75t_L g2980 ( 
.A(n_2295),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2470),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2340),
.B(n_253),
.Y(n_2982)
);

A2O1A1Ixp33_ASAP7_75t_L g2983 ( 
.A1(n_2588),
.A2(n_255),
.B(n_253),
.C(n_254),
.Y(n_2983)
);

NOR2xp33_ASAP7_75t_SL g2984 ( 
.A(n_2638),
.B(n_254),
.Y(n_2984)
);

AND2x4_ASAP7_75t_L g2985 ( 
.A(n_2677),
.B(n_255),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_SL g2986 ( 
.A(n_2352),
.B(n_256),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2706),
.Y(n_2987)
);

INVxp67_ASAP7_75t_SL g2988 ( 
.A(n_2589),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2569),
.B(n_256),
.Y(n_2989)
);

INVx4_ASAP7_75t_L g2990 ( 
.A(n_2577),
.Y(n_2990)
);

INVx1_ASAP7_75t_SL g2991 ( 
.A(n_2446),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2685),
.Y(n_2992)
);

OR2x2_ASAP7_75t_L g2993 ( 
.A(n_2315),
.B(n_257),
.Y(n_2993)
);

INVx1_ASAP7_75t_SL g2994 ( 
.A(n_2352),
.Y(n_2994)
);

CKINVDCx5p33_ASAP7_75t_R g2995 ( 
.A(n_2388),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2513),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2614),
.B(n_257),
.Y(n_2997)
);

AOI22xp33_ASAP7_75t_L g2998 ( 
.A1(n_2600),
.A2(n_2445),
.B1(n_2598),
.B2(n_2483),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2274),
.B(n_259),
.Y(n_2999)
);

NOR2xp33_ASAP7_75t_L g3000 ( 
.A(n_2303),
.B(n_259),
.Y(n_3000)
);

BUFx2_ASAP7_75t_L g3001 ( 
.A(n_2574),
.Y(n_3001)
);

INVx4_ASAP7_75t_L g3002 ( 
.A(n_2403),
.Y(n_3002)
);

AND2x4_ASAP7_75t_L g3003 ( 
.A(n_2677),
.B(n_260),
.Y(n_3003)
);

NAND3xp33_ASAP7_75t_SL g3004 ( 
.A(n_2406),
.B(n_260),
.C(n_261),
.Y(n_3004)
);

BUFx12f_ASAP7_75t_L g3005 ( 
.A(n_2388),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2686),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2691),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2696),
.Y(n_3008)
);

BUFx6f_ASAP7_75t_L g3009 ( 
.A(n_2527),
.Y(n_3009)
);

INVx3_ASAP7_75t_L g3010 ( 
.A(n_2712),
.Y(n_3010)
);

INVx3_ASAP7_75t_L g3011 ( 
.A(n_2712),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2558),
.B(n_261),
.Y(n_3012)
);

HB1xp67_ASAP7_75t_L g3013 ( 
.A(n_2559),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2498),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2697),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2545),
.B(n_262),
.Y(n_3016)
);

BUFx12f_ASAP7_75t_L g3017 ( 
.A(n_2257),
.Y(n_3017)
);

HB1xp67_ASAP7_75t_L g3018 ( 
.A(n_2559),
.Y(n_3018)
);

HB1xp67_ASAP7_75t_L g3019 ( 
.A(n_2559),
.Y(n_3019)
);

INVx3_ASAP7_75t_L g3020 ( 
.A(n_2605),
.Y(n_3020)
);

AND2x4_ASAP7_75t_L g3021 ( 
.A(n_2412),
.B(n_262),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2682),
.B(n_264),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2307),
.B(n_264),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2317),
.B(n_266),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2717),
.Y(n_3025)
);

BUFx2_ASAP7_75t_L g3026 ( 
.A(n_2574),
.Y(n_3026)
);

BUFx3_ASAP7_75t_L g3027 ( 
.A(n_2265),
.Y(n_3027)
);

NOR2xp33_ASAP7_75t_L g3028 ( 
.A(n_2289),
.B(n_266),
.Y(n_3028)
);

OR2x6_ASAP7_75t_L g3029 ( 
.A(n_2511),
.B(n_267),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2500),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2718),
.Y(n_3031)
);

INVxp67_ASAP7_75t_L g3032 ( 
.A(n_2426),
.Y(n_3032)
);

NOR3xp33_ASAP7_75t_L g3033 ( 
.A(n_2619),
.B(n_267),
.C(n_268),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2608),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2491),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2256),
.B(n_268),
.Y(n_3036)
);

AND2x2_ASAP7_75t_L g3037 ( 
.A(n_2550),
.B(n_270),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_2645),
.Y(n_3038)
);

INVx2_ASAP7_75t_SL g3039 ( 
.A(n_2716),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2491),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2353),
.Y(n_3041)
);

INVx3_ASAP7_75t_L g3042 ( 
.A(n_2412),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2327),
.B(n_270),
.Y(n_3043)
);

OAI22xp5_ASAP7_75t_L g3044 ( 
.A1(n_2485),
.A2(n_273),
.B1(n_271),
.B2(n_272),
.Y(n_3044)
);

INVx3_ASAP7_75t_L g3045 ( 
.A(n_2439),
.Y(n_3045)
);

AND2x4_ASAP7_75t_L g3046 ( 
.A(n_2439),
.B(n_271),
.Y(n_3046)
);

INVx3_ASAP7_75t_L g3047 ( 
.A(n_2423),
.Y(n_3047)
);

INVx5_ASAP7_75t_L g3048 ( 
.A(n_2349),
.Y(n_3048)
);

CKINVDCx5p33_ASAP7_75t_R g3049 ( 
.A(n_2531),
.Y(n_3049)
);

BUFx3_ASAP7_75t_L g3050 ( 
.A(n_2543),
.Y(n_3050)
);

INVx2_ASAP7_75t_L g3051 ( 
.A(n_2646),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_SL g3052 ( 
.A(n_2334),
.B(n_272),
.Y(n_3052)
);

INVx2_ASAP7_75t_SL g3053 ( 
.A(n_2487),
.Y(n_3053)
);

NOR2xp33_ASAP7_75t_L g3054 ( 
.A(n_2322),
.B(n_275),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_L g3055 ( 
.A(n_2525),
.B(n_275),
.Y(n_3055)
);

AND2x6_ASAP7_75t_L g3056 ( 
.A(n_2280),
.B(n_276),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2692),
.Y(n_3057)
);

INVx3_ASAP7_75t_L g3058 ( 
.A(n_2423),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2557),
.Y(n_3059)
);

AOI22xp5_ASAP7_75t_L g3060 ( 
.A1(n_2600),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2557),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2499),
.Y(n_3062)
);

BUFx2_ASAP7_75t_L g3063 ( 
.A(n_2432),
.Y(n_3063)
);

AOI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_2598),
.A2(n_281),
.B1(n_277),
.B2(n_280),
.Y(n_3064)
);

BUFx3_ASAP7_75t_L g3065 ( 
.A(n_2309),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2656),
.Y(n_3066)
);

AND2x2_ASAP7_75t_L g3067 ( 
.A(n_2373),
.B(n_280),
.Y(n_3067)
);

INVx3_ASAP7_75t_L g3068 ( 
.A(n_2443),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2644),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2649),
.Y(n_3070)
);

AND2x2_ASAP7_75t_L g3071 ( 
.A(n_2408),
.B(n_2271),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2549),
.B(n_282),
.Y(n_3072)
);

INVx5_ASAP7_75t_L g3073 ( 
.A(n_2349),
.Y(n_3073)
);

INVx3_ASAP7_75t_L g3074 ( 
.A(n_2443),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2564),
.B(n_282),
.Y(n_3075)
);

BUFx6f_ASAP7_75t_L g3076 ( 
.A(n_2527),
.Y(n_3076)
);

XNOR2x1_ASAP7_75t_L g3077 ( 
.A(n_2678),
.B(n_283),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2658),
.Y(n_3078)
);

INVx4_ASAP7_75t_L g3079 ( 
.A(n_2529),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2667),
.Y(n_3080)
);

AOI22xp5_ASAP7_75t_L g3081 ( 
.A1(n_2334),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_2476),
.Y(n_3082)
);

AOI22xp33_ASAP7_75t_L g3083 ( 
.A1(n_2464),
.A2(n_287),
.B1(n_284),
.B2(n_286),
.Y(n_3083)
);

HB1xp67_ASAP7_75t_L g3084 ( 
.A(n_2544),
.Y(n_3084)
);

NOR2xp33_ASAP7_75t_L g3085 ( 
.A(n_2299),
.B(n_287),
.Y(n_3085)
);

NOR2xp33_ASAP7_75t_L g3086 ( 
.A(n_2308),
.B(n_288),
.Y(n_3086)
);

CKINVDCx6p67_ASAP7_75t_R g3087 ( 
.A(n_2432),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2571),
.B(n_289),
.Y(n_3088)
);

OR2x2_ASAP7_75t_L g3089 ( 
.A(n_2407),
.B(n_289),
.Y(n_3089)
);

OR2x6_ASAP7_75t_L g3090 ( 
.A(n_2478),
.B(n_290),
.Y(n_3090)
);

CKINVDCx11_ASAP7_75t_R g3091 ( 
.A(n_2478),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2579),
.B(n_290),
.Y(n_3092)
);

INVx1_ASAP7_75t_SL g3093 ( 
.A(n_2591),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2410),
.B(n_291),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2418),
.B(n_291),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2427),
.Y(n_3096)
);

AOI22xp33_ASAP7_75t_L g3097 ( 
.A1(n_2556),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2398),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2603),
.Y(n_3099)
);

AOI22xp33_ASAP7_75t_L g3100 ( 
.A1(n_2619),
.A2(n_295),
.B1(n_292),
.B2(n_294),
.Y(n_3100)
);

INVx1_ASAP7_75t_SL g3101 ( 
.A(n_2505),
.Y(n_3101)
);

AOI221xp5_ASAP7_75t_SL g3102 ( 
.A1(n_2592),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.C(n_299),
.Y(n_3102)
);

AOI22xp5_ASAP7_75t_L g3103 ( 
.A1(n_2456),
.A2(n_299),
.B1(n_296),
.B2(n_297),
.Y(n_3103)
);

INVx2_ASAP7_75t_L g3104 ( 
.A(n_2488),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2663),
.Y(n_3105)
);

AOI22xp5_ASAP7_75t_L g3106 ( 
.A1(n_2471),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2536),
.Y(n_3107)
);

INVxp67_ASAP7_75t_L g3108 ( 
.A(n_2366),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2597),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2611),
.Y(n_3110)
);

AND2x2_ASAP7_75t_L g3111 ( 
.A(n_2408),
.B(n_2539),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2447),
.B(n_301),
.Y(n_3112)
);

INVxp67_ASAP7_75t_L g3113 ( 
.A(n_2329),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2453),
.B(n_302),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2831),
.Y(n_3115)
);

BUFx6f_ASAP7_75t_L g3116 ( 
.A(n_2757),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2831),
.Y(n_3117)
);

INVx3_ASAP7_75t_L g3118 ( 
.A(n_2757),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2835),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2835),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_3071),
.B(n_2521),
.Y(n_3121)
);

AO21x1_ASAP7_75t_L g3122 ( 
.A1(n_2798),
.A2(n_2539),
.B(n_2615),
.Y(n_3122)
);

INVxp67_ASAP7_75t_SL g3123 ( 
.A(n_2988),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2800),
.Y(n_3124)
);

BUFx2_ASAP7_75t_L g3125 ( 
.A(n_3056),
.Y(n_3125)
);

INVx2_ASAP7_75t_SL g3126 ( 
.A(n_2730),
.Y(n_3126)
);

AND2x4_ASAP7_75t_L g3127 ( 
.A(n_2948),
.B(n_2461),
.Y(n_3127)
);

BUFx3_ASAP7_75t_L g3128 ( 
.A(n_2899),
.Y(n_3128)
);

AOI21xp5_ASAP7_75t_L g3129 ( 
.A1(n_2941),
.A2(n_2368),
.B(n_2671),
.Y(n_3129)
);

AOI221xp5_ASAP7_75t_L g3130 ( 
.A1(n_2820),
.A2(n_2435),
.B1(n_2444),
.B2(n_2688),
.C(n_2452),
.Y(n_3130)
);

BUFx6f_ASAP7_75t_L g3131 ( 
.A(n_2860),
.Y(n_3131)
);

AOI21xp5_ASAP7_75t_L g3132 ( 
.A1(n_3098),
.A2(n_2448),
.B(n_2516),
.Y(n_3132)
);

NAND2xp33_ASAP7_75t_L g3133 ( 
.A(n_2930),
.B(n_2529),
.Y(n_3133)
);

NOR2xp33_ASAP7_75t_L g3134 ( 
.A(n_2770),
.B(n_2290),
.Y(n_3134)
);

INVx5_ASAP7_75t_L g3135 ( 
.A(n_3056),
.Y(n_3135)
);

NOR2xp33_ASAP7_75t_L g3136 ( 
.A(n_3063),
.B(n_2621),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2725),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2818),
.Y(n_3138)
);

AOI221xp5_ASAP7_75t_L g3139 ( 
.A1(n_2729),
.A2(n_2618),
.B1(n_2593),
.B2(n_2517),
.C(n_2515),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2836),
.Y(n_3140)
);

BUFx3_ASAP7_75t_L g3141 ( 
.A(n_2762),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2884),
.B(n_2433),
.Y(n_3142)
);

BUFx12f_ASAP7_75t_L g3143 ( 
.A(n_2812),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2844),
.Y(n_3144)
);

NOR2xp67_ASAP7_75t_L g3145 ( 
.A(n_3002),
.B(n_2402),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2765),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_2742),
.B(n_2486),
.Y(n_3147)
);

AND2x2_ASAP7_75t_L g3148 ( 
.A(n_2832),
.B(n_2721),
.Y(n_3148)
);

CKINVDCx16_ASAP7_75t_R g3149 ( 
.A(n_2811),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_2777),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_2778),
.Y(n_3151)
);

AND2x2_ASAP7_75t_L g3152 ( 
.A(n_2759),
.B(n_2449),
.Y(n_3152)
);

AOI21xp5_ASAP7_75t_L g3153 ( 
.A1(n_3098),
.A2(n_2568),
.B(n_2560),
.Y(n_3153)
);

BUFx2_ASAP7_75t_L g3154 ( 
.A(n_3056),
.Y(n_3154)
);

AND2x2_ASAP7_75t_L g3155 ( 
.A(n_2772),
.B(n_2329),
.Y(n_3155)
);

INVx3_ASAP7_75t_L g3156 ( 
.A(n_2860),
.Y(n_3156)
);

AND2x6_ASAP7_75t_L g3157 ( 
.A(n_2740),
.B(n_2560),
.Y(n_3157)
);

AND2x4_ASAP7_75t_L g3158 ( 
.A(n_2948),
.B(n_2461),
.Y(n_3158)
);

AOI21xp5_ASAP7_75t_L g3159 ( 
.A1(n_2952),
.A2(n_2568),
.B(n_2560),
.Y(n_3159)
);

BUFx12f_ASAP7_75t_L g3160 ( 
.A(n_2750),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_2845),
.B(n_2856),
.Y(n_3161)
);

INVx5_ASAP7_75t_L g3162 ( 
.A(n_3056),
.Y(n_3162)
);

AOI21xp33_ASAP7_75t_L g3163 ( 
.A1(n_2876),
.A2(n_2612),
.B(n_2609),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2862),
.Y(n_3164)
);

OAI22xp33_ASAP7_75t_L g3165 ( 
.A1(n_2839),
.A2(n_2610),
.B1(n_2615),
.B2(n_2635),
.Y(n_3165)
);

INVx6_ASAP7_75t_L g3166 ( 
.A(n_2762),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2865),
.Y(n_3167)
);

OR2x2_ASAP7_75t_L g3168 ( 
.A(n_2768),
.B(n_2383),
.Y(n_3168)
);

OR2x6_ASAP7_75t_L g3169 ( 
.A(n_3001),
.B(n_2467),
.Y(n_3169)
);

OR2x6_ASAP7_75t_L g3170 ( 
.A(n_3026),
.B(n_2434),
.Y(n_3170)
);

OAI22xp33_ASAP7_75t_L g3171 ( 
.A1(n_3090),
.A2(n_2610),
.B1(n_2350),
.B2(n_2390),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_SL g3172 ( 
.A(n_2804),
.B(n_2529),
.Y(n_3172)
);

INVx1_ASAP7_75t_SL g3173 ( 
.A(n_3091),
.Y(n_3173)
);

HB1xp67_ASAP7_75t_L g3174 ( 
.A(n_3084),
.Y(n_3174)
);

BUFx2_ASAP7_75t_L g3175 ( 
.A(n_3090),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2871),
.Y(n_3176)
);

INVx3_ASAP7_75t_L g3177 ( 
.A(n_3002),
.Y(n_3177)
);

BUFx10_ASAP7_75t_L g3178 ( 
.A(n_2961),
.Y(n_3178)
);

INVx2_ASAP7_75t_SL g3179 ( 
.A(n_2852),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_2815),
.Y(n_3180)
);

INVx6_ASAP7_75t_L g3181 ( 
.A(n_2852),
.Y(n_3181)
);

INVx3_ASAP7_75t_L g3182 ( 
.A(n_2918),
.Y(n_3182)
);

CKINVDCx5p33_ASAP7_75t_R g3183 ( 
.A(n_2951),
.Y(n_3183)
);

INVx1_ASAP7_75t_SL g3184 ( 
.A(n_2758),
.Y(n_3184)
);

BUFx2_ASAP7_75t_L g3185 ( 
.A(n_3013),
.Y(n_3185)
);

INVx4_ASAP7_75t_L g3186 ( 
.A(n_2901),
.Y(n_3186)
);

INVx2_ASAP7_75t_L g3187 ( 
.A(n_2827),
.Y(n_3187)
);

INVx4_ASAP7_75t_L g3188 ( 
.A(n_2737),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2873),
.B(n_3111),
.Y(n_3189)
);

CKINVDCx20_ASAP7_75t_R g3190 ( 
.A(n_2738),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_3087),
.B(n_2269),
.Y(n_3191)
);

HB1xp67_ASAP7_75t_L g3192 ( 
.A(n_2779),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_3037),
.B(n_2606),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2879),
.Y(n_3194)
);

BUFx2_ASAP7_75t_L g3195 ( 
.A(n_3018),
.Y(n_3195)
);

BUFx2_ASAP7_75t_L g3196 ( 
.A(n_3019),
.Y(n_3196)
);

AOI22xp33_ASAP7_75t_L g3197 ( 
.A1(n_2736),
.A2(n_2546),
.B1(n_2489),
.B2(n_2472),
.Y(n_3197)
);

CKINVDCx16_ASAP7_75t_R g3198 ( 
.A(n_2803),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2894),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2895),
.Y(n_3200)
);

INVx3_ASAP7_75t_L g3201 ( 
.A(n_2918),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2910),
.Y(n_3202)
);

AOI21xp5_ASAP7_75t_L g3203 ( 
.A1(n_3105),
.A2(n_2628),
.B(n_2568),
.Y(n_3203)
);

OAI221xp5_ASAP7_75t_L g3204 ( 
.A1(n_2998),
.A2(n_2512),
.B1(n_2538),
.B2(n_2707),
.C(n_2496),
.Y(n_3204)
);

INVx4_ASAP7_75t_L g3205 ( 
.A(n_2769),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2916),
.Y(n_3206)
);

INVx2_ASAP7_75t_L g3207 ( 
.A(n_2837),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_2764),
.B(n_2587),
.Y(n_3208)
);

AOI22xp33_ASAP7_75t_L g3209 ( 
.A1(n_3033),
.A2(n_2616),
.B1(n_2596),
.B2(n_2502),
.Y(n_3209)
);

INVx3_ASAP7_75t_L g3210 ( 
.A(n_2990),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2922),
.Y(n_3211)
);

BUFx2_ASAP7_75t_L g3212 ( 
.A(n_2813),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_2854),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2940),
.Y(n_3214)
);

INVx4_ASAP7_75t_L g3215 ( 
.A(n_2783),
.Y(n_3215)
);

BUFx6f_ASAP7_75t_L g3216 ( 
.A(n_2799),
.Y(n_3216)
);

BUFx2_ASAP7_75t_L g3217 ( 
.A(n_2830),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2775),
.B(n_2650),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_2791),
.B(n_2631),
.Y(n_3219)
);

BUFx3_ASAP7_75t_L g3220 ( 
.A(n_3050),
.Y(n_3220)
);

NOR2xp33_ASAP7_75t_L g3221 ( 
.A(n_2751),
.B(n_2320),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_2925),
.Y(n_3222)
);

INVx2_ASAP7_75t_L g3223 ( 
.A(n_2958),
.Y(n_3223)
);

AND2x2_ASAP7_75t_L g3224 ( 
.A(n_2735),
.B(n_2632),
.Y(n_3224)
);

BUFx6f_ASAP7_75t_L g3225 ( 
.A(n_2904),
.Y(n_3225)
);

BUFx2_ASAP7_75t_L g3226 ( 
.A(n_2868),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_2926),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2929),
.Y(n_3228)
);

BUFx2_ASAP7_75t_L g3229 ( 
.A(n_2891),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2727),
.B(n_2636),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2932),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2782),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_2790),
.Y(n_3233)
);

INVx3_ASAP7_75t_L g3234 ( 
.A(n_2990),
.Y(n_3234)
);

BUFx6f_ASAP7_75t_L g3235 ( 
.A(n_2752),
.Y(n_3235)
);

BUFx2_ASAP7_75t_L g3236 ( 
.A(n_2950),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2936),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_2748),
.Y(n_3238)
);

CKINVDCx5p33_ASAP7_75t_R g3239 ( 
.A(n_2745),
.Y(n_3239)
);

INVx2_ASAP7_75t_SL g3240 ( 
.A(n_2980),
.Y(n_3240)
);

AND2x4_ASAP7_75t_L g3241 ( 
.A(n_3048),
.B(n_2475),
.Y(n_3241)
);

INVx4_ASAP7_75t_L g3242 ( 
.A(n_2841),
.Y(n_3242)
);

OAI22xp5_ASAP7_75t_L g3243 ( 
.A1(n_2994),
.A2(n_2627),
.B1(n_2640),
.B2(n_2379),
.Y(n_3243)
);

NOR2xp33_ASAP7_75t_L g3244 ( 
.A(n_3059),
.B(n_2328),
.Y(n_3244)
);

INVx1_ASAP7_75t_SL g3245 ( 
.A(n_3093),
.Y(n_3245)
);

BUFx6f_ASAP7_75t_SL g3246 ( 
.A(n_2979),
.Y(n_3246)
);

AND2x4_ASAP7_75t_L g3247 ( 
.A(n_3048),
.B(n_2475),
.Y(n_3247)
);

BUFx3_ASAP7_75t_L g3248 ( 
.A(n_2889),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_3069),
.Y(n_3249)
);

BUFx2_ASAP7_75t_L g3250 ( 
.A(n_2752),
.Y(n_3250)
);

INVx2_ASAP7_75t_L g3251 ( 
.A(n_3070),
.Y(n_3251)
);

INVx1_ASAP7_75t_SL g3252 ( 
.A(n_2763),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_3078),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_2753),
.Y(n_3254)
);

BUFx2_ASAP7_75t_L g3255 ( 
.A(n_2752),
.Y(n_3255)
);

AND2x4_ASAP7_75t_L g3256 ( 
.A(n_3048),
.B(n_2530),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2760),
.Y(n_3257)
);

BUFx3_ASAP7_75t_L g3258 ( 
.A(n_2915),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2771),
.Y(n_3259)
);

CKINVDCx14_ASAP7_75t_R g3260 ( 
.A(n_2870),
.Y(n_3260)
);

INVxp67_ASAP7_75t_L g3261 ( 
.A(n_2756),
.Y(n_3261)
);

CKINVDCx5p33_ASAP7_75t_R g3262 ( 
.A(n_3005),
.Y(n_3262)
);

AND2x2_ASAP7_75t_L g3263 ( 
.A(n_2767),
.B(n_2622),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_2776),
.Y(n_3264)
);

BUFx6f_ASAP7_75t_L g3265 ( 
.A(n_2766),
.Y(n_3265)
);

AOI21xp5_ASAP7_75t_L g3266 ( 
.A1(n_3105),
.A2(n_2661),
.B(n_2628),
.Y(n_3266)
);

INVx3_ASAP7_75t_L g3267 ( 
.A(n_2980),
.Y(n_3267)
);

CKINVDCx8_ASAP7_75t_R g3268 ( 
.A(n_2863),
.Y(n_3268)
);

OR2x2_ASAP7_75t_L g3269 ( 
.A(n_2991),
.B(n_2622),
.Y(n_3269)
);

AND2x4_ASAP7_75t_L g3270 ( 
.A(n_3073),
.B(n_2530),
.Y(n_3270)
);

AOI22xp5_ASAP7_75t_L g3271 ( 
.A1(n_2833),
.A2(n_2492),
.B1(n_2639),
.B2(n_2668),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_2792),
.Y(n_3272)
);

AND2x4_ASAP7_75t_L g3273 ( 
.A(n_3073),
.B(n_2672),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_2959),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_2795),
.Y(n_3275)
);

BUFx2_ASAP7_75t_L g3276 ( 
.A(n_2766),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_2909),
.B(n_2629),
.Y(n_3277)
);

BUFx6f_ASAP7_75t_L g3278 ( 
.A(n_2766),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_2727),
.B(n_2630),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_2963),
.Y(n_3280)
);

AND2x2_ASAP7_75t_L g3281 ( 
.A(n_2843),
.B(n_2633),
.Y(n_3281)
);

CKINVDCx5p33_ASAP7_75t_R g3282 ( 
.A(n_3049),
.Y(n_3282)
);

BUFx2_ASAP7_75t_L g3283 ( 
.A(n_2787),
.Y(n_3283)
);

BUFx2_ASAP7_75t_L g3284 ( 
.A(n_2787),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_2732),
.B(n_2595),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_2732),
.B(n_2595),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_2806),
.Y(n_3287)
);

AND2x4_ASAP7_75t_L g3288 ( 
.A(n_3073),
.B(n_2617),
.Y(n_3288)
);

HB1xp67_ASAP7_75t_L g3289 ( 
.A(n_2807),
.Y(n_3289)
);

INVx2_ASAP7_75t_SL g3290 ( 
.A(n_2921),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_3080),
.Y(n_3291)
);

NOR2xp33_ASAP7_75t_L g3292 ( 
.A(n_3061),
.B(n_2601),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3109),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_2734),
.B(n_2601),
.Y(n_3294)
);

INVx2_ASAP7_75t_L g3295 ( 
.A(n_2808),
.Y(n_3295)
);

INVx3_ASAP7_75t_L g3296 ( 
.A(n_3020),
.Y(n_3296)
);

AOI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_2992),
.A2(n_2661),
.B(n_2628),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3109),
.Y(n_3298)
);

CKINVDCx8_ASAP7_75t_R g3299 ( 
.A(n_2863),
.Y(n_3299)
);

AOI21xp5_ASAP7_75t_L g3300 ( 
.A1(n_3006),
.A2(n_2661),
.B(n_2674),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_2734),
.B(n_2660),
.Y(n_3301)
);

AOI22xp5_ASAP7_75t_L g3302 ( 
.A1(n_2896),
.A2(n_2651),
.B1(n_2421),
.B2(n_2357),
.Y(n_3302)
);

INVx2_ASAP7_75t_L g3303 ( 
.A(n_2858),
.Y(n_3303)
);

AOI22xp33_ASAP7_75t_SL g3304 ( 
.A1(n_2944),
.A2(n_2548),
.B1(n_2460),
.B2(n_2602),
.Y(n_3304)
);

OAI22xp33_ASAP7_75t_L g3305 ( 
.A1(n_3029),
.A2(n_2984),
.B1(n_3064),
.B2(n_2878),
.Y(n_3305)
);

OR2x6_ASAP7_75t_L g3306 ( 
.A(n_3029),
.B(n_2528),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_2867),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_2821),
.B(n_2647),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_2821),
.B(n_2528),
.Y(n_3309)
);

NOR2xp33_ASAP7_75t_L g3310 ( 
.A(n_3062),
.B(n_2652),
.Y(n_3310)
);

OAI221xp5_ASAP7_75t_L g3311 ( 
.A1(n_2954),
.A2(n_2648),
.B1(n_2264),
.B2(n_2254),
.C(n_2358),
.Y(n_3311)
);

INVx2_ASAP7_75t_SL g3312 ( 
.A(n_2938),
.Y(n_3312)
);

INVx5_ASAP7_75t_L g3313 ( 
.A(n_2787),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_2869),
.Y(n_3314)
);

AND2x4_ASAP7_75t_L g3315 ( 
.A(n_2749),
.B(n_2280),
.Y(n_3315)
);

AOI21xp5_ASAP7_75t_L g3316 ( 
.A1(n_3007),
.A2(n_2670),
.B(n_2343),
.Y(n_3316)
);

INVx2_ASAP7_75t_L g3317 ( 
.A(n_2875),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_2902),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_2822),
.B(n_2584),
.Y(n_3319)
);

NAND2x1p5_ASAP7_75t_L g3320 ( 
.A(n_2817),
.B(n_2576),
.Y(n_3320)
);

A2O1A1Ixp33_ASAP7_75t_L g3321 ( 
.A1(n_2797),
.A2(n_2648),
.B(n_2343),
.C(n_2567),
.Y(n_3321)
);

BUFx3_ASAP7_75t_L g3322 ( 
.A(n_2975),
.Y(n_3322)
);

AOI22xp5_ASAP7_75t_L g3323 ( 
.A1(n_2802),
.A2(n_2584),
.B1(n_2669),
.B2(n_2358),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_2822),
.Y(n_3324)
);

INVx5_ASAP7_75t_L g3325 ( 
.A(n_2874),
.Y(n_3325)
);

INVx2_ASAP7_75t_SL g3326 ( 
.A(n_3020),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_2911),
.Y(n_3327)
);

AOI22xp5_ASAP7_75t_L g3328 ( 
.A1(n_2819),
.A2(n_2739),
.B1(n_2970),
.B2(n_2733),
.Y(n_3328)
);

AOI21x1_ASAP7_75t_L g3329 ( 
.A1(n_2731),
.A2(n_2653),
.B(n_2376),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_3034),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_2829),
.B(n_2584),
.Y(n_3331)
);

BUFx3_ASAP7_75t_L g3332 ( 
.A(n_3017),
.Y(n_3332)
);

A2O1A1Ixp33_ASAP7_75t_L g3333 ( 
.A1(n_2969),
.A2(n_2316),
.B(n_2298),
.C(n_2723),
.Y(n_3333)
);

INVx2_ASAP7_75t_SL g3334 ( 
.A(n_2877),
.Y(n_3334)
);

INVx3_ASAP7_75t_L g3335 ( 
.A(n_3065),
.Y(n_3335)
);

HB1xp67_ASAP7_75t_L g3336 ( 
.A(n_2969),
.Y(n_3336)
);

AND2x4_ASAP7_75t_L g3337 ( 
.A(n_2749),
.B(n_2280),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_2829),
.Y(n_3338)
);

INVx3_ASAP7_75t_L g3339 ( 
.A(n_3042),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3099),
.Y(n_3340)
);

AND2x2_ASAP7_75t_L g3341 ( 
.A(n_2796),
.B(n_303),
.Y(n_3341)
);

BUFx2_ASAP7_75t_L g3342 ( 
.A(n_2874),
.Y(n_3342)
);

BUFx3_ASAP7_75t_L g3343 ( 
.A(n_3027),
.Y(n_3343)
);

BUFx2_ASAP7_75t_L g3344 ( 
.A(n_2874),
.Y(n_3344)
);

AND2x2_ASAP7_75t_L g3345 ( 
.A(n_3067),
.B(n_304),
.Y(n_3345)
);

BUFx12f_ASAP7_75t_L g3346 ( 
.A(n_2995),
.Y(n_3346)
);

BUFx2_ASAP7_75t_L g3347 ( 
.A(n_2898),
.Y(n_3347)
);

OAI221xp5_ASAP7_75t_L g3348 ( 
.A1(n_3100),
.A2(n_2379),
.B1(n_2666),
.B2(n_2665),
.C(n_2655),
.Y(n_3348)
);

INVx1_ASAP7_75t_SL g3349 ( 
.A(n_3101),
.Y(n_3349)
);

BUFx8_ASAP7_75t_L g3350 ( 
.A(n_2788),
.Y(n_3350)
);

AND2x4_ASAP7_75t_L g3351 ( 
.A(n_2784),
.B(n_2296),
.Y(n_3351)
);

AOI22xp5_ASAP7_75t_L g3352 ( 
.A1(n_3054),
.A2(n_2584),
.B1(n_2298),
.B2(n_2316),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_2913),
.Y(n_3353)
);

AOI22xp33_ASAP7_75t_L g3354 ( 
.A1(n_2823),
.A2(n_2642),
.B1(n_2662),
.B2(n_2676),
.Y(n_3354)
);

AND2x4_ASAP7_75t_L g3355 ( 
.A(n_2784),
.B(n_3042),
.Y(n_3355)
);

AOI22xp33_ASAP7_75t_L g3356 ( 
.A1(n_3004),
.A2(n_2389),
.B1(n_2624),
.B2(n_2623),
.Y(n_3356)
);

A2O1A1Ixp33_ASAP7_75t_SL g3357 ( 
.A1(n_2931),
.A2(n_2654),
.B(n_2626),
.C(n_2664),
.Y(n_3357)
);

BUFx3_ASAP7_75t_L g3358 ( 
.A(n_2881),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_SL g3359 ( 
.A(n_2985),
.B(n_2576),
.Y(n_3359)
);

INVx3_ASAP7_75t_L g3360 ( 
.A(n_3045),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3099),
.Y(n_3361)
);

INVx2_ASAP7_75t_L g3362 ( 
.A(n_2919),
.Y(n_3362)
);

BUFx2_ASAP7_75t_L g3363 ( 
.A(n_2898),
.Y(n_3363)
);

AOI22xp5_ASAP7_75t_L g3364 ( 
.A1(n_2905),
.A2(n_2389),
.B1(n_2457),
.B2(n_2573),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_2978),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_SL g3366 ( 
.A(n_2985),
.B(n_2576),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_2981),
.Y(n_3367)
);

BUFx2_ASAP7_75t_L g3368 ( 
.A(n_2898),
.Y(n_3368)
);

BUFx6f_ASAP7_75t_L g3369 ( 
.A(n_2903),
.Y(n_3369)
);

NAND3x1_ASAP7_75t_L g3370 ( 
.A(n_3000),
.B(n_2641),
.C(n_2626),
.Y(n_3370)
);

BUFx6f_ASAP7_75t_L g3371 ( 
.A(n_2903),
.Y(n_3371)
);

AOI21xp5_ASAP7_75t_L g3372 ( 
.A1(n_3008),
.A2(n_2675),
.B(n_2296),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3096),
.B(n_2389),
.Y(n_3373)
);

AND2x4_ASAP7_75t_L g3374 ( 
.A(n_3045),
.B(n_2726),
.Y(n_3374)
);

AND2x2_ASAP7_75t_L g3375 ( 
.A(n_2814),
.B(n_304),
.Y(n_3375)
);

BUFx2_ASAP7_75t_SL g3376 ( 
.A(n_2754),
.Y(n_3376)
);

INVx5_ASAP7_75t_L g3377 ( 
.A(n_2903),
.Y(n_3377)
);

OAI22xp5_ASAP7_75t_L g3378 ( 
.A1(n_3083),
.A2(n_2457),
.B1(n_2659),
.B2(n_2657),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_2949),
.B(n_2389),
.Y(n_3379)
);

OAI22xp5_ASAP7_75t_L g3380 ( 
.A1(n_3060),
.A2(n_2659),
.B1(n_2657),
.B2(n_2376),
.Y(n_3380)
);

NAND2x1p5_ASAP7_75t_L g3381 ( 
.A(n_2726),
.B(n_2657),
.Y(n_3381)
);

NAND2x1p5_ASAP7_75t_L g3382 ( 
.A(n_2741),
.B(n_2659),
.Y(n_3382)
);

INVx2_ASAP7_75t_L g3383 ( 
.A(n_2996),
.Y(n_3383)
);

AND2x2_ASAP7_75t_L g3384 ( 
.A(n_3021),
.B(n_305),
.Y(n_3384)
);

INVx1_ASAP7_75t_SL g3385 ( 
.A(n_2887),
.Y(n_3385)
);

BUFx4f_ASAP7_75t_L g3386 ( 
.A(n_2761),
.Y(n_3386)
);

BUFx2_ASAP7_75t_SL g3387 ( 
.A(n_2885),
.Y(n_3387)
);

AND2x4_ASAP7_75t_L g3388 ( 
.A(n_2741),
.B(n_2296),
.Y(n_3388)
);

AOI22xp33_ASAP7_75t_L g3389 ( 
.A1(n_3015),
.A2(n_2360),
.B1(n_2364),
.B2(n_2347),
.Y(n_3389)
);

INVx3_ASAP7_75t_L g3390 ( 
.A(n_2897),
.Y(n_3390)
);

AND2x4_ASAP7_75t_L g3391 ( 
.A(n_2744),
.B(n_2680),
.Y(n_3391)
);

AND2x4_ASAP7_75t_L g3392 ( 
.A(n_2934),
.B(n_2680),
.Y(n_3392)
);

BUFx12f_ASAP7_75t_L g3393 ( 
.A(n_3053),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3038),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_2957),
.B(n_306),
.Y(n_3395)
);

OAI21xp33_ASAP7_75t_L g3396 ( 
.A1(n_2946),
.A2(n_2380),
.B(n_2395),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_2912),
.B(n_306),
.Y(n_3397)
);

AOI22xp33_ASAP7_75t_SL g3398 ( 
.A1(n_3077),
.A2(n_2347),
.B1(n_2689),
.B2(n_2680),
.Y(n_3398)
);

INVx3_ASAP7_75t_L g3399 ( 
.A(n_2744),
.Y(n_3399)
);

INVx2_ASAP7_75t_L g3400 ( 
.A(n_3051),
.Y(n_3400)
);

AOI22xp33_ASAP7_75t_L g3401 ( 
.A1(n_3025),
.A2(n_2347),
.B1(n_2573),
.B2(n_2689),
.Y(n_3401)
);

OAI22xp33_ASAP7_75t_L g3402 ( 
.A1(n_2933),
.A2(n_2689),
.B1(n_2347),
.B2(n_309),
.Y(n_3402)
);

AO22x1_ASAP7_75t_L g3403 ( 
.A1(n_2740),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3066),
.Y(n_3404)
);

HB1xp67_ASAP7_75t_L g3405 ( 
.A(n_3003),
.Y(n_3405)
);

AOI21xp5_ASAP7_75t_L g3406 ( 
.A1(n_3031),
.A2(n_3041),
.B(n_2923),
.Y(n_3406)
);

BUFx6f_ASAP7_75t_L g3407 ( 
.A(n_2907),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_3110),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_2774),
.Y(n_3409)
);

OR2x6_ASAP7_75t_L g3410 ( 
.A(n_2809),
.B(n_307),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_2781),
.Y(n_3411)
);

NOR2xp33_ASAP7_75t_L g3412 ( 
.A(n_3032),
.B(n_308),
.Y(n_3412)
);

NAND2xp33_ASAP7_75t_L g3413 ( 
.A(n_2930),
.B(n_310),
.Y(n_3413)
);

INVx2_ASAP7_75t_SL g3414 ( 
.A(n_3021),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_2786),
.Y(n_3415)
);

AND2x4_ASAP7_75t_L g3416 ( 
.A(n_2851),
.B(n_2794),
.Y(n_3416)
);

OAI22xp5_ASAP7_75t_L g3417 ( 
.A1(n_2937),
.A2(n_313),
.B1(n_310),
.B2(n_311),
.Y(n_3417)
);

BUFx12f_ASAP7_75t_L g3418 ( 
.A(n_2785),
.Y(n_3418)
);

INVx4_ASAP7_75t_L g3419 ( 
.A(n_2851),
.Y(n_3419)
);

OAI22xp5_ASAP7_75t_L g3420 ( 
.A1(n_3304),
.A2(n_2971),
.B1(n_2883),
.B2(n_2960),
.Y(n_3420)
);

INVx2_ASAP7_75t_L g3421 ( 
.A(n_3249),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_L g3422 ( 
.A(n_3189),
.B(n_3035),
.Y(n_3422)
);

OA21x2_ASAP7_75t_L g3423 ( 
.A1(n_3132),
.A2(n_3102),
.B(n_2892),
.Y(n_3423)
);

HB1xp67_ASAP7_75t_L g3424 ( 
.A(n_3174),
.Y(n_3424)
);

OAI21x1_ASAP7_75t_L g3425 ( 
.A1(n_3329),
.A2(n_2747),
.B(n_3047),
.Y(n_3425)
);

OAI21x1_ASAP7_75t_L g3426 ( 
.A1(n_3372),
.A2(n_3058),
.B(n_3047),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3324),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3338),
.Y(n_3428)
);

OAI21x1_ASAP7_75t_L g3429 ( 
.A1(n_3159),
.A2(n_3068),
.B(n_3058),
.Y(n_3429)
);

NOR2xp33_ASAP7_75t_L g3430 ( 
.A(n_3268),
.B(n_2793),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_3124),
.B(n_3040),
.Y(n_3431)
);

OAI21x1_ASAP7_75t_L g3432 ( 
.A1(n_3153),
.A2(n_3074),
.B(n_3068),
.Y(n_3432)
);

BUFx6f_ASAP7_75t_L g3433 ( 
.A(n_3131),
.Y(n_3433)
);

AO21x2_ASAP7_75t_L g3434 ( 
.A1(n_3163),
.A2(n_3052),
.B(n_3044),
.Y(n_3434)
);

OAI222xp33_ASAP7_75t_L g3435 ( 
.A1(n_3299),
.A2(n_2943),
.B1(n_3081),
.B2(n_2973),
.C1(n_2986),
.C2(n_2977),
.Y(n_3435)
);

OAI21x1_ASAP7_75t_L g3436 ( 
.A1(n_3203),
.A2(n_3074),
.B(n_2840),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_3115),
.Y(n_3437)
);

OAI21x1_ASAP7_75t_L g3438 ( 
.A1(n_3266),
.A2(n_2840),
.B(n_2794),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3117),
.Y(n_3439)
);

INVx4_ASAP7_75t_L g3440 ( 
.A(n_3135),
.Y(n_3440)
);

BUFx3_ASAP7_75t_L g3441 ( 
.A(n_3186),
.Y(n_3441)
);

OA21x2_ASAP7_75t_L g3442 ( 
.A1(n_3129),
.A2(n_3108),
.B(n_2983),
.Y(n_3442)
);

NAND3xp33_ASAP7_75t_L g3443 ( 
.A(n_3134),
.B(n_2947),
.C(n_2780),
.Y(n_3443)
);

AOI22xp33_ASAP7_75t_L g3444 ( 
.A1(n_3171),
.A2(n_2789),
.B1(n_2864),
.B2(n_2846),
.Y(n_3444)
);

OAI21x1_ASAP7_75t_L g3445 ( 
.A1(n_3370),
.A2(n_2914),
.B(n_2890),
.Y(n_3445)
);

OAI21xp5_ASAP7_75t_L g3446 ( 
.A1(n_3139),
.A2(n_2920),
.B(n_2962),
.Y(n_3446)
);

AOI22xp33_ASAP7_75t_L g3447 ( 
.A1(n_3122),
.A2(n_3003),
.B1(n_2805),
.B2(n_2828),
.Y(n_3447)
);

INVx1_ASAP7_75t_SL g3448 ( 
.A(n_3376),
.Y(n_3448)
);

AOI211xp5_ASAP7_75t_L g3449 ( 
.A1(n_3305),
.A2(n_2927),
.B(n_2810),
.C(n_3028),
.Y(n_3449)
);

OR2x2_ASAP7_75t_L g3450 ( 
.A(n_3192),
.B(n_2886),
.Y(n_3450)
);

A2O1A1Ixp33_ASAP7_75t_L g3451 ( 
.A1(n_3413),
.A2(n_2805),
.B(n_2828),
.C(n_2785),
.Y(n_3451)
);

AOI21xp5_ASAP7_75t_L g3452 ( 
.A1(n_3321),
.A2(n_2935),
.B(n_2907),
.Y(n_3452)
);

OAI21x1_ASAP7_75t_L g3453 ( 
.A1(n_3297),
.A2(n_2914),
.B(n_2890),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3138),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_3251),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3140),
.Y(n_3456)
);

HB1xp67_ASAP7_75t_L g3457 ( 
.A(n_3289),
.Y(n_3457)
);

AND2x4_ASAP7_75t_L g3458 ( 
.A(n_3135),
.B(n_2850),
.Y(n_3458)
);

AOI221xp5_ASAP7_75t_L g3459 ( 
.A1(n_3165),
.A2(n_2724),
.B1(n_2855),
.B2(n_2997),
.C(n_3057),
.Y(n_3459)
);

HB1xp67_ASAP7_75t_L g3460 ( 
.A(n_3336),
.Y(n_3460)
);

O2A1O1Ixp33_ASAP7_75t_L g3461 ( 
.A1(n_3121),
.A2(n_3142),
.B(n_3357),
.C(n_2882),
.Y(n_3461)
);

AOI22xp33_ASAP7_75t_L g3462 ( 
.A1(n_3130),
.A2(n_2850),
.B1(n_3086),
.B2(n_3085),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3144),
.Y(n_3463)
);

OAI21x1_ASAP7_75t_L g3464 ( 
.A1(n_3300),
.A2(n_3316),
.B(n_3406),
.Y(n_3464)
);

OAI21x1_ASAP7_75t_L g3465 ( 
.A1(n_3379),
.A2(n_3401),
.B(n_3380),
.Y(n_3465)
);

NOR2xp33_ASAP7_75t_L g3466 ( 
.A(n_3175),
.B(n_2826),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_3164),
.B(n_2967),
.Y(n_3467)
);

INVx3_ASAP7_75t_L g3468 ( 
.A(n_3135),
.Y(n_3468)
);

NAND2xp33_ASAP7_75t_L g3469 ( 
.A(n_3157),
.B(n_2930),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3119),
.Y(n_3470)
);

OAI21x1_ASAP7_75t_L g3471 ( 
.A1(n_3319),
.A2(n_3010),
.B(n_2955),
.Y(n_3471)
);

AOI21xp5_ASAP7_75t_L g3472 ( 
.A1(n_3333),
.A2(n_2935),
.B(n_2907),
.Y(n_3472)
);

OA21x2_ASAP7_75t_L g3473 ( 
.A1(n_3354),
.A2(n_3114),
.B(n_3112),
.Y(n_3473)
);

NOR2xp33_ASAP7_75t_L g3474 ( 
.A(n_3175),
.B(n_3039),
.Y(n_3474)
);

OAI21x1_ASAP7_75t_L g3475 ( 
.A1(n_3331),
.A2(n_3010),
.B(n_2955),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3120),
.Y(n_3476)
);

OAI21x1_ASAP7_75t_L g3477 ( 
.A1(n_3378),
.A2(n_3011),
.B(n_3082),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3167),
.B(n_2974),
.Y(n_3478)
);

OAI221xp5_ASAP7_75t_L g3479 ( 
.A1(n_3328),
.A2(n_2728),
.B1(n_2972),
.B2(n_2880),
.C(n_2872),
.Y(n_3479)
);

AND2x2_ASAP7_75t_L g3480 ( 
.A(n_3193),
.B(n_3046),
.Y(n_3480)
);

OAI21x1_ASAP7_75t_L g3481 ( 
.A1(n_3373),
.A2(n_3011),
.B(n_3104),
.Y(n_3481)
);

NOR2x1_ASAP7_75t_SL g3482 ( 
.A(n_3162),
.B(n_3359),
.Y(n_3482)
);

OAI21x1_ASAP7_75t_L g3483 ( 
.A1(n_3366),
.A2(n_3107),
.B(n_2987),
.Y(n_3483)
);

BUFx2_ASAP7_75t_SL g3484 ( 
.A(n_3246),
.Y(n_3484)
);

INVx2_ASAP7_75t_L g3485 ( 
.A(n_3253),
.Y(n_3485)
);

INVx2_ASAP7_75t_SL g3486 ( 
.A(n_3166),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3293),
.Y(n_3487)
);

AO21x2_ASAP7_75t_L g3488 ( 
.A1(n_3402),
.A2(n_2906),
.B(n_2917),
.Y(n_3488)
);

OAI21x1_ASAP7_75t_L g3489 ( 
.A1(n_3320),
.A2(n_2976),
.B(n_2743),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3298),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3340),
.Y(n_3491)
);

BUFx2_ASAP7_75t_L g3492 ( 
.A(n_3418),
.Y(n_3492)
);

INVxp67_ASAP7_75t_SL g3493 ( 
.A(n_3123),
.Y(n_3493)
);

OAI222xp33_ASAP7_75t_L g3494 ( 
.A1(n_3410),
.A2(n_2755),
.B1(n_3046),
.B2(n_3113),
.C1(n_2965),
.C2(n_3106),
.Y(n_3494)
);

OAI21x1_ASAP7_75t_SL g3495 ( 
.A1(n_3414),
.A2(n_3079),
.B(n_3103),
.Y(n_3495)
);

OAI21x1_ASAP7_75t_L g3496 ( 
.A1(n_3361),
.A2(n_3030),
.B(n_3014),
.Y(n_3496)
);

AOI21xp5_ASAP7_75t_L g3497 ( 
.A1(n_3133),
.A2(n_2945),
.B(n_2935),
.Y(n_3497)
);

OAI21x1_ASAP7_75t_L g3498 ( 
.A1(n_3381),
.A2(n_2893),
.B(n_2888),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3176),
.B(n_2746),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3194),
.B(n_2801),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3199),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3200),
.Y(n_3502)
);

AND2x4_ASAP7_75t_L g3503 ( 
.A(n_3162),
.B(n_3079),
.Y(n_3503)
);

INVx2_ASAP7_75t_SL g3504 ( 
.A(n_3166),
.Y(n_3504)
);

BUFx2_ASAP7_75t_L g3505 ( 
.A(n_3260),
.Y(n_3505)
);

INVx1_ASAP7_75t_SL g3506 ( 
.A(n_3387),
.Y(n_3506)
);

OAI21x1_ASAP7_75t_L g3507 ( 
.A1(n_3382),
.A2(n_2928),
.B(n_2924),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3202),
.Y(n_3508)
);

OAI21x1_ASAP7_75t_L g3509 ( 
.A1(n_3364),
.A2(n_3294),
.B(n_3389),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3206),
.Y(n_3510)
);

AOI22xp33_ASAP7_75t_L g3511 ( 
.A1(n_3148),
.A2(n_2900),
.B1(n_3043),
.B2(n_2956),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3211),
.Y(n_3512)
);

OAI22xp33_ASAP7_75t_L g3513 ( 
.A1(n_3410),
.A2(n_3198),
.B1(n_3386),
.B2(n_3306),
.Y(n_3513)
);

NOR2xp33_ASAP7_75t_L g3514 ( 
.A(n_3205),
.B(n_3022),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3137),
.Y(n_3515)
);

OA21x2_ASAP7_75t_L g3516 ( 
.A1(n_3125),
.A2(n_3072),
.B(n_3055),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3214),
.Y(n_3517)
);

AND2x4_ASAP7_75t_L g3518 ( 
.A(n_3162),
.B(n_2945),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3291),
.B(n_2816),
.Y(n_3519)
);

OAI21x1_ASAP7_75t_L g3520 ( 
.A1(n_3285),
.A2(n_2942),
.B(n_2939),
.Y(n_3520)
);

OAI21xp5_ASAP7_75t_L g3521 ( 
.A1(n_3197),
.A2(n_3097),
.B(n_2966),
.Y(n_3521)
);

AND2x2_ASAP7_75t_L g3522 ( 
.A(n_3277),
.B(n_3281),
.Y(n_3522)
);

AO21x2_ASAP7_75t_L g3523 ( 
.A1(n_3208),
.A2(n_2866),
.B(n_3075),
.Y(n_3523)
);

HB1xp67_ASAP7_75t_L g3524 ( 
.A(n_3405),
.Y(n_3524)
);

AO21x2_ASAP7_75t_L g3525 ( 
.A1(n_3271),
.A2(n_3092),
.B(n_3088),
.Y(n_3525)
);

OAI21x1_ASAP7_75t_L g3526 ( 
.A1(n_3286),
.A2(n_2825),
.B(n_2824),
.Y(n_3526)
);

OAI21x1_ASAP7_75t_L g3527 ( 
.A1(n_3399),
.A2(n_2838),
.B(n_2834),
.Y(n_3527)
);

BUFx6f_ASAP7_75t_L g3528 ( 
.A(n_3131),
.Y(n_3528)
);

O2A1O1Ixp5_ASAP7_75t_L g3529 ( 
.A1(n_3172),
.A2(n_3094),
.B(n_3095),
.C(n_2773),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3146),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3161),
.Y(n_3531)
);

AOI21xp5_ASAP7_75t_L g3532 ( 
.A1(n_3311),
.A2(n_2964),
.B(n_2945),
.Y(n_3532)
);

OAI21x1_ASAP7_75t_L g3533 ( 
.A1(n_3356),
.A2(n_2849),
.B(n_2848),
.Y(n_3533)
);

BUFx2_ASAP7_75t_L g3534 ( 
.A(n_3157),
.Y(n_3534)
);

AO21x2_ASAP7_75t_L g3535 ( 
.A1(n_3396),
.A2(n_2857),
.B(n_2853),
.Y(n_3535)
);

OAI21xp5_ASAP7_75t_L g3536 ( 
.A1(n_3204),
.A2(n_2968),
.B(n_2953),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_3224),
.B(n_3384),
.Y(n_3537)
);

NAND2x1p5_ASAP7_75t_L g3538 ( 
.A(n_3141),
.B(n_2964),
.Y(n_3538)
);

O2A1O1Ixp33_ASAP7_75t_SL g3539 ( 
.A1(n_3179),
.A2(n_2999),
.B(n_3023),
.C(n_3036),
.Y(n_3539)
);

NAND2x1p5_ASAP7_75t_L g3540 ( 
.A(n_3332),
.B(n_3188),
.Y(n_3540)
);

NAND2x1p5_ASAP7_75t_L g3541 ( 
.A(n_3215),
.B(n_2964),
.Y(n_3541)
);

AND2x4_ASAP7_75t_L g3542 ( 
.A(n_3125),
.B(n_3009),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3218),
.B(n_2859),
.Y(n_3543)
);

OR2x2_ASAP7_75t_L g3544 ( 
.A(n_3254),
.B(n_2993),
.Y(n_3544)
);

BUFx2_ASAP7_75t_L g3545 ( 
.A(n_3157),
.Y(n_3545)
);

INVx2_ASAP7_75t_L g3546 ( 
.A(n_3150),
.Y(n_3546)
);

OR2x2_ASAP7_75t_L g3547 ( 
.A(n_3264),
.B(n_2861),
.Y(n_3547)
);

INVxp67_ASAP7_75t_SL g3548 ( 
.A(n_3154),
.Y(n_3548)
);

AOI21x1_ASAP7_75t_L g3549 ( 
.A1(n_3154),
.A2(n_2982),
.B(n_3016),
.Y(n_3549)
);

BUFx3_ASAP7_75t_L g3550 ( 
.A(n_3128),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3238),
.Y(n_3551)
);

OAI21x1_ASAP7_75t_L g3552 ( 
.A1(n_3232),
.A2(n_2847),
.B(n_2842),
.Y(n_3552)
);

OAI21x1_ASAP7_75t_L g3553 ( 
.A1(n_3233),
.A2(n_2908),
.B(n_3024),
.Y(n_3553)
);

INVxp67_ASAP7_75t_SL g3554 ( 
.A(n_3185),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3257),
.Y(n_3555)
);

CKINVDCx5p33_ASAP7_75t_R g3556 ( 
.A(n_3190),
.Y(n_3556)
);

AOI21x1_ASAP7_75t_L g3557 ( 
.A1(n_3250),
.A2(n_2989),
.B(n_3012),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3222),
.B(n_3089),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3227),
.B(n_3228),
.Y(n_3559)
);

AND2x4_ASAP7_75t_L g3560 ( 
.A(n_3374),
.B(n_3009),
.Y(n_3560)
);

OAI21xp5_ASAP7_75t_L g3561 ( 
.A1(n_3417),
.A2(n_2930),
.B(n_3009),
.Y(n_3561)
);

NOR2xp33_ASAP7_75t_L g3562 ( 
.A(n_3242),
.B(n_313),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3231),
.B(n_3076),
.Y(n_3563)
);

AO21x2_ASAP7_75t_L g3564 ( 
.A1(n_3395),
.A2(n_2930),
.B(n_3076),
.Y(n_3564)
);

AOI222xp33_ASAP7_75t_L g3565 ( 
.A1(n_3136),
.A2(n_316),
.B1(n_318),
.B2(n_314),
.C1(n_315),
.C2(n_317),
.Y(n_3565)
);

NAND2x1p5_ASAP7_75t_L g3566 ( 
.A(n_3267),
.B(n_3076),
.Y(n_3566)
);

AND2x2_ASAP7_75t_L g3567 ( 
.A(n_3375),
.B(n_314),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3259),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3237),
.B(n_317),
.Y(n_3569)
);

INVx2_ASAP7_75t_SL g3570 ( 
.A(n_3181),
.Y(n_3570)
);

INVx2_ASAP7_75t_L g3571 ( 
.A(n_3151),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3274),
.B(n_319),
.Y(n_3572)
);

NOR2xp33_ASAP7_75t_L g3573 ( 
.A(n_3245),
.B(n_319),
.Y(n_3573)
);

AO21x2_ASAP7_75t_L g3574 ( 
.A1(n_3323),
.A2(n_320),
.B(n_321),
.Y(n_3574)
);

NOR2xp33_ASAP7_75t_SL g3575 ( 
.A(n_3181),
.B(n_320),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3180),
.Y(n_3576)
);

AOI21xp5_ASAP7_75t_L g3577 ( 
.A1(n_3348),
.A2(n_655),
.B(n_650),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3280),
.B(n_321),
.Y(n_3578)
);

OAI21x1_ASAP7_75t_L g3579 ( 
.A1(n_3187),
.A2(n_660),
.B(n_658),
.Y(n_3579)
);

AO31x2_ASAP7_75t_L g3580 ( 
.A1(n_3243),
.A2(n_662),
.A3(n_664),
.B(n_661),
.Y(n_3580)
);

AOI22xp33_ASAP7_75t_L g3581 ( 
.A1(n_3152),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_3581)
);

O2A1O1Ixp33_ASAP7_75t_L g3582 ( 
.A1(n_3409),
.A2(n_3411),
.B(n_3415),
.C(n_3397),
.Y(n_3582)
);

OAI21x1_ASAP7_75t_L g3583 ( 
.A1(n_3207),
.A2(n_3223),
.B(n_3213),
.Y(n_3583)
);

OAI21x1_ASAP7_75t_L g3584 ( 
.A1(n_3330),
.A2(n_666),
.B(n_665),
.Y(n_3584)
);

AND2x4_ASAP7_75t_L g3585 ( 
.A(n_3374),
.B(n_3355),
.Y(n_3585)
);

OAI21x1_ASAP7_75t_SL g3586 ( 
.A1(n_3419),
.A2(n_325),
.B(n_326),
.Y(n_3586)
);

AOI21xp5_ASAP7_75t_L g3587 ( 
.A1(n_3308),
.A2(n_668),
.B(n_667),
.Y(n_3587)
);

AO21x2_ASAP7_75t_L g3588 ( 
.A1(n_3352),
.A2(n_326),
.B(n_327),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_3272),
.Y(n_3589)
);

NOR2x1_ASAP7_75t_L g3590 ( 
.A(n_3182),
.B(n_327),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3365),
.Y(n_3591)
);

AND2x2_ASAP7_75t_L g3592 ( 
.A(n_3341),
.B(n_328),
.Y(n_3592)
);

AND2x4_ASAP7_75t_L g3593 ( 
.A(n_3355),
.B(n_329),
.Y(n_3593)
);

AOI22x1_ASAP7_75t_L g3594 ( 
.A1(n_3201),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.Y(n_3594)
);

AOI22xp33_ASAP7_75t_L g3595 ( 
.A1(n_3398),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.Y(n_3595)
);

OAI21x1_ASAP7_75t_L g3596 ( 
.A1(n_3275),
.A2(n_670),
.B(n_669),
.Y(n_3596)
);

BUFx2_ASAP7_75t_L g3597 ( 
.A(n_3358),
.Y(n_3597)
);

OAI21x1_ASAP7_75t_L g3598 ( 
.A1(n_3287),
.A2(n_673),
.B(n_672),
.Y(n_3598)
);

NOR2x1_ASAP7_75t_L g3599 ( 
.A(n_3306),
.B(n_3248),
.Y(n_3599)
);

AO21x2_ASAP7_75t_L g3600 ( 
.A1(n_3302),
.A2(n_333),
.B(n_334),
.Y(n_3600)
);

INVx2_ASAP7_75t_L g3601 ( 
.A(n_3295),
.Y(n_3601)
);

AND2x2_ASAP7_75t_L g3602 ( 
.A(n_3263),
.B(n_333),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3367),
.Y(n_3603)
);

AND2x2_ASAP7_75t_L g3604 ( 
.A(n_3155),
.B(n_335),
.Y(n_3604)
);

OA21x2_ASAP7_75t_L g3605 ( 
.A1(n_3230),
.A2(n_685),
.B(n_682),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_3303),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3394),
.Y(n_3607)
);

BUFx3_ASAP7_75t_L g3608 ( 
.A(n_3220),
.Y(n_3608)
);

CKINVDCx11_ASAP7_75t_R g3609 ( 
.A(n_3143),
.Y(n_3609)
);

OAI21x1_ASAP7_75t_L g3610 ( 
.A1(n_3307),
.A2(n_687),
.B(n_686),
.Y(n_3610)
);

AND2x2_ASAP7_75t_L g3611 ( 
.A(n_3345),
.B(n_336),
.Y(n_3611)
);

OAI21x1_ASAP7_75t_L g3612 ( 
.A1(n_3314),
.A2(n_691),
.B(n_689),
.Y(n_3612)
);

BUFx8_ASAP7_75t_L g3613 ( 
.A(n_3160),
.Y(n_3613)
);

OAI21x1_ASAP7_75t_L g3614 ( 
.A1(n_3317),
.A2(n_3327),
.B(n_3318),
.Y(n_3614)
);

AOI22xp33_ASAP7_75t_L g3615 ( 
.A1(n_3185),
.A2(n_340),
.B1(n_337),
.B2(n_338),
.Y(n_3615)
);

OA21x2_ASAP7_75t_L g3616 ( 
.A1(n_3250),
.A2(n_693),
.B(n_692),
.Y(n_3616)
);

AOI21xp5_ASAP7_75t_L g3617 ( 
.A1(n_3255),
.A2(n_696),
.B(n_694),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3404),
.Y(n_3618)
);

OAI21x1_ASAP7_75t_L g3619 ( 
.A1(n_3353),
.A2(n_698),
.B(n_697),
.Y(n_3619)
);

OAI21xp5_ASAP7_75t_L g3620 ( 
.A1(n_3209),
.A2(n_337),
.B(n_340),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3362),
.Y(n_3621)
);

NOR2xp33_ASAP7_75t_SL g3622 ( 
.A(n_3173),
.B(n_343),
.Y(n_3622)
);

AOI22xp33_ASAP7_75t_L g3623 ( 
.A1(n_3195),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_3623)
);

OAI21x1_ASAP7_75t_L g3624 ( 
.A1(n_3383),
.A2(n_700),
.B(n_699),
.Y(n_3624)
);

AOI22xp33_ASAP7_75t_SL g3625 ( 
.A1(n_3195),
.A2(n_3196),
.B1(n_3236),
.B2(n_3229),
.Y(n_3625)
);

AO21x2_ASAP7_75t_L g3626 ( 
.A1(n_3309),
.A2(n_344),
.B(n_345),
.Y(n_3626)
);

OAI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_3310),
.A2(n_346),
.B(n_347),
.Y(n_3627)
);

O2A1O1Ixp33_ASAP7_75t_SL g3628 ( 
.A1(n_3385),
.A2(n_348),
.B(n_346),
.C(n_347),
.Y(n_3628)
);

OAI21x1_ASAP7_75t_L g3629 ( 
.A1(n_3400),
.A2(n_707),
.B(n_706),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3408),
.Y(n_3630)
);

OA21x2_ASAP7_75t_L g3631 ( 
.A1(n_3255),
.A2(n_709),
.B(n_708),
.Y(n_3631)
);

INVx2_ASAP7_75t_L g3632 ( 
.A(n_3219),
.Y(n_3632)
);

OAI21x1_ASAP7_75t_L g3633 ( 
.A1(n_3339),
.A2(n_713),
.B(n_710),
.Y(n_3633)
);

OA21x2_ASAP7_75t_L g3634 ( 
.A1(n_3276),
.A2(n_716),
.B(n_714),
.Y(n_3634)
);

OAI22xp33_ASAP7_75t_L g3635 ( 
.A1(n_3169),
.A2(n_351),
.B1(n_349),
.B2(n_350),
.Y(n_3635)
);

NAND2xp33_ASAP7_75t_L g3636 ( 
.A(n_3116),
.B(n_350),
.Y(n_3636)
);

NAND2xp33_ASAP7_75t_L g3637 ( 
.A(n_3116),
.B(n_351),
.Y(n_3637)
);

OAI21x1_ASAP7_75t_SL g3638 ( 
.A1(n_3334),
.A2(n_352),
.B(n_353),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_3184),
.B(n_353),
.Y(n_3639)
);

BUFx6f_ASAP7_75t_L g3640 ( 
.A(n_3235),
.Y(n_3640)
);

OAI21x1_ASAP7_75t_L g3641 ( 
.A1(n_3360),
.A2(n_720),
.B(n_719),
.Y(n_3641)
);

INVx2_ASAP7_75t_L g3642 ( 
.A(n_3279),
.Y(n_3642)
);

NAND2x1p5_ASAP7_75t_L g3643 ( 
.A(n_3343),
.B(n_355),
.Y(n_3643)
);

AND2x4_ASAP7_75t_L g3644 ( 
.A(n_3416),
.B(n_355),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3301),
.Y(n_3645)
);

OAI21x1_ASAP7_75t_L g3646 ( 
.A1(n_3156),
.A2(n_723),
.B(n_721),
.Y(n_3646)
);

INVx2_ASAP7_75t_L g3647 ( 
.A(n_3235),
.Y(n_3647)
);

NOR2xp67_ASAP7_75t_L g3648 ( 
.A(n_3177),
.B(n_356),
.Y(n_3648)
);

OAI21x1_ASAP7_75t_L g3649 ( 
.A1(n_3292),
.A2(n_725),
.B(n_724),
.Y(n_3649)
);

OA21x2_ASAP7_75t_L g3650 ( 
.A1(n_3276),
.A2(n_730),
.B(n_726),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3196),
.Y(n_3651)
);

OAI22xp5_ASAP7_75t_L g3652 ( 
.A1(n_3169),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3212),
.Y(n_3653)
);

OAI21x1_ASAP7_75t_L g3654 ( 
.A1(n_3296),
.A2(n_3234),
.B(n_3210),
.Y(n_3654)
);

OAI21x1_ASAP7_75t_SL g3655 ( 
.A1(n_3326),
.A2(n_357),
.B(n_358),
.Y(n_3655)
);

AND2x4_ASAP7_75t_L g3656 ( 
.A(n_3416),
.B(n_3241),
.Y(n_3656)
);

OAI21x1_ASAP7_75t_L g3657 ( 
.A1(n_3390),
.A2(n_732),
.B(n_731),
.Y(n_3657)
);

A2O1A1Ixp33_ASAP7_75t_L g3658 ( 
.A1(n_3412),
.A2(n_361),
.B(n_359),
.C(n_360),
.Y(n_3658)
);

OAI21xp5_ASAP7_75t_L g3659 ( 
.A1(n_3261),
.A2(n_360),
.B(n_363),
.Y(n_3659)
);

NAND2x1p5_ASAP7_75t_L g3660 ( 
.A(n_3258),
.B(n_364),
.Y(n_3660)
);

OAI21x1_ASAP7_75t_L g3661 ( 
.A1(n_3269),
.A2(n_3168),
.B(n_3118),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3147),
.Y(n_3662)
);

OAI22xp33_ASAP7_75t_SL g3663 ( 
.A1(n_3575),
.A2(n_3252),
.B1(n_3212),
.B2(n_3226),
.Y(n_3663)
);

BUFx2_ASAP7_75t_L g3664 ( 
.A(n_3493),
.Y(n_3664)
);

OAI21xp5_ASAP7_75t_L g3665 ( 
.A1(n_3443),
.A2(n_3244),
.B(n_3221),
.Y(n_3665)
);

OR2x6_ASAP7_75t_L g3666 ( 
.A(n_3484),
.B(n_3403),
.Y(n_3666)
);

CKINVDCx20_ASAP7_75t_R g3667 ( 
.A(n_3609),
.Y(n_3667)
);

OAI22xp5_ASAP7_75t_SL g3668 ( 
.A1(n_3505),
.A2(n_3183),
.B1(n_3149),
.B2(n_3262),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3515),
.Y(n_3669)
);

AOI22xp33_ASAP7_75t_SL g3670 ( 
.A1(n_3448),
.A2(n_3236),
.B1(n_3229),
.B2(n_3226),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3501),
.Y(n_3671)
);

AND2x4_ASAP7_75t_SL g3672 ( 
.A(n_3585),
.B(n_3178),
.Y(n_3672)
);

CKINVDCx5p33_ASAP7_75t_R g3673 ( 
.A(n_3613),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3501),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3502),
.Y(n_3675)
);

AOI21xp33_ASAP7_75t_L g3676 ( 
.A1(n_3461),
.A2(n_3349),
.B(n_3217),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3502),
.Y(n_3677)
);

OAI21x1_ASAP7_75t_L g3678 ( 
.A1(n_3425),
.A2(n_3335),
.B(n_3145),
.Y(n_3678)
);

AND2x4_ASAP7_75t_L g3679 ( 
.A(n_3585),
.B(n_3217),
.Y(n_3679)
);

CKINVDCx8_ASAP7_75t_R g3680 ( 
.A(n_3556),
.Y(n_3680)
);

AND2x2_ASAP7_75t_L g3681 ( 
.A(n_3522),
.B(n_3283),
.Y(n_3681)
);

INVx2_ASAP7_75t_L g3682 ( 
.A(n_3530),
.Y(n_3682)
);

AND2x4_ASAP7_75t_L g3683 ( 
.A(n_3554),
.B(n_3283),
.Y(n_3683)
);

AOI22xp5_ASAP7_75t_L g3684 ( 
.A1(n_3420),
.A2(n_3191),
.B1(n_3126),
.B2(n_3350),
.Y(n_3684)
);

AND2x4_ASAP7_75t_L g3685 ( 
.A(n_3656),
.B(n_3284),
.Y(n_3685)
);

AND2x4_ASAP7_75t_L g3686 ( 
.A(n_3656),
.B(n_3284),
.Y(n_3686)
);

CKINVDCx11_ASAP7_75t_R g3687 ( 
.A(n_3441),
.Y(n_3687)
);

AND2x4_ASAP7_75t_L g3688 ( 
.A(n_3651),
.B(n_3342),
.Y(n_3688)
);

AOI221xp5_ASAP7_75t_L g3689 ( 
.A1(n_3582),
.A2(n_3312),
.B1(n_3290),
.B2(n_3240),
.C(n_3225),
.Y(n_3689)
);

OAI22xp5_ASAP7_75t_L g3690 ( 
.A1(n_3451),
.A2(n_3170),
.B1(n_3247),
.B2(n_3241),
.Y(n_3690)
);

INVxp67_ASAP7_75t_L g3691 ( 
.A(n_3597),
.Y(n_3691)
);

A2O1A1Ixp33_ASAP7_75t_L g3692 ( 
.A1(n_3627),
.A2(n_3158),
.B(n_3127),
.C(n_3247),
.Y(n_3692)
);

AOI221xp5_ASAP7_75t_L g3693 ( 
.A1(n_3459),
.A2(n_3225),
.B1(n_3322),
.B2(n_3158),
.C(n_3127),
.Y(n_3693)
);

OR2x2_ASAP7_75t_L g3694 ( 
.A(n_3424),
.B(n_3170),
.Y(n_3694)
);

NAND2xp33_ASAP7_75t_SL g3695 ( 
.A(n_3534),
.B(n_3545),
.Y(n_3695)
);

OAI221xp5_ASAP7_75t_L g3696 ( 
.A1(n_3449),
.A2(n_3216),
.B1(n_3282),
.B2(n_3239),
.C(n_3342),
.Y(n_3696)
);

AND2x2_ASAP7_75t_L g3697 ( 
.A(n_3537),
.B(n_3344),
.Y(n_3697)
);

AND2x2_ASAP7_75t_L g3698 ( 
.A(n_3662),
.B(n_3344),
.Y(n_3698)
);

OR2x2_ASAP7_75t_L g3699 ( 
.A(n_3457),
.B(n_3632),
.Y(n_3699)
);

OAI21xp33_ASAP7_75t_SL g3700 ( 
.A1(n_3506),
.A2(n_3288),
.B(n_3270),
.Y(n_3700)
);

AOI22xp33_ASAP7_75t_L g3701 ( 
.A1(n_3444),
.A2(n_3256),
.B1(n_3270),
.B2(n_3288),
.Y(n_3701)
);

AOI22xp33_ASAP7_75t_L g3702 ( 
.A1(n_3447),
.A2(n_3256),
.B1(n_3273),
.B2(n_3393),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3645),
.B(n_3347),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_3645),
.B(n_3347),
.Y(n_3704)
);

AND2x2_ASAP7_75t_L g3705 ( 
.A(n_3480),
.B(n_3531),
.Y(n_3705)
);

AND2x2_ASAP7_75t_L g3706 ( 
.A(n_3642),
.B(n_3363),
.Y(n_3706)
);

BUFx4f_ASAP7_75t_SL g3707 ( 
.A(n_3613),
.Y(n_3707)
);

OAI22xp33_ASAP7_75t_SL g3708 ( 
.A1(n_3622),
.A2(n_3363),
.B1(n_3368),
.B2(n_3273),
.Y(n_3708)
);

AOI22xp33_ASAP7_75t_SL g3709 ( 
.A1(n_3482),
.A2(n_3368),
.B1(n_3315),
.B2(n_3351),
.Y(n_3709)
);

HB1xp67_ASAP7_75t_L g3710 ( 
.A(n_3460),
.Y(n_3710)
);

AOI22xp33_ASAP7_75t_L g3711 ( 
.A1(n_3479),
.A2(n_3462),
.B1(n_3446),
.B2(n_3521),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3508),
.Y(n_3712)
);

INVx2_ASAP7_75t_L g3713 ( 
.A(n_3546),
.Y(n_3713)
);

AOI22xp5_ASAP7_75t_L g3714 ( 
.A1(n_3565),
.A2(n_3346),
.B1(n_3315),
.B2(n_3337),
.Y(n_3714)
);

INVx2_ASAP7_75t_SL g3715 ( 
.A(n_3550),
.Y(n_3715)
);

AOI21x1_ASAP7_75t_L g3716 ( 
.A1(n_3549),
.A2(n_3351),
.B(n_3337),
.Y(n_3716)
);

OAI22xp5_ASAP7_75t_L g3717 ( 
.A1(n_3595),
.A2(n_3648),
.B1(n_3513),
.B2(n_3659),
.Y(n_3717)
);

OAI21x1_ASAP7_75t_L g3718 ( 
.A1(n_3452),
.A2(n_3325),
.B(n_3313),
.Y(n_3718)
);

AOI22xp5_ASAP7_75t_L g3719 ( 
.A1(n_3635),
.A2(n_3392),
.B1(n_3216),
.B2(n_3391),
.Y(n_3719)
);

NAND2xp33_ASAP7_75t_R g3720 ( 
.A(n_3492),
.B(n_364),
.Y(n_3720)
);

BUFx4f_ASAP7_75t_SL g3721 ( 
.A(n_3608),
.Y(n_3721)
);

AOI22xp33_ASAP7_75t_L g3722 ( 
.A1(n_3536),
.A2(n_3391),
.B1(n_3388),
.B2(n_3325),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3508),
.Y(n_3723)
);

INVx1_ASAP7_75t_SL g3724 ( 
.A(n_3540),
.Y(n_3724)
);

AND2x2_ASAP7_75t_L g3725 ( 
.A(n_3454),
.B(n_3388),
.Y(n_3725)
);

INVx2_ASAP7_75t_L g3726 ( 
.A(n_3571),
.Y(n_3726)
);

BUFx2_ASAP7_75t_L g3727 ( 
.A(n_3599),
.Y(n_3727)
);

AOI22xp33_ASAP7_75t_L g3728 ( 
.A1(n_3620),
.A2(n_3594),
.B1(n_3434),
.B2(n_3652),
.Y(n_3728)
);

INVx2_ASAP7_75t_L g3729 ( 
.A(n_3576),
.Y(n_3729)
);

OAI22xp33_ASAP7_75t_L g3730 ( 
.A1(n_3660),
.A2(n_3325),
.B1(n_3377),
.B2(n_3313),
.Y(n_3730)
);

AND2x2_ASAP7_75t_L g3731 ( 
.A(n_3456),
.B(n_3313),
.Y(n_3731)
);

INVx2_ASAP7_75t_L g3732 ( 
.A(n_3589),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3510),
.Y(n_3733)
);

CKINVDCx6p67_ASAP7_75t_R g3734 ( 
.A(n_3644),
.Y(n_3734)
);

AOI22xp33_ASAP7_75t_L g3735 ( 
.A1(n_3594),
.A2(n_3377),
.B1(n_3278),
.B2(n_3369),
.Y(n_3735)
);

OAI22xp5_ASAP7_75t_L g3736 ( 
.A1(n_3625),
.A2(n_3377),
.B1(n_3278),
.B2(n_3369),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3510),
.Y(n_3737)
);

OR2x2_ASAP7_75t_L g3738 ( 
.A(n_3450),
.B(n_3265),
.Y(n_3738)
);

OAI22xp5_ASAP7_75t_L g3739 ( 
.A1(n_3643),
.A2(n_3407),
.B1(n_3371),
.B2(n_3265),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3512),
.Y(n_3740)
);

AOI22xp33_ASAP7_75t_L g3741 ( 
.A1(n_3511),
.A2(n_3488),
.B1(n_3644),
.B2(n_3593),
.Y(n_3741)
);

O2A1O1Ixp33_ASAP7_75t_L g3742 ( 
.A1(n_3435),
.A2(n_367),
.B(n_365),
.C(n_366),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3512),
.Y(n_3743)
);

AND2x2_ASAP7_75t_SL g3744 ( 
.A(n_3469),
.B(n_3371),
.Y(n_3744)
);

AOI21xp33_ASAP7_75t_L g3745 ( 
.A1(n_3473),
.A2(n_3495),
.B(n_3525),
.Y(n_3745)
);

OAI21xp5_ASAP7_75t_L g3746 ( 
.A1(n_3529),
.A2(n_365),
.B(n_366),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3463),
.Y(n_3747)
);

AOI21xp5_ASAP7_75t_SL g3748 ( 
.A1(n_3458),
.A2(n_3407),
.B(n_368),
.Y(n_3748)
);

AND2x4_ASAP7_75t_L g3749 ( 
.A(n_3651),
.B(n_369),
.Y(n_3749)
);

OAI21xp5_ASAP7_75t_L g3750 ( 
.A1(n_3590),
.A2(n_369),
.B(n_370),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3517),
.Y(n_3751)
);

NAND3xp33_ASAP7_75t_L g3752 ( 
.A(n_3473),
.B(n_370),
.C(n_371),
.Y(n_3752)
);

OAI21x1_ASAP7_75t_L g3753 ( 
.A1(n_3472),
.A2(n_736),
.B(n_733),
.Y(n_3753)
);

OAI22xp5_ASAP7_75t_L g3754 ( 
.A1(n_3593),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_3754)
);

AOI22xp33_ASAP7_75t_SL g3755 ( 
.A1(n_3482),
.A2(n_376),
.B1(n_373),
.B2(n_374),
.Y(n_3755)
);

INVxp67_ASAP7_75t_SL g3756 ( 
.A(n_3563),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3551),
.Y(n_3757)
);

NAND2xp33_ASAP7_75t_R g3758 ( 
.A(n_3562),
.B(n_3458),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3555),
.Y(n_3759)
);

CKINVDCx11_ASAP7_75t_R g3760 ( 
.A(n_3433),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3591),
.B(n_377),
.Y(n_3761)
);

NOR2xp33_ASAP7_75t_L g3762 ( 
.A(n_3486),
.B(n_377),
.Y(n_3762)
);

INVx2_ASAP7_75t_L g3763 ( 
.A(n_3601),
.Y(n_3763)
);

AOI21xp5_ASAP7_75t_L g3764 ( 
.A1(n_3539),
.A2(n_378),
.B(n_379),
.Y(n_3764)
);

NOR3xp33_ASAP7_75t_SL g3765 ( 
.A(n_3494),
.B(n_379),
.C(n_380),
.Y(n_3765)
);

NAND2x1p5_ASAP7_75t_L g3766 ( 
.A(n_3504),
.B(n_3570),
.Y(n_3766)
);

AND2x4_ASAP7_75t_L g3767 ( 
.A(n_3653),
.B(n_380),
.Y(n_3767)
);

AOI22x1_ASAP7_75t_L g3768 ( 
.A1(n_3586),
.A2(n_383),
.B1(n_381),
.B2(n_382),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3606),
.Y(n_3769)
);

A2O1A1Ixp33_ASAP7_75t_L g3770 ( 
.A1(n_3658),
.A2(n_384),
.B(n_381),
.C(n_382),
.Y(n_3770)
);

AOI22xp33_ASAP7_75t_L g3771 ( 
.A1(n_3604),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_3771)
);

OR2x6_ASAP7_75t_L g3772 ( 
.A(n_3654),
.B(n_387),
.Y(n_3772)
);

OR2x6_ASAP7_75t_L g3773 ( 
.A(n_3541),
.B(n_387),
.Y(n_3773)
);

AOI22xp33_ASAP7_75t_L g3774 ( 
.A1(n_3466),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_3774)
);

AOI221xp5_ASAP7_75t_L g3775 ( 
.A1(n_3543),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.C(n_391),
.Y(n_3775)
);

AOI22xp33_ASAP7_75t_SL g3776 ( 
.A1(n_3548),
.A2(n_394),
.B1(n_391),
.B2(n_392),
.Y(n_3776)
);

CKINVDCx16_ASAP7_75t_R g3777 ( 
.A(n_3430),
.Y(n_3777)
);

AOI22xp33_ASAP7_75t_L g3778 ( 
.A1(n_3611),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_3778)
);

NAND2xp33_ASAP7_75t_SL g3779 ( 
.A(n_3440),
.B(n_395),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3602),
.B(n_397),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3421),
.Y(n_3781)
);

INVx1_ASAP7_75t_L g3782 ( 
.A(n_3568),
.Y(n_3782)
);

AO21x2_ASAP7_75t_L g3783 ( 
.A1(n_3535),
.A2(n_397),
.B(n_398),
.Y(n_3783)
);

AOI22xp33_ASAP7_75t_L g3784 ( 
.A1(n_3592),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3524),
.B(n_3455),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3591),
.B(n_399),
.Y(n_3786)
);

BUFx2_ASAP7_75t_L g3787 ( 
.A(n_3560),
.Y(n_3787)
);

INVx2_ASAP7_75t_L g3788 ( 
.A(n_3485),
.Y(n_3788)
);

OAI22xp5_ASAP7_75t_L g3789 ( 
.A1(n_3615),
.A2(n_404),
.B1(n_400),
.B2(n_401),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_3603),
.B(n_401),
.Y(n_3790)
);

AOI22xp33_ASAP7_75t_L g3791 ( 
.A1(n_3567),
.A2(n_408),
.B1(n_404),
.B2(n_407),
.Y(n_3791)
);

OAI21x1_ASAP7_75t_L g3792 ( 
.A1(n_3464),
.A2(n_741),
.B(n_738),
.Y(n_3792)
);

AOI22xp33_ASAP7_75t_SL g3793 ( 
.A1(n_3616),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_3793)
);

AOI22xp33_ASAP7_75t_SL g3794 ( 
.A1(n_3616),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_3794)
);

INVx1_ASAP7_75t_SL g3795 ( 
.A(n_3538),
.Y(n_3795)
);

AOI22xp33_ASAP7_75t_L g3796 ( 
.A1(n_3588),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.Y(n_3796)
);

OA21x2_ASAP7_75t_L g3797 ( 
.A1(n_3509),
.A2(n_412),
.B(n_413),
.Y(n_3797)
);

OAI21x1_ASAP7_75t_SL g3798 ( 
.A1(n_3638),
.A2(n_413),
.B(n_414),
.Y(n_3798)
);

OAI211xp5_ASAP7_75t_L g3799 ( 
.A1(n_3581),
.A2(n_416),
.B(n_414),
.C(n_415),
.Y(n_3799)
);

AOI22x1_ASAP7_75t_L g3800 ( 
.A1(n_3440),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_3800)
);

OR2x2_ASAP7_75t_L g3801 ( 
.A(n_3621),
.B(n_419),
.Y(n_3801)
);

AOI22xp33_ASAP7_75t_L g3802 ( 
.A1(n_3574),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.Y(n_3802)
);

NOR4xp25_ASAP7_75t_L g3803 ( 
.A(n_3639),
.B(n_423),
.C(n_420),
.D(n_422),
.Y(n_3803)
);

BUFx3_ASAP7_75t_L g3804 ( 
.A(n_3433),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_3621),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3427),
.Y(n_3806)
);

INVx3_ASAP7_75t_L g3807 ( 
.A(n_3468),
.Y(n_3807)
);

AOI221xp5_ASAP7_75t_L g3808 ( 
.A1(n_3573),
.A2(n_3499),
.B1(n_3422),
.B2(n_3558),
.C(n_3519),
.Y(n_3808)
);

AOI22xp33_ASAP7_75t_SL g3809 ( 
.A1(n_3631),
.A2(n_3650),
.B1(n_3634),
.B2(n_3468),
.Y(n_3809)
);

AND2x4_ASAP7_75t_L g3810 ( 
.A(n_3653),
.B(n_424),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3427),
.Y(n_3811)
);

OAI22xp5_ASAP7_75t_L g3812 ( 
.A1(n_3623),
.A2(n_427),
.B1(n_425),
.B2(n_426),
.Y(n_3812)
);

OR2x6_ASAP7_75t_L g3813 ( 
.A(n_3503),
.B(n_3655),
.Y(n_3813)
);

OR2x2_ASAP7_75t_L g3814 ( 
.A(n_3630),
.B(n_428),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3428),
.Y(n_3815)
);

BUFx6f_ASAP7_75t_L g3816 ( 
.A(n_3433),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3428),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3437),
.Y(n_3818)
);

INVx2_ASAP7_75t_L g3819 ( 
.A(n_3630),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3603),
.B(n_428),
.Y(n_3820)
);

OAI22xp33_ASAP7_75t_L g3821 ( 
.A1(n_3631),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.Y(n_3821)
);

AND2x2_ASAP7_75t_L g3822 ( 
.A(n_3607),
.B(n_430),
.Y(n_3822)
);

HB1xp67_ASAP7_75t_L g3823 ( 
.A(n_3661),
.Y(n_3823)
);

INVx2_ASAP7_75t_SL g3824 ( 
.A(n_3528),
.Y(n_3824)
);

AO21x2_ASAP7_75t_L g3825 ( 
.A1(n_3557),
.A2(n_432),
.B(n_433),
.Y(n_3825)
);

INVx2_ASAP7_75t_SL g3826 ( 
.A(n_3528),
.Y(n_3826)
);

AOI22xp33_ASAP7_75t_SL g3827 ( 
.A1(n_3634),
.A2(n_436),
.B1(n_432),
.B2(n_434),
.Y(n_3827)
);

AND2x2_ASAP7_75t_L g3828 ( 
.A(n_3607),
.B(n_434),
.Y(n_3828)
);

NAND3xp33_ASAP7_75t_SL g3829 ( 
.A(n_3514),
.B(n_437),
.C(n_438),
.Y(n_3829)
);

NAND2xp33_ASAP7_75t_R g3830 ( 
.A(n_3765),
.B(n_3650),
.Y(n_3830)
);

INVx3_ASAP7_75t_L g3831 ( 
.A(n_3807),
.Y(n_3831)
);

INVx2_ASAP7_75t_L g3832 ( 
.A(n_3664),
.Y(n_3832)
);

A2O1A1Ixp33_ASAP7_75t_L g3833 ( 
.A1(n_3700),
.A2(n_3637),
.B(n_3636),
.C(n_3474),
.Y(n_3833)
);

CKINVDCx5p33_ASAP7_75t_R g3834 ( 
.A(n_3687),
.Y(n_3834)
);

BUFx2_ASAP7_75t_SL g3835 ( 
.A(n_3724),
.Y(n_3835)
);

OAI22xp33_ASAP7_75t_SL g3836 ( 
.A1(n_3666),
.A2(n_3618),
.B1(n_3559),
.B2(n_3491),
.Y(n_3836)
);

NOR2xp33_ASAP7_75t_R g3837 ( 
.A(n_3707),
.B(n_3673),
.Y(n_3837)
);

INVx3_ASAP7_75t_L g3838 ( 
.A(n_3807),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3747),
.Y(n_3839)
);

AOI22xp33_ASAP7_75t_L g3840 ( 
.A1(n_3711),
.A2(n_3442),
.B1(n_3600),
.B2(n_3523),
.Y(n_3840)
);

AND2x2_ASAP7_75t_L g3841 ( 
.A(n_3697),
.B(n_3437),
.Y(n_3841)
);

INVx2_ASAP7_75t_L g3842 ( 
.A(n_3785),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3751),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_3710),
.B(n_3618),
.Y(n_3844)
);

INVxp67_ASAP7_75t_L g3845 ( 
.A(n_3715),
.Y(n_3845)
);

NOR2xp33_ASAP7_75t_L g3846 ( 
.A(n_3777),
.B(n_3544),
.Y(n_3846)
);

AO21x1_ASAP7_75t_L g3847 ( 
.A1(n_3663),
.A2(n_3491),
.B(n_3470),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3699),
.B(n_3439),
.Y(n_3848)
);

INVx3_ASAP7_75t_L g3849 ( 
.A(n_3679),
.Y(n_3849)
);

CKINVDCx16_ASAP7_75t_R g3850 ( 
.A(n_3667),
.Y(n_3850)
);

CKINVDCx8_ASAP7_75t_R g3851 ( 
.A(n_3666),
.Y(n_3851)
);

OAI21xp5_ASAP7_75t_SL g3852 ( 
.A1(n_3693),
.A2(n_3503),
.B(n_3561),
.Y(n_3852)
);

OR2x2_ASAP7_75t_L g3853 ( 
.A(n_3681),
.B(n_3439),
.Y(n_3853)
);

AND2x4_ASAP7_75t_L g3854 ( 
.A(n_3683),
.B(n_3470),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3805),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3806),
.Y(n_3856)
);

INVx2_ASAP7_75t_L g3857 ( 
.A(n_3819),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3757),
.Y(n_3858)
);

HB1xp67_ASAP7_75t_L g3859 ( 
.A(n_3691),
.Y(n_3859)
);

INVx2_ASAP7_75t_L g3860 ( 
.A(n_3669),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3705),
.B(n_3476),
.Y(n_3861)
);

CKINVDCx20_ASAP7_75t_R g3862 ( 
.A(n_3721),
.Y(n_3862)
);

OAI22xp5_ASAP7_75t_L g3863 ( 
.A1(n_3734),
.A2(n_3560),
.B1(n_3547),
.B2(n_3572),
.Y(n_3863)
);

OR2x6_ASAP7_75t_L g3864 ( 
.A(n_3813),
.B(n_3528),
.Y(n_3864)
);

AND2x2_ASAP7_75t_L g3865 ( 
.A(n_3756),
.B(n_3476),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3759),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3682),
.Y(n_3867)
);

OAI21xp33_ASAP7_75t_L g3868 ( 
.A1(n_3741),
.A2(n_3578),
.B(n_3569),
.Y(n_3868)
);

AND2x2_ASAP7_75t_L g3869 ( 
.A(n_3679),
.B(n_3487),
.Y(n_3869)
);

INVx3_ASAP7_75t_L g3870 ( 
.A(n_3744),
.Y(n_3870)
);

INVx2_ASAP7_75t_SL g3871 ( 
.A(n_3672),
.Y(n_3871)
);

BUFx4f_ASAP7_75t_SL g3872 ( 
.A(n_3694),
.Y(n_3872)
);

CKINVDCx5p33_ASAP7_75t_R g3873 ( 
.A(n_3680),
.Y(n_3873)
);

OR2x2_ASAP7_75t_SL g3874 ( 
.A(n_3758),
.B(n_3516),
.Y(n_3874)
);

AND2x2_ASAP7_75t_L g3875 ( 
.A(n_3683),
.B(n_3487),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3713),
.Y(n_3876)
);

BUFx4f_ASAP7_75t_SL g3877 ( 
.A(n_3727),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3782),
.Y(n_3878)
);

INVxp67_ASAP7_75t_L g3879 ( 
.A(n_3720),
.Y(n_3879)
);

AND2x2_ASAP7_75t_L g3880 ( 
.A(n_3706),
.B(n_3490),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3671),
.Y(n_3881)
);

AO31x2_ASAP7_75t_L g3882 ( 
.A1(n_3736),
.A2(n_3692),
.A3(n_3690),
.B(n_3787),
.Y(n_3882)
);

CKINVDCx20_ASAP7_75t_R g3883 ( 
.A(n_3668),
.Y(n_3883)
);

NOR2xp67_ASAP7_75t_L g3884 ( 
.A(n_3696),
.B(n_3532),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3674),
.Y(n_3885)
);

NOR2xp33_ASAP7_75t_R g3886 ( 
.A(n_3695),
.B(n_438),
.Y(n_3886)
);

OR2x6_ASAP7_75t_L g3887 ( 
.A(n_3813),
.B(n_3445),
.Y(n_3887)
);

CKINVDCx16_ASAP7_75t_R g3888 ( 
.A(n_3684),
.Y(n_3888)
);

AND2x4_ASAP7_75t_L g3889 ( 
.A(n_3688),
.B(n_3490),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_3675),
.B(n_3431),
.Y(n_3890)
);

OR2x2_ASAP7_75t_L g3891 ( 
.A(n_3726),
.B(n_3467),
.Y(n_3891)
);

BUFx3_ASAP7_75t_L g3892 ( 
.A(n_3766),
.Y(n_3892)
);

AOI221xp5_ASAP7_75t_L g3893 ( 
.A1(n_3803),
.A2(n_3628),
.B1(n_3500),
.B2(n_3478),
.C(n_3626),
.Y(n_3893)
);

OAI21x1_ASAP7_75t_L g3894 ( 
.A1(n_3716),
.A2(n_3527),
.B(n_3465),
.Y(n_3894)
);

AND2x2_ASAP7_75t_L g3895 ( 
.A(n_3725),
.B(n_3516),
.Y(n_3895)
);

OR2x2_ASAP7_75t_L g3896 ( 
.A(n_3729),
.B(n_3583),
.Y(n_3896)
);

BUFx6f_ASAP7_75t_L g3897 ( 
.A(n_3816),
.Y(n_3897)
);

NAND3xp33_ASAP7_75t_L g3898 ( 
.A(n_3745),
.B(n_3442),
.C(n_3577),
.Y(n_3898)
);

HB1xp67_ASAP7_75t_L g3899 ( 
.A(n_3732),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3677),
.Y(n_3900)
);

NOR2xp33_ASAP7_75t_R g3901 ( 
.A(n_3760),
.B(n_439),
.Y(n_3901)
);

NAND2xp33_ASAP7_75t_R g3902 ( 
.A(n_3773),
.B(n_3605),
.Y(n_3902)
);

INVx2_ASAP7_75t_L g3903 ( 
.A(n_3763),
.Y(n_3903)
);

AND2x2_ASAP7_75t_L g3904 ( 
.A(n_3698),
.B(n_3542),
.Y(n_3904)
);

XOR2xp5_ASAP7_75t_L g3905 ( 
.A(n_3738),
.B(n_3566),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3769),
.Y(n_3906)
);

AND2x4_ASAP7_75t_L g3907 ( 
.A(n_3688),
.B(n_3542),
.Y(n_3907)
);

INVx3_ASAP7_75t_L g3908 ( 
.A(n_3685),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3712),
.B(n_3614),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3723),
.Y(n_3910)
);

INVx2_ASAP7_75t_L g3911 ( 
.A(n_3781),
.Y(n_3911)
);

OR2x6_ASAP7_75t_L g3912 ( 
.A(n_3748),
.B(n_3518),
.Y(n_3912)
);

OR2x2_ASAP7_75t_L g3913 ( 
.A(n_3842),
.B(n_3733),
.Y(n_3913)
);

OR2x6_ASAP7_75t_L g3914 ( 
.A(n_3887),
.B(n_3772),
.Y(n_3914)
);

BUFx6f_ASAP7_75t_L g3915 ( 
.A(n_3897),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_3896),
.Y(n_3916)
);

OA21x2_ASAP7_75t_L g3917 ( 
.A1(n_3894),
.A2(n_3752),
.B(n_3823),
.Y(n_3917)
);

INVxp67_ASAP7_75t_SL g3918 ( 
.A(n_3899),
.Y(n_3918)
);

AND2x2_ASAP7_75t_L g3919 ( 
.A(n_3895),
.B(n_3869),
.Y(n_3919)
);

AND2x2_ASAP7_75t_L g3920 ( 
.A(n_3875),
.B(n_3737),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3856),
.Y(n_3921)
);

AND2x2_ASAP7_75t_L g3922 ( 
.A(n_3841),
.B(n_3740),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3856),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3855),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3839),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3843),
.Y(n_3926)
);

AND2x2_ASAP7_75t_L g3927 ( 
.A(n_3861),
.B(n_3743),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3881),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3880),
.B(n_3811),
.Y(n_3929)
);

INVx2_ASAP7_75t_L g3930 ( 
.A(n_3857),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3885),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3889),
.B(n_3815),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3900),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3865),
.B(n_3817),
.Y(n_3934)
);

NOR2xp33_ASAP7_75t_L g3935 ( 
.A(n_3851),
.B(n_3665),
.Y(n_3935)
);

INVx2_ASAP7_75t_L g3936 ( 
.A(n_3860),
.Y(n_3936)
);

AND2x2_ASAP7_75t_L g3937 ( 
.A(n_3889),
.B(n_3818),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3910),
.Y(n_3938)
);

CKINVDCx5p33_ASAP7_75t_R g3939 ( 
.A(n_3837),
.Y(n_3939)
);

HB1xp67_ASAP7_75t_L g3940 ( 
.A(n_3832),
.Y(n_3940)
);

BUFx3_ASAP7_75t_L g3941 ( 
.A(n_3871),
.Y(n_3941)
);

INVx2_ASAP7_75t_L g3942 ( 
.A(n_3867),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3876),
.Y(n_3943)
);

INVx2_ASAP7_75t_L g3944 ( 
.A(n_3903),
.Y(n_3944)
);

AND2x2_ASAP7_75t_L g3945 ( 
.A(n_3854),
.B(n_3849),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3858),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3866),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3906),
.Y(n_3948)
);

AND2x2_ASAP7_75t_L g3949 ( 
.A(n_3854),
.B(n_3788),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3878),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3844),
.Y(n_3951)
);

AND2x2_ASAP7_75t_L g3952 ( 
.A(n_3849),
.B(n_3809),
.Y(n_3952)
);

INVxp67_ASAP7_75t_L g3953 ( 
.A(n_3835),
.Y(n_3953)
);

INVx2_ASAP7_75t_L g3954 ( 
.A(n_3911),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3848),
.B(n_3808),
.Y(n_3955)
);

INVx2_ASAP7_75t_L g3956 ( 
.A(n_3909),
.Y(n_3956)
);

AND2x4_ASAP7_75t_L g3957 ( 
.A(n_3887),
.B(n_3685),
.Y(n_3957)
);

AND2x2_ASAP7_75t_L g3958 ( 
.A(n_3908),
.B(n_3853),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3891),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3890),
.Y(n_3960)
);

INVx2_ASAP7_75t_L g3961 ( 
.A(n_3831),
.Y(n_3961)
);

BUFx2_ASAP7_75t_L g3962 ( 
.A(n_3877),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3859),
.Y(n_3963)
);

AND2x2_ASAP7_75t_L g3964 ( 
.A(n_3908),
.B(n_3797),
.Y(n_3964)
);

BUFx3_ASAP7_75t_L g3965 ( 
.A(n_3892),
.Y(n_3965)
);

INVx2_ASAP7_75t_L g3966 ( 
.A(n_3831),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3847),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3874),
.Y(n_3968)
);

AND2x2_ASAP7_75t_L g3969 ( 
.A(n_3904),
.B(n_3797),
.Y(n_3969)
);

INVx2_ASAP7_75t_L g3970 ( 
.A(n_3838),
.Y(n_3970)
);

INVx2_ASAP7_75t_L g3971 ( 
.A(n_3838),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3836),
.Y(n_3972)
);

BUFx6f_ASAP7_75t_L g3973 ( 
.A(n_3897),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_3864),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3864),
.Y(n_3975)
);

AND2x2_ASAP7_75t_L g3976 ( 
.A(n_3945),
.B(n_3907),
.Y(n_3976)
);

OA211x2_ASAP7_75t_L g3977 ( 
.A1(n_3953),
.A2(n_3879),
.B(n_3689),
.C(n_3845),
.Y(n_3977)
);

AND2x2_ASAP7_75t_L g3978 ( 
.A(n_3945),
.B(n_3919),
.Y(n_3978)
);

OAI22xp5_ASAP7_75t_L g3979 ( 
.A1(n_3914),
.A2(n_3835),
.B1(n_3888),
.B2(n_3872),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_SL g3980 ( 
.A(n_3962),
.B(n_3886),
.Y(n_3980)
);

NAND3xp33_ASAP7_75t_L g3981 ( 
.A(n_3967),
.B(n_3902),
.C(n_3840),
.Y(n_3981)
);

AOI22xp33_ASAP7_75t_L g3982 ( 
.A1(n_3914),
.A2(n_3717),
.B1(n_3884),
.B2(n_3868),
.Y(n_3982)
);

NAND4xp25_ASAP7_75t_L g3983 ( 
.A(n_3935),
.B(n_3714),
.C(n_3701),
.D(n_3830),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_3918),
.B(n_3960),
.Y(n_3984)
);

NAND3xp33_ASAP7_75t_L g3985 ( 
.A(n_3967),
.B(n_3893),
.C(n_3676),
.Y(n_3985)
);

OA21x2_ASAP7_75t_L g3986 ( 
.A1(n_3968),
.A2(n_3852),
.B(n_3898),
.Y(n_3986)
);

OAI221xp5_ASAP7_75t_L g3987 ( 
.A1(n_3914),
.A2(n_3833),
.B1(n_3728),
.B2(n_3863),
.C(n_3670),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3960),
.B(n_3882),
.Y(n_3988)
);

NAND3xp33_ASAP7_75t_L g3989 ( 
.A(n_3972),
.B(n_3846),
.C(n_3794),
.Y(n_3989)
);

NAND3xp33_ASAP7_75t_L g3990 ( 
.A(n_3972),
.B(n_3827),
.C(n_3793),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_L g3991 ( 
.A(n_3969),
.B(n_3882),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_L g3992 ( 
.A(n_3969),
.B(n_3882),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_L g3993 ( 
.A(n_3951),
.B(n_3703),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3956),
.B(n_3704),
.Y(n_3994)
);

OAI22xp5_ASAP7_75t_L g3995 ( 
.A1(n_3914),
.A2(n_3870),
.B1(n_3772),
.B2(n_3883),
.Y(n_3995)
);

AOI21xp5_ASAP7_75t_SL g3996 ( 
.A1(n_3965),
.A2(n_3708),
.B(n_3912),
.Y(n_3996)
);

AOI221xp5_ASAP7_75t_L g3997 ( 
.A1(n_3968),
.A2(n_3742),
.B1(n_3754),
.B2(n_3901),
.C(n_3829),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_L g3998 ( 
.A(n_3952),
.B(n_3907),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_L g3999 ( 
.A(n_3952),
.B(n_3749),
.Y(n_3999)
);

AND2x2_ASAP7_75t_L g4000 ( 
.A(n_3919),
.B(n_3686),
.Y(n_4000)
);

AND2x2_ASAP7_75t_L g4001 ( 
.A(n_3958),
.B(n_3686),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3928),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_L g4003 ( 
.A(n_3959),
.B(n_3749),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_L g4004 ( 
.A(n_3959),
.B(n_3767),
.Y(n_4004)
);

OAI21xp5_ASAP7_75t_SL g4005 ( 
.A1(n_3962),
.A2(n_3870),
.B(n_3755),
.Y(n_4005)
);

AND2x2_ASAP7_75t_L g4006 ( 
.A(n_3958),
.B(n_3905),
.Y(n_4006)
);

AND2x2_ASAP7_75t_L g4007 ( 
.A(n_3932),
.B(n_3937),
.Y(n_4007)
);

AND2x2_ASAP7_75t_L g4008 ( 
.A(n_3932),
.B(n_3850),
.Y(n_4008)
);

NAND3xp33_ASAP7_75t_L g4009 ( 
.A(n_3963),
.B(n_3776),
.C(n_3762),
.Y(n_4009)
);

AND2x2_ASAP7_75t_L g4010 ( 
.A(n_3937),
.B(n_3897),
.Y(n_4010)
);

OAI22xp5_ASAP7_75t_L g4011 ( 
.A1(n_3941),
.A2(n_3773),
.B1(n_3912),
.B2(n_3702),
.Y(n_4011)
);

AND2x2_ASAP7_75t_L g4012 ( 
.A(n_3949),
.B(n_3731),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3927),
.B(n_3767),
.Y(n_4013)
);

OAI221xp5_ASAP7_75t_L g4014 ( 
.A1(n_3955),
.A2(n_3719),
.B1(n_3750),
.B2(n_3722),
.C(n_3746),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_L g4015 ( 
.A(n_3927),
.B(n_3810),
.Y(n_4015)
);

NAND3xp33_ASAP7_75t_L g4016 ( 
.A(n_3974),
.B(n_3802),
.C(n_3796),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_L g4017 ( 
.A(n_3956),
.B(n_3783),
.Y(n_4017)
);

OAI221xp5_ASAP7_75t_L g4018 ( 
.A1(n_3941),
.A2(n_3779),
.B1(n_3768),
.B2(n_3774),
.C(n_3778),
.Y(n_4018)
);

NAND3xp33_ASAP7_75t_L g4019 ( 
.A(n_3974),
.B(n_3764),
.C(n_3800),
.Y(n_4019)
);

OAI21xp5_ASAP7_75t_SL g4020 ( 
.A1(n_3957),
.A2(n_3730),
.B(n_3709),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_3922),
.B(n_3810),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3922),
.B(n_3822),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_3929),
.B(n_3828),
.Y(n_4023)
);

NAND4xp25_ASAP7_75t_SL g4024 ( 
.A(n_3975),
.B(n_3862),
.C(n_3735),
.D(n_3780),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_L g4025 ( 
.A(n_3929),
.B(n_3825),
.Y(n_4025)
);

AND2x2_ASAP7_75t_L g4026 ( 
.A(n_3949),
.B(n_3804),
.Y(n_4026)
);

NAND3xp33_ASAP7_75t_L g4027 ( 
.A(n_3975),
.B(n_3775),
.C(n_3761),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_L g4028 ( 
.A(n_3920),
.B(n_3801),
.Y(n_4028)
);

NAND2xp5_ASAP7_75t_L g4029 ( 
.A(n_3920),
.B(n_3814),
.Y(n_4029)
);

AOI22xp33_ASAP7_75t_L g4030 ( 
.A1(n_3957),
.A2(n_3798),
.B1(n_3821),
.B2(n_3771),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3940),
.B(n_3786),
.Y(n_4031)
);

INVx2_ASAP7_75t_L g4032 ( 
.A(n_3916),
.Y(n_4032)
);

NOR3xp33_ASAP7_75t_SL g4033 ( 
.A(n_3939),
.B(n_3834),
.C(n_3873),
.Y(n_4033)
);

NOR3xp33_ASAP7_75t_L g4034 ( 
.A(n_3964),
.B(n_3799),
.C(n_3739),
.Y(n_4034)
);

AND2x2_ASAP7_75t_L g4035 ( 
.A(n_3957),
.B(n_3824),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_3984),
.Y(n_4036)
);

INVx2_ASAP7_75t_L g4037 ( 
.A(n_4032),
.Y(n_4037)
);

OR2x2_ASAP7_75t_L g4038 ( 
.A(n_3994),
.B(n_3913),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_4002),
.Y(n_4039)
);

AND2x2_ASAP7_75t_L g4040 ( 
.A(n_3978),
.B(n_3965),
.Y(n_4040)
);

OR2x2_ASAP7_75t_L g4041 ( 
.A(n_3994),
.B(n_3913),
.Y(n_4041)
);

AND2x4_ASAP7_75t_L g4042 ( 
.A(n_3981),
.B(n_3964),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_4025),
.B(n_3916),
.Y(n_4043)
);

INVx2_ASAP7_75t_L g4044 ( 
.A(n_4017),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3993),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_4003),
.Y(n_4046)
);

HB1xp67_ASAP7_75t_L g4047 ( 
.A(n_3988),
.Y(n_4047)
);

CKINVDCx16_ASAP7_75t_R g4048 ( 
.A(n_3979),
.Y(n_4048)
);

HB1xp67_ASAP7_75t_L g4049 ( 
.A(n_4017),
.Y(n_4049)
);

AND2x2_ASAP7_75t_L g4050 ( 
.A(n_4007),
.B(n_3961),
.Y(n_4050)
);

NOR2xp33_ASAP7_75t_L g4051 ( 
.A(n_3983),
.B(n_3939),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_4004),
.Y(n_4052)
);

NOR2xp67_ASAP7_75t_L g4053 ( 
.A(n_3979),
.B(n_3961),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_4031),
.Y(n_4054)
);

INVx3_ASAP7_75t_L g4055 ( 
.A(n_3986),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_3985),
.B(n_3928),
.Y(n_4056)
);

HB1xp67_ASAP7_75t_L g4057 ( 
.A(n_3986),
.Y(n_4057)
);

INVx2_ASAP7_75t_SL g4058 ( 
.A(n_4026),
.Y(n_4058)
);

INVx2_ASAP7_75t_L g4059 ( 
.A(n_4012),
.Y(n_4059)
);

INVx2_ASAP7_75t_L g4060 ( 
.A(n_4000),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3998),
.Y(n_4061)
);

AND2x2_ASAP7_75t_L g4062 ( 
.A(n_4010),
.B(n_3966),
.Y(n_4062)
);

OR2x2_ASAP7_75t_L g4063 ( 
.A(n_3991),
.B(n_3934),
.Y(n_4063)
);

INVx2_ASAP7_75t_SL g4064 ( 
.A(n_4035),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_4028),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_3992),
.B(n_3931),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_4029),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_4022),
.Y(n_4068)
);

INVx2_ASAP7_75t_L g4069 ( 
.A(n_4001),
.Y(n_4069)
);

INVxp67_ASAP7_75t_L g4070 ( 
.A(n_3980),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_L g4071 ( 
.A(n_4034),
.B(n_3931),
.Y(n_4071)
);

AND2x2_ASAP7_75t_L g4072 ( 
.A(n_3976),
.B(n_3966),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_4006),
.B(n_3970),
.Y(n_4073)
);

OR2x2_ASAP7_75t_L g4074 ( 
.A(n_4038),
.B(n_3995),
.Y(n_4074)
);

OR2x2_ASAP7_75t_L g4075 ( 
.A(n_4041),
.B(n_3995),
.Y(n_4075)
);

OR2x2_ASAP7_75t_L g4076 ( 
.A(n_4043),
.B(n_4023),
.Y(n_4076)
);

OR2x2_ASAP7_75t_L g4077 ( 
.A(n_4063),
.B(n_3999),
.Y(n_4077)
);

INVx2_ASAP7_75t_SL g4078 ( 
.A(n_4040),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_4048),
.B(n_4008),
.Y(n_4079)
);

AND2x2_ASAP7_75t_L g4080 ( 
.A(n_4070),
.B(n_3982),
.Y(n_4080)
);

INVx2_ASAP7_75t_L g4081 ( 
.A(n_4037),
.Y(n_4081)
);

AND2x2_ASAP7_75t_L g4082 ( 
.A(n_4053),
.B(n_3996),
.Y(n_4082)
);

AND2x2_ASAP7_75t_L g4083 ( 
.A(n_4073),
.B(n_4064),
.Y(n_4083)
);

AND2x2_ASAP7_75t_L g4084 ( 
.A(n_4073),
.B(n_4020),
.Y(n_4084)
);

INVx1_ASAP7_75t_SL g4085 ( 
.A(n_4057),
.Y(n_4085)
);

AND2x2_ASAP7_75t_L g4086 ( 
.A(n_4064),
.B(n_4011),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_4036),
.Y(n_4087)
);

AND2x2_ASAP7_75t_L g4088 ( 
.A(n_4069),
.B(n_4011),
.Y(n_4088)
);

HB1xp67_ASAP7_75t_L g4089 ( 
.A(n_4044),
.Y(n_4089)
);

AND2x4_ASAP7_75t_L g4090 ( 
.A(n_4055),
.B(n_3989),
.Y(n_4090)
);

NAND2x1p5_ASAP7_75t_SL g4091 ( 
.A(n_4044),
.B(n_3977),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_4045),
.Y(n_4092)
);

OR2x2_ASAP7_75t_L g4093 ( 
.A(n_4066),
.B(n_4013),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_4069),
.B(n_4015),
.Y(n_4094)
);

AND2x2_ASAP7_75t_L g4095 ( 
.A(n_4060),
.B(n_4021),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_4049),
.B(n_3933),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_4054),
.Y(n_4097)
);

INVx2_ASAP7_75t_L g4098 ( 
.A(n_4037),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_4039),
.Y(n_4099)
);

AND2x2_ASAP7_75t_SL g4100 ( 
.A(n_4057),
.B(n_4055),
.Y(n_4100)
);

NOR2xp67_ASAP7_75t_L g4101 ( 
.A(n_4055),
.B(n_4024),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_4065),
.Y(n_4102)
);

NAND2x1_ASAP7_75t_SL g4103 ( 
.A(n_4051),
.B(n_4042),
.Y(n_4103)
);

INVxp67_ASAP7_75t_L g4104 ( 
.A(n_4051),
.Y(n_4104)
);

HB1xp67_ASAP7_75t_L g4105 ( 
.A(n_4049),
.Y(n_4105)
);

INVx1_ASAP7_75t_L g4106 ( 
.A(n_4067),
.Y(n_4106)
);

INVx2_ASAP7_75t_L g4107 ( 
.A(n_4059),
.Y(n_4107)
);

OR2x2_ASAP7_75t_L g4108 ( 
.A(n_4071),
.B(n_3924),
.Y(n_4108)
);

NAND2x1p5_ASAP7_75t_L g4109 ( 
.A(n_4058),
.B(n_3678),
.Y(n_4109)
);

OAI211xp5_ASAP7_75t_L g4110 ( 
.A1(n_4056),
.A2(n_4005),
.B(n_3987),
.C(n_3997),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_4078),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_4090),
.B(n_4061),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_4085),
.Y(n_4113)
);

INVx2_ASAP7_75t_SL g4114 ( 
.A(n_4083),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_4085),
.Y(n_4115)
);

OR2x2_ASAP7_75t_L g4116 ( 
.A(n_4074),
.B(n_4042),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_L g4117 ( 
.A(n_4090),
.B(n_4080),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_4105),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_4105),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_4090),
.B(n_4042),
.Y(n_4120)
);

OAI21xp33_ASAP7_75t_L g4121 ( 
.A1(n_4110),
.A2(n_3990),
.B(n_4047),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_4100),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_4100),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_4102),
.Y(n_4124)
);

INVx2_ASAP7_75t_L g4125 ( 
.A(n_4081),
.Y(n_4125)
);

HB1xp67_ASAP7_75t_L g4126 ( 
.A(n_4087),
.Y(n_4126)
);

AOI211xp5_ASAP7_75t_L g4127 ( 
.A1(n_4110),
.A2(n_4009),
.B(n_4018),
.C(n_4014),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_4106),
.Y(n_4128)
);

NAND2x1p5_ASAP7_75t_L g4129 ( 
.A(n_4101),
.B(n_4058),
.Y(n_4129)
);

OR2x2_ASAP7_75t_L g4130 ( 
.A(n_4075),
.B(n_4047),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_4092),
.B(n_4068),
.Y(n_4131)
);

INVx1_ASAP7_75t_SL g4132 ( 
.A(n_4103),
.Y(n_4132)
);

NOR2x1_ASAP7_75t_L g4133 ( 
.A(n_4082),
.B(n_4019),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_4097),
.Y(n_4134)
);

OAI31xp33_ASAP7_75t_L g4135 ( 
.A1(n_4104),
.A2(n_4016),
.A3(n_4027),
.B(n_4030),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_4096),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_L g4137 ( 
.A(n_4127),
.B(n_4079),
.Y(n_4137)
);

AOI22xp5_ASAP7_75t_L g4138 ( 
.A1(n_4127),
.A2(n_4104),
.B1(n_4086),
.B2(n_4084),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_4113),
.Y(n_4139)
);

OR2x2_ASAP7_75t_L g4140 ( 
.A(n_4130),
.B(n_4107),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_4115),
.Y(n_4141)
);

INVx1_ASAP7_75t_SL g4142 ( 
.A(n_4132),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_4135),
.B(n_4088),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_4135),
.B(n_4099),
.Y(n_4144)
);

AND2x4_ASAP7_75t_L g4145 ( 
.A(n_4114),
.B(n_4033),
.Y(n_4145)
);

OAI22xp5_ASAP7_75t_L g4146 ( 
.A1(n_4129),
.A2(n_4077),
.B1(n_4076),
.B2(n_4093),
.Y(n_4146)
);

O2A1O1Ixp33_ASAP7_75t_L g4147 ( 
.A1(n_4121),
.A2(n_4109),
.B(n_4089),
.C(n_4096),
.Y(n_4147)
);

AOI22xp5_ASAP7_75t_L g4148 ( 
.A1(n_4121),
.A2(n_4107),
.B1(n_4052),
.B2(n_4046),
.Y(n_4148)
);

OAI21xp5_ASAP7_75t_L g4149 ( 
.A1(n_4133),
.A2(n_4109),
.B(n_4089),
.Y(n_4149)
);

INVx3_ASAP7_75t_L g4150 ( 
.A(n_4111),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_4118),
.Y(n_4151)
);

AND2x2_ASAP7_75t_L g4152 ( 
.A(n_4116),
.B(n_4094),
.Y(n_4152)
);

OAI221xp5_ASAP7_75t_L g4153 ( 
.A1(n_4120),
.A2(n_4108),
.B1(n_4091),
.B2(n_4098),
.C(n_4081),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_4119),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_4126),
.Y(n_4155)
);

AND2x4_ASAP7_75t_L g4156 ( 
.A(n_4117),
.B(n_4122),
.Y(n_4156)
);

HB1xp67_ASAP7_75t_L g4157 ( 
.A(n_4125),
.Y(n_4157)
);

NOR2x1_ASAP7_75t_L g4158 ( 
.A(n_4142),
.B(n_4123),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_L g4159 ( 
.A(n_4138),
.B(n_4136),
.Y(n_4159)
);

OAI21xp5_ASAP7_75t_L g4160 ( 
.A1(n_4137),
.A2(n_4112),
.B(n_4124),
.Y(n_4160)
);

A2O1A1Ixp33_ASAP7_75t_L g4161 ( 
.A1(n_4145),
.A2(n_4134),
.B(n_4128),
.C(n_4131),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_4143),
.B(n_4095),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_4156),
.B(n_4098),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_4156),
.B(n_4091),
.Y(n_4164)
);

AND2x2_ASAP7_75t_L g4165 ( 
.A(n_4145),
.B(n_4060),
.Y(n_4165)
);

AOI22xp33_ASAP7_75t_L g4166 ( 
.A1(n_4153),
.A2(n_3917),
.B1(n_4059),
.B2(n_3971),
.Y(n_4166)
);

AOI21xp5_ASAP7_75t_SL g4167 ( 
.A1(n_4147),
.A2(n_4144),
.B(n_4141),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_4140),
.Y(n_4168)
);

AOI221xp5_ASAP7_75t_L g4169 ( 
.A1(n_4155),
.A2(n_3926),
.B1(n_3947),
.B2(n_3946),
.C(n_3925),
.Y(n_4169)
);

INVx1_ASAP7_75t_SL g4170 ( 
.A(n_4150),
.Y(n_4170)
);

AND2x4_ASAP7_75t_L g4171 ( 
.A(n_4139),
.B(n_4050),
.Y(n_4171)
);

INVx1_ASAP7_75t_SL g4172 ( 
.A(n_4157),
.Y(n_4172)
);

OAI22xp5_ASAP7_75t_L g4173 ( 
.A1(n_4148),
.A2(n_4050),
.B1(n_4062),
.B2(n_4072),
.Y(n_4173)
);

NAND3xp33_ASAP7_75t_L g4174 ( 
.A(n_4151),
.B(n_3784),
.C(n_3791),
.Y(n_4174)
);

INVx2_ASAP7_75t_L g4175 ( 
.A(n_4152),
.Y(n_4175)
);

AND2x2_ASAP7_75t_L g4176 ( 
.A(n_4146),
.B(n_3950),
.Y(n_4176)
);

AOI211xp5_ASAP7_75t_L g4177 ( 
.A1(n_4154),
.A2(n_3812),
.B(n_3789),
.C(n_3770),
.Y(n_4177)
);

XOR2x2_ASAP7_75t_L g4178 ( 
.A(n_4149),
.B(n_3917),
.Y(n_4178)
);

AND2x4_ASAP7_75t_L g4179 ( 
.A(n_4145),
.B(n_3933),
.Y(n_4179)
);

NAND2x1p5_ASAP7_75t_L g4180 ( 
.A(n_4142),
.B(n_3795),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_4180),
.Y(n_4181)
);

NAND3xp33_ASAP7_75t_L g4182 ( 
.A(n_4158),
.B(n_3820),
.C(n_3790),
.Y(n_4182)
);

AOI21xp5_ASAP7_75t_L g4183 ( 
.A1(n_4164),
.A2(n_3917),
.B(n_3938),
.Y(n_4183)
);

NAND2x1_ASAP7_75t_L g4184 ( 
.A(n_4179),
.B(n_3917),
.Y(n_4184)
);

AND2x4_ASAP7_75t_L g4185 ( 
.A(n_4170),
.B(n_3938),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_L g4186 ( 
.A(n_4172),
.B(n_3921),
.Y(n_4186)
);

AOI21xp5_ASAP7_75t_L g4187 ( 
.A1(n_4167),
.A2(n_3507),
.B(n_3498),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4163),
.Y(n_4188)
);

AOI21xp33_ASAP7_75t_L g4189 ( 
.A1(n_4159),
.A2(n_440),
.B(n_441),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_SL g4190 ( 
.A(n_4179),
.B(n_3915),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_SL g4191 ( 
.A(n_4160),
.B(n_3915),
.Y(n_4191)
);

OR2x2_ASAP7_75t_L g4192 ( 
.A(n_4168),
.B(n_3921),
.Y(n_4192)
);

OR2x2_ASAP7_75t_L g4193 ( 
.A(n_4175),
.B(n_3923),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4171),
.Y(n_4194)
);

AOI222xp33_ASAP7_75t_L g4195 ( 
.A1(n_4162),
.A2(n_3923),
.B1(n_3971),
.B2(n_3970),
.C1(n_3924),
.C2(n_3930),
.Y(n_4195)
);

NAND2xp5_ASAP7_75t_L g4196 ( 
.A(n_4176),
.B(n_3930),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_4171),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_4165),
.B(n_3936),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4174),
.Y(n_4199)
);

AOI21xp33_ASAP7_75t_SL g4200 ( 
.A1(n_4161),
.A2(n_440),
.B(n_441),
.Y(n_4200)
);

INVx2_ASAP7_75t_SL g4201 ( 
.A(n_4178),
.Y(n_4201)
);

OAI21xp33_ASAP7_75t_L g4202 ( 
.A1(n_4166),
.A2(n_3826),
.B(n_3915),
.Y(n_4202)
);

AOI22xp33_ASAP7_75t_SL g4203 ( 
.A1(n_4173),
.A2(n_3973),
.B1(n_3915),
.B2(n_3816),
.Y(n_4203)
);

AND2x2_ASAP7_75t_L g4204 ( 
.A(n_4169),
.B(n_3936),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4177),
.Y(n_4205)
);

NAND4xp25_ASAP7_75t_L g4206 ( 
.A(n_4164),
.B(n_3617),
.C(n_3587),
.D(n_3518),
.Y(n_4206)
);

AOI22xp5_ASAP7_75t_L g4207 ( 
.A1(n_4201),
.A2(n_3915),
.B1(n_3973),
.B2(n_3943),
.Y(n_4207)
);

AOI211xp5_ASAP7_75t_L g4208 ( 
.A1(n_4200),
.A2(n_3973),
.B(n_3649),
.C(n_3657),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_SL g4209 ( 
.A(n_4181),
.B(n_3973),
.Y(n_4209)
);

OAI32xp33_ASAP7_75t_L g4210 ( 
.A1(n_4205),
.A2(n_3942),
.A3(n_3948),
.B1(n_3944),
.B2(n_3943),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_4188),
.Y(n_4211)
);

AOI22xp33_ASAP7_75t_L g4212 ( 
.A1(n_4199),
.A2(n_3973),
.B1(n_3944),
.B2(n_3948),
.Y(n_4212)
);

AOI21xp33_ASAP7_75t_SL g4213 ( 
.A1(n_4189),
.A2(n_442),
.B(n_443),
.Y(n_4213)
);

NOR2xp33_ASAP7_75t_L g4214 ( 
.A(n_4194),
.B(n_442),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_4197),
.Y(n_4215)
);

AOI211xp5_ASAP7_75t_L g4216 ( 
.A1(n_4187),
.A2(n_3753),
.B(n_3646),
.C(n_3520),
.Y(n_4216)
);

O2A1O1Ixp33_ASAP7_75t_L g4217 ( 
.A1(n_4191),
.A2(n_4186),
.B(n_4190),
.C(n_4185),
.Y(n_4217)
);

AOI211xp5_ASAP7_75t_L g4218 ( 
.A1(n_4185),
.A2(n_3526),
.B(n_3533),
.C(n_3633),
.Y(n_4218)
);

AOI211xp5_ASAP7_75t_L g4219 ( 
.A1(n_4182),
.A2(n_3641),
.B(n_3792),
.C(n_3718),
.Y(n_4219)
);

INVx2_ASAP7_75t_SL g4220 ( 
.A(n_4193),
.Y(n_4220)
);

OAI321xp33_ASAP7_75t_L g4221 ( 
.A1(n_4202),
.A2(n_3640),
.A3(n_3816),
.B1(n_3647),
.B2(n_3942),
.C(n_3954),
.Y(n_4221)
);

AOI211xp5_ASAP7_75t_L g4222 ( 
.A1(n_4192),
.A2(n_4206),
.B(n_4183),
.C(n_4204),
.Y(n_4222)
);

OAI322xp33_ASAP7_75t_L g4223 ( 
.A1(n_4184),
.A2(n_3954),
.A3(n_3580),
.B1(n_447),
.B2(n_448),
.C1(n_449),
.C2(n_451),
.Y(n_4223)
);

AOI221xp5_ASAP7_75t_L g4224 ( 
.A1(n_4203),
.A2(n_3564),
.B1(n_3497),
.B2(n_3640),
.C(n_452),
.Y(n_4224)
);

NAND3xp33_ASAP7_75t_SL g4225 ( 
.A(n_4195),
.B(n_445),
.C(n_446),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4198),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_4196),
.B(n_446),
.Y(n_4227)
);

NAND5xp2_ASAP7_75t_L g4228 ( 
.A(n_4205),
.B(n_447),
.C(n_453),
.D(n_454),
.E(n_456),
.Y(n_4228)
);

AOI31xp33_ASAP7_75t_L g4229 ( 
.A1(n_4205),
.A2(n_456),
.A3(n_453),
.B(n_454),
.Y(n_4229)
);

INVx2_ASAP7_75t_L g4230 ( 
.A(n_4181),
.Y(n_4230)
);

AOI22xp5_ASAP7_75t_L g4231 ( 
.A1(n_4201),
.A2(n_3489),
.B1(n_3605),
.B2(n_3553),
.Y(n_4231)
);

OAI22x1_ASAP7_75t_L g4232 ( 
.A1(n_4205),
.A2(n_3580),
.B1(n_3423),
.B2(n_459),
.Y(n_4232)
);

AOI222xp33_ASAP7_75t_L g4233 ( 
.A1(n_4205),
.A2(n_3483),
.B1(n_3552),
.B2(n_3496),
.C1(n_3640),
.C2(n_3475),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_4188),
.Y(n_4234)
);

NOR2xp33_ASAP7_75t_SL g4235 ( 
.A(n_4181),
.B(n_457),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_L g4236 ( 
.A(n_4201),
.B(n_458),
.Y(n_4236)
);

INVxp67_ASAP7_75t_SL g4237 ( 
.A(n_4188),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_L g4238 ( 
.A(n_4230),
.B(n_458),
.Y(n_4238)
);

AOI211xp5_ASAP7_75t_L g4239 ( 
.A1(n_4213),
.A2(n_462),
.B(n_460),
.C(n_461),
.Y(n_4239)
);

AOI22xp5_ASAP7_75t_L g4240 ( 
.A1(n_4235),
.A2(n_3423),
.B1(n_3429),
.B2(n_3453),
.Y(n_4240)
);

AOI22xp5_ASAP7_75t_L g4241 ( 
.A1(n_4214),
.A2(n_3432),
.B1(n_3438),
.B2(n_3436),
.Y(n_4241)
);

AND4x1_ASAP7_75t_L g4242 ( 
.A(n_4236),
.B(n_462),
.C(n_460),
.D(n_461),
.Y(n_4242)
);

OAI211xp5_ASAP7_75t_SL g4243 ( 
.A1(n_4215),
.A2(n_466),
.B(n_464),
.C(n_465),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_L g4244 ( 
.A(n_4237),
.B(n_465),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4229),
.Y(n_4245)
);

OAI21xp5_ASAP7_75t_L g4246 ( 
.A1(n_4225),
.A2(n_3584),
.B(n_3579),
.Y(n_4246)
);

OAI211xp5_ASAP7_75t_SL g4247 ( 
.A1(n_4211),
.A2(n_469),
.B(n_466),
.C(n_468),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_SL g4248 ( 
.A(n_4234),
.B(n_3596),
.Y(n_4248)
);

AOI22xp5_ASAP7_75t_L g4249 ( 
.A1(n_4226),
.A2(n_3426),
.B1(n_3471),
.B2(n_3481),
.Y(n_4249)
);

AOI21xp5_ASAP7_75t_L g4250 ( 
.A1(n_4227),
.A2(n_3610),
.B(n_3598),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_4222),
.B(n_468),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_L g4252 ( 
.A(n_4224),
.B(n_4208),
.Y(n_4252)
);

NOR3xp33_ASAP7_75t_L g4253 ( 
.A(n_4228),
.B(n_469),
.C(n_470),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_4220),
.B(n_470),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4217),
.Y(n_4255)
);

NOR4xp25_ASAP7_75t_L g4256 ( 
.A(n_4209),
.B(n_473),
.C(n_471),
.D(n_472),
.Y(n_4256)
);

OA22x2_ASAP7_75t_L g4257 ( 
.A1(n_4207),
.A2(n_3612),
.B1(n_3624),
.B2(n_3619),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_L g4258 ( 
.A(n_4233),
.B(n_471),
.Y(n_4258)
);

XNOR2x1_ASAP7_75t_SL g4259 ( 
.A(n_4232),
.B(n_4221),
.Y(n_4259)
);

AND2x2_ASAP7_75t_L g4260 ( 
.A(n_4212),
.B(n_475),
.Y(n_4260)
);

NOR2xp33_ASAP7_75t_L g4261 ( 
.A(n_4210),
.B(n_476),
.Y(n_4261)
);

NAND4xp25_ASAP7_75t_L g4262 ( 
.A(n_4231),
.B(n_478),
.C(n_476),
.D(n_477),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_L g4263 ( 
.A(n_4216),
.B(n_4219),
.Y(n_4263)
);

AND4x1_ASAP7_75t_L g4264 ( 
.A(n_4218),
.B(n_482),
.C(n_479),
.D(n_481),
.Y(n_4264)
);

NAND3xp33_ASAP7_75t_L g4265 ( 
.A(n_4255),
.B(n_4223),
.C(n_479),
.Y(n_4265)
);

NAND4xp25_ASAP7_75t_L g4266 ( 
.A(n_4245),
.B(n_4223),
.C(n_484),
.D(n_485),
.Y(n_4266)
);

NAND5xp2_ASAP7_75t_L g4267 ( 
.A(n_4239),
.B(n_483),
.C(n_484),
.D(n_485),
.E(n_486),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_SL g4268 ( 
.A(n_4251),
.B(n_3629),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_SL g4269 ( 
.A(n_4260),
.B(n_486),
.Y(n_4269)
);

NOR3xp33_ASAP7_75t_L g4270 ( 
.A(n_4244),
.B(n_488),
.C(n_489),
.Y(n_4270)
);

NAND4xp25_ASAP7_75t_L g4271 ( 
.A(n_4252),
.B(n_4253),
.C(n_4261),
.D(n_4262),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_4256),
.B(n_488),
.Y(n_4272)
);

AOI21xp5_ASAP7_75t_L g4273 ( 
.A1(n_4238),
.A2(n_491),
.B(n_492),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_4254),
.Y(n_4274)
);

NAND4xp75_ASAP7_75t_L g4275 ( 
.A(n_4258),
.B(n_4263),
.C(n_4248),
.D(n_4259),
.Y(n_4275)
);

NOR3xp33_ASAP7_75t_L g4276 ( 
.A(n_4247),
.B(n_491),
.C(n_492),
.Y(n_4276)
);

NOR3xp33_ASAP7_75t_SL g4277 ( 
.A(n_4243),
.B(n_493),
.C(n_494),
.Y(n_4277)
);

O2A1O1Ixp33_ASAP7_75t_L g4278 ( 
.A1(n_4242),
.A2(n_495),
.B(n_496),
.C(n_497),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_4264),
.B(n_495),
.Y(n_4279)
);

NOR3x1_ASAP7_75t_L g4280 ( 
.A(n_4246),
.B(n_496),
.C(n_498),
.Y(n_4280)
);

NAND3xp33_ASAP7_75t_L g4281 ( 
.A(n_4241),
.B(n_498),
.C(n_499),
.Y(n_4281)
);

NOR2xp33_ASAP7_75t_L g4282 ( 
.A(n_4250),
.B(n_499),
.Y(n_4282)
);

NOR3xp33_ASAP7_75t_L g4283 ( 
.A(n_4240),
.B(n_500),
.C(n_501),
.Y(n_4283)
);

NAND3xp33_ASAP7_75t_L g4284 ( 
.A(n_4249),
.B(n_501),
.C(n_502),
.Y(n_4284)
);

NOR4xp25_ASAP7_75t_L g4285 ( 
.A(n_4257),
.B(n_504),
.C(n_505),
.D(n_507),
.Y(n_4285)
);

OAI211xp5_ASAP7_75t_L g4286 ( 
.A1(n_4255),
.A2(n_505),
.B(n_508),
.C(n_509),
.Y(n_4286)
);

OAI221xp5_ASAP7_75t_L g4287 ( 
.A1(n_4256),
.A2(n_509),
.B1(n_510),
.B2(n_511),
.C(n_512),
.Y(n_4287)
);

NOR2x1_ASAP7_75t_L g4288 ( 
.A(n_4255),
.B(n_510),
.Y(n_4288)
);

NOR5xp2_ASAP7_75t_L g4289 ( 
.A(n_4255),
.B(n_511),
.C(n_513),
.D(n_514),
.E(n_515),
.Y(n_4289)
);

OAI211xp5_ASAP7_75t_L g4290 ( 
.A1(n_4278),
.A2(n_513),
.B(n_516),
.C(n_517),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4279),
.Y(n_4291)
);

AOI21xp5_ASAP7_75t_L g4292 ( 
.A1(n_4272),
.A2(n_516),
.B(n_518),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4288),
.Y(n_4293)
);

NAND4xp75_ASAP7_75t_L g4294 ( 
.A(n_4280),
.B(n_518),
.C(n_519),
.D(n_520),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_4286),
.Y(n_4295)
);

NOR2x1_ASAP7_75t_L g4296 ( 
.A(n_4275),
.B(n_519),
.Y(n_4296)
);

NOR2x1_ASAP7_75t_L g4297 ( 
.A(n_4271),
.B(n_520),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4269),
.Y(n_4298)
);

NAND4xp75_ASAP7_75t_L g4299 ( 
.A(n_4273),
.B(n_521),
.C(n_522),
.D(n_524),
.Y(n_4299)
);

NAND2xp5_ASAP7_75t_L g4300 ( 
.A(n_4285),
.B(n_521),
.Y(n_4300)
);

NOR3xp33_ASAP7_75t_L g4301 ( 
.A(n_4287),
.B(n_522),
.C(n_524),
.Y(n_4301)
);

NOR3xp33_ASAP7_75t_L g4302 ( 
.A(n_4266),
.B(n_4270),
.C(n_4265),
.Y(n_4302)
);

HB1xp67_ASAP7_75t_L g4303 ( 
.A(n_4274),
.Y(n_4303)
);

AND2x4_ASAP7_75t_L g4304 ( 
.A(n_4277),
.B(n_525),
.Y(n_4304)
);

OAI222xp33_ASAP7_75t_L g4305 ( 
.A1(n_4268),
.A2(n_3580),
.B1(n_527),
.B2(n_528),
.C1(n_529),
.C2(n_530),
.Y(n_4305)
);

NAND2xp5_ASAP7_75t_L g4306 ( 
.A(n_4276),
.B(n_526),
.Y(n_4306)
);

OAI22x1_ASAP7_75t_L g4307 ( 
.A1(n_4282),
.A2(n_4281),
.B1(n_4284),
.B2(n_4267),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4283),
.Y(n_4308)
);

INVx2_ASAP7_75t_L g4309 ( 
.A(n_4289),
.Y(n_4309)
);

NOR2x1_ASAP7_75t_L g4310 ( 
.A(n_4288),
.B(n_526),
.Y(n_4310)
);

NOR2x1_ASAP7_75t_L g4311 ( 
.A(n_4288),
.B(n_527),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4279),
.Y(n_4312)
);

AOI22xp5_ASAP7_75t_L g4313 ( 
.A1(n_4276),
.A2(n_3477),
.B1(n_532),
.B2(n_533),
.Y(n_4313)
);

AOI22xp5_ASAP7_75t_L g4314 ( 
.A1(n_4276),
.A2(n_531),
.B1(n_534),
.B2(n_535),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_L g4315 ( 
.A(n_4304),
.B(n_531),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4296),
.Y(n_4316)
);

NOR3xp33_ASAP7_75t_L g4317 ( 
.A(n_4290),
.B(n_535),
.C(n_536),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4304),
.Y(n_4318)
);

INVx2_ASAP7_75t_L g4319 ( 
.A(n_4309),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4294),
.Y(n_4320)
);

AND2x2_ASAP7_75t_L g4321 ( 
.A(n_4295),
.B(n_4301),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4310),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4311),
.Y(n_4323)
);

OAI22xp33_ASAP7_75t_L g4324 ( 
.A1(n_4300),
.A2(n_536),
.B1(n_537),
.B2(n_538),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_4297),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4299),
.Y(n_4326)
);

INVxp67_ASAP7_75t_SL g4327 ( 
.A(n_4306),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4303),
.Y(n_4328)
);

HB1xp67_ASAP7_75t_L g4329 ( 
.A(n_4308),
.Y(n_4329)
);

OR2x2_ASAP7_75t_L g4330 ( 
.A(n_4291),
.B(n_537),
.Y(n_4330)
);

INVx2_ASAP7_75t_L g4331 ( 
.A(n_4298),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4314),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_SL g4333 ( 
.A(n_4302),
.B(n_539),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_4307),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4293),
.Y(n_4335)
);

INVx2_ASAP7_75t_L g4336 ( 
.A(n_4312),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_4292),
.B(n_540),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4315),
.Y(n_4338)
);

OR2x2_ASAP7_75t_L g4339 ( 
.A(n_4315),
.B(n_4313),
.Y(n_4339)
);

HB1xp67_ASAP7_75t_L g4340 ( 
.A(n_4334),
.Y(n_4340)
);

NOR4xp75_ASAP7_75t_SL g4341 ( 
.A(n_4337),
.B(n_4317),
.C(n_4324),
.D(n_4333),
.Y(n_4341)
);

NOR4xp25_ASAP7_75t_L g4342 ( 
.A(n_4328),
.B(n_4305),
.C(n_542),
.D(n_543),
.Y(n_4342)
);

NAND3xp33_ASAP7_75t_L g4343 ( 
.A(n_4318),
.B(n_540),
.C(n_542),
.Y(n_4343)
);

HB1xp67_ASAP7_75t_L g4344 ( 
.A(n_4319),
.Y(n_4344)
);

INVx2_ASAP7_75t_L g4345 ( 
.A(n_4331),
.Y(n_4345)
);

BUFx2_ASAP7_75t_L g4346 ( 
.A(n_4320),
.Y(n_4346)
);

AOI221xp5_ASAP7_75t_SL g4347 ( 
.A1(n_4316),
.A2(n_544),
.B1(n_545),
.B2(n_547),
.C(n_548),
.Y(n_4347)
);

AND2x4_ASAP7_75t_L g4348 ( 
.A(n_4336),
.B(n_544),
.Y(n_4348)
);

HB1xp67_ASAP7_75t_L g4349 ( 
.A(n_4321),
.Y(n_4349)
);

NOR3xp33_ASAP7_75t_L g4350 ( 
.A(n_4337),
.B(n_547),
.C(n_549),
.Y(n_4350)
);

OR5x1_ASAP7_75t_L g4351 ( 
.A(n_4329),
.B(n_550),
.C(n_551),
.D(n_552),
.E(n_553),
.Y(n_4351)
);

OR2x2_ASAP7_75t_L g4352 ( 
.A(n_4330),
.B(n_550),
.Y(n_4352)
);

INVx1_ASAP7_75t_SL g4353 ( 
.A(n_4335),
.Y(n_4353)
);

OR2x2_ASAP7_75t_L g4354 ( 
.A(n_4345),
.B(n_4326),
.Y(n_4354)
);

NOR2xp33_ASAP7_75t_R g4355 ( 
.A(n_4338),
.B(n_4322),
.Y(n_4355)
);

OAI221xp5_ASAP7_75t_L g4356 ( 
.A1(n_4347),
.A2(n_4342),
.B1(n_4340),
.B2(n_4350),
.C(n_4353),
.Y(n_4356)
);

NAND2xp33_ASAP7_75t_SL g4357 ( 
.A(n_4344),
.B(n_4325),
.Y(n_4357)
);

OAI221xp5_ASAP7_75t_L g4358 ( 
.A1(n_4343),
.A2(n_4332),
.B1(n_4327),
.B2(n_4323),
.C(n_557),
.Y(n_4358)
);

CKINVDCx5p33_ASAP7_75t_R g4359 ( 
.A(n_4346),
.Y(n_4359)
);

CKINVDCx16_ASAP7_75t_R g4360 ( 
.A(n_4348),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4348),
.Y(n_4361)
);

CKINVDCx5p33_ASAP7_75t_R g4362 ( 
.A(n_4349),
.Y(n_4362)
);

BUFx2_ASAP7_75t_R g4363 ( 
.A(n_4352),
.Y(n_4363)
);

NOR2xp33_ASAP7_75t_R g4364 ( 
.A(n_4339),
.B(n_553),
.Y(n_4364)
);

CKINVDCx5p33_ASAP7_75t_R g4365 ( 
.A(n_4341),
.Y(n_4365)
);

BUFx2_ASAP7_75t_L g4366 ( 
.A(n_4351),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_L g4367 ( 
.A(n_4345),
.B(n_554),
.Y(n_4367)
);

OAI221xp5_ASAP7_75t_L g4368 ( 
.A1(n_4357),
.A2(n_554),
.B1(n_555),
.B2(n_558),
.C(n_560),
.Y(n_4368)
);

NAND2xp5_ASAP7_75t_L g4369 ( 
.A(n_4362),
.B(n_558),
.Y(n_4369)
);

CKINVDCx5p33_ASAP7_75t_R g4370 ( 
.A(n_4364),
.Y(n_4370)
);

O2A1O1Ixp33_ASAP7_75t_L g4371 ( 
.A1(n_4367),
.A2(n_560),
.B(n_561),
.C(n_562),
.Y(n_4371)
);

BUFx2_ASAP7_75t_L g4372 ( 
.A(n_4359),
.Y(n_4372)
);

AOI22xp33_ASAP7_75t_L g4373 ( 
.A1(n_4366),
.A2(n_563),
.B1(n_564),
.B2(n_565),
.Y(n_4373)
);

AOI22xp33_ASAP7_75t_R g4374 ( 
.A1(n_4355),
.A2(n_563),
.B1(n_564),
.B2(n_566),
.Y(n_4374)
);

AOI221xp5_ASAP7_75t_L g4375 ( 
.A1(n_4356),
.A2(n_566),
.B1(n_568),
.B2(n_569),
.C(n_570),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4354),
.Y(n_4376)
);

NAND4xp25_ASAP7_75t_L g4377 ( 
.A(n_4358),
.B(n_568),
.C(n_569),
.D(n_570),
.Y(n_4377)
);

HB1xp67_ASAP7_75t_SL g4378 ( 
.A(n_4363),
.Y(n_4378)
);

AO22x2_ASAP7_75t_L g4379 ( 
.A1(n_4376),
.A2(n_4361),
.B1(n_4360),
.B2(n_4365),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4378),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_4369),
.Y(n_4381)
);

BUFx2_ASAP7_75t_L g4382 ( 
.A(n_4372),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_4368),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_4371),
.Y(n_4384)
);

OAI21x1_ASAP7_75t_L g4385 ( 
.A1(n_4377),
.A2(n_571),
.B(n_572),
.Y(n_4385)
);

INVx1_ASAP7_75t_SL g4386 ( 
.A(n_4370),
.Y(n_4386)
);

AO22x2_ASAP7_75t_L g4387 ( 
.A1(n_4380),
.A2(n_4374),
.B1(n_4375),
.B2(n_4373),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_L g4388 ( 
.A(n_4379),
.B(n_572),
.Y(n_4388)
);

INVx2_ASAP7_75t_L g4389 ( 
.A(n_4379),
.Y(n_4389)
);

AOI21xp5_ASAP7_75t_L g4390 ( 
.A1(n_4383),
.A2(n_573),
.B(n_575),
.Y(n_4390)
);

CKINVDCx20_ASAP7_75t_R g4391 ( 
.A(n_4382),
.Y(n_4391)
);

OAI22xp5_ASAP7_75t_L g4392 ( 
.A1(n_4384),
.A2(n_573),
.B1(n_575),
.B2(n_576),
.Y(n_4392)
);

AOI21xp5_ASAP7_75t_L g4393 ( 
.A1(n_4386),
.A2(n_576),
.B(n_577),
.Y(n_4393)
);

XNOR2xp5_ASAP7_75t_L g4394 ( 
.A(n_4391),
.B(n_4385),
.Y(n_4394)
);

OR2x2_ASAP7_75t_SL g4395 ( 
.A(n_4389),
.B(n_4381),
.Y(n_4395)
);

OAI22xp5_ASAP7_75t_L g4396 ( 
.A1(n_4394),
.A2(n_4388),
.B1(n_4387),
.B2(n_4390),
.Y(n_4396)
);

HB1xp67_ASAP7_75t_L g4397 ( 
.A(n_4396),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4397),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_4398),
.Y(n_4399)
);

AOI22xp5_ASAP7_75t_L g4400 ( 
.A1(n_4399),
.A2(n_4395),
.B1(n_4393),
.B2(n_4392),
.Y(n_4400)
);

AOI211xp5_ASAP7_75t_L g4401 ( 
.A1(n_4400),
.A2(n_578),
.B(n_580),
.C(n_581),
.Y(n_4401)
);


endmodule