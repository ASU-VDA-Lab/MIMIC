module real_jpeg_24371_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g98 ( 
.A(n_0),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_0),
.Y(n_99)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_0),
.Y(n_117)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_0),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_2),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_2),
.A2(n_35),
.B1(n_56),
.B2(n_57),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_2),
.A2(n_35),
.B1(n_73),
.B2(n_75),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_4),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_14)
);

CKINVDCx12_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_7),
.A2(n_10),
.B1(n_24),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_7),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_7),
.A2(n_30),
.B1(n_32),
.B2(n_130),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_7),
.A2(n_56),
.B1(n_57),
.B2(n_130),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_7),
.A2(n_73),
.B1(n_75),
.B2(n_130),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_8),
.A2(n_30),
.B1(n_32),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_8),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_8),
.A2(n_28),
.B1(n_52),
.B2(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_8),
.A2(n_52),
.B1(n_73),
.B2(n_75),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_13),
.A2(n_23),
.B1(n_24),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_13),
.A2(n_40),
.B1(n_56),
.B2(n_57),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_13),
.A2(n_40),
.B1(n_73),
.B2(n_75),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_13),
.A2(n_30),
.B1(n_32),
.B2(n_40),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_13),
.A2(n_26),
.B(n_36),
.C(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_13),
.B(n_29),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_13),
.A2(n_32),
.B(n_55),
.C(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_13),
.B(n_71),
.C(n_73),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_13),
.B(n_53),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_13),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_13),
.B(n_69),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_324),
.Y(n_16)
);

OAI221xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_41),
.B1(n_45),
.B2(n_321),
.C(n_323),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_18),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_18),
.B(n_322),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_18),
.B(n_41),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_37),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_19),
.A2(n_29),
.B(n_142),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_20),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_21),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_29),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_22)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_24),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_32),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_25),
.A2(n_32),
.B(n_40),
.Y(n_198)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_39),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_29),
.B(n_33),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_29),
.B(n_129),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_30),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_30),
.A2(n_32),
.B1(n_55),
.B2(n_59),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_38),
.B(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_40),
.A2(n_56),
.B(n_59),
.Y(n_221)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_41),
.A2(n_96),
.B1(n_105),
.B2(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B(n_44),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_42),
.A2(n_84),
.B(n_316),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_310),
.B(n_320),
.Y(n_45)
);

OAI211xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_131),
.B(n_147),
.C(n_309),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_106),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_48),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_48),
.B(n_106),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_48),
.B(n_133),
.Y(n_309)
);

FAx1_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_81),
.CI(n_95),
.CON(n_48),
.SN(n_48)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_49),
.A2(n_50),
.B(n_64),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_64),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_53),
.B(n_60),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_53),
.B(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_54),
.B(n_63),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_54),
.B(n_140),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_54),
.A2(n_61),
.B(n_140),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_54)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_57),
.B1(n_70),
.B2(n_71),
.Y(n_79)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_57),
.B(n_238),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_60),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_60),
.B(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_61),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_76),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_65),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_66),
.A2(n_68),
.B(n_92),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_67),
.B(n_78),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_68),
.A2(n_77),
.B(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_69),
.B(n_225),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_75),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_73),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_73),
.B(n_263),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_77),
.B(n_235),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_78),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_93),
.B2(n_94),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_82),
.A2(n_93),
.B1(n_135),
.B2(n_145),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_82),
.B(n_87),
.C(n_90),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_82),
.B(n_135),
.C(n_146),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_83),
.B(n_168),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_84),
.B(n_128),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_88),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_89),
.B(n_191),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_90),
.A2(n_91),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_90),
.B(n_180),
.C(n_182),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_90),
.A2(n_91),
.B1(n_182),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_91),
.B(n_138),
.C(n_141),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_101),
.B(n_105),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_96),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_96),
.A2(n_102),
.B1(n_110),
.B2(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_96),
.B(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_96),
.A2(n_110),
.B1(n_220),
.B2(n_280),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B(n_100),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_97),
.A2(n_161),
.B(n_162),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_97),
.B(n_100),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_97),
.B(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_99),
.B(n_120),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_99),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_102),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_104),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_104),
.B(n_224),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.C(n_112),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_111),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_112),
.B(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_122),
.C(n_126),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_114),
.B(n_121),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_115),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_119),
.A2(n_161),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_119),
.B(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_122),
.A2(n_126),
.B1(n_127),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_124),
.B(n_184),
.Y(n_277)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_SL g147 ( 
.A(n_132),
.B(n_148),
.C(n_149),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_146),
.Y(n_133)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_141),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_139),
.B(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_142),
.Y(n_316)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_172),
.B(n_308),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_169),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_151),
.B(n_169),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_157),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_152),
.B(n_155),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_157),
.B(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_166),
.C(n_167),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_158),
.A2(n_159),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_164),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_163),
.B(n_248),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_165),
.B(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_166),
.A2(n_167),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_166),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_166),
.A2(n_297),
.B1(n_315),
.B2(n_317),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_166),
.B(n_312),
.C(n_317),
.Y(n_322)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_167),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_303),
.B(n_307),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_214),
.B(n_289),
.C(n_302),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_202),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_175),
.B(n_202),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_188),
.B2(n_201),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_186),
.B2(n_187),
.Y(n_177)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_178),
.B(n_187),
.C(n_201),
.Y(n_290)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_181),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_SL g192 ( 
.A(n_185),
.Y(n_192)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_196),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_189)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_190),
.B(n_195),
.C(n_196),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_193),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_199),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.C(n_209),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_203),
.A2(n_204),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_209),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_209),
.Y(n_218)
);

FAx1_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.CI(n_213),
.CON(n_209),
.SN(n_209)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_212),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_288),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_229),
.B(n_287),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_226),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_217),
.B(n_226),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.C(n_222),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_218),
.B(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_219),
.B(n_222),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_220),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_282),
.B(n_286),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_273),
.B(n_281),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_252),
.B(n_272),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_239),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_233),
.B(n_239),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_234),
.A2(n_236),
.B1(n_237),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_246),
.B2(n_251),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_242),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_245),
.C(n_251),
.Y(n_274)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_243),
.Y(n_245)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_246),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_250),
.B(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_260),
.B(n_271),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_254),
.B(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

INVx3_ASAP7_75t_SL g256 ( 
.A(n_257),
.Y(n_256)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_257),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_267),
.B(n_270),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_268),
.B(n_269),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_274),
.B(n_275),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_279),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_278),
.C(n_279),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_283),
.B(n_284),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_290),
.B(n_291),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_301),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_299),
.B2(n_300),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_300),
.C(n_301),
.Y(n_304)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_304),
.B(n_305),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_319),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_319),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_318),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_314),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_315),
.Y(n_317)
);


endmodule