module fake_netlist_1_4574_n_517 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_517);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_517;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g74 ( .A(n_22), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_25), .Y(n_75) );
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_17), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_23), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_64), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_2), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_65), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_39), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_57), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_3), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_47), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_15), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_72), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_4), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_35), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_40), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_55), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_4), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_53), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_43), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_8), .Y(n_94) );
INVxp33_ASAP7_75t_L g95 ( .A(n_33), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_42), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_67), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_73), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_19), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_70), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_29), .Y(n_101) );
HB1xp67_ASAP7_75t_L g102 ( .A(n_26), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_61), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_20), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_44), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_52), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_48), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_83), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_81), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_102), .B(n_83), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g111 ( .A(n_79), .B(n_0), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_81), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_75), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_75), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_77), .Y(n_115) );
AND2x4_ASAP7_75t_L g116 ( .A(n_85), .B(n_0), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g117 ( .A(n_77), .B(n_1), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_91), .B(n_1), .Y(n_118) );
AND2x4_ASAP7_75t_L g119 ( .A(n_85), .B(n_2), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g120 ( .A1(n_101), .A2(n_3), .B1(n_5), .B2(n_6), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_84), .B(n_5), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_80), .Y(n_122) );
NOR2x1_ASAP7_75t_L g123 ( .A(n_93), .B(n_6), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_80), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_94), .B(n_7), .Y(n_125) );
OA21x2_ASAP7_75t_L g126 ( .A1(n_82), .A2(n_36), .B(n_69), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_82), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_88), .Y(n_128) );
INVx6_ASAP7_75t_L g129 ( .A(n_95), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_88), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_116), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_116), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_115), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_116), .B(n_97), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_115), .Y(n_135) );
INVx4_ASAP7_75t_L g136 ( .A(n_116), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_129), .B(n_76), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_129), .B(n_96), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_116), .Y(n_139) );
INVx2_ASAP7_75t_SL g140 ( .A(n_129), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_129), .B(n_87), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_129), .B(n_74), .Y(n_142) );
AND2x6_ASAP7_75t_L g143 ( .A(n_119), .B(n_97), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_119), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_108), .B(n_94), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_119), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_119), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_129), .B(n_78), .Y(n_148) );
AND2x6_ASAP7_75t_L g149 ( .A(n_119), .B(n_98), .Y(n_149) );
AND2x2_ASAP7_75t_SL g150 ( .A(n_121), .B(n_99), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_124), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_115), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_124), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_124), .B(n_99), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_124), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_124), .Y(n_156) );
INVx5_ASAP7_75t_L g157 ( .A(n_134), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_150), .B(n_118), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_145), .B(n_118), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_151), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_153), .Y(n_161) );
BUFx2_ASAP7_75t_L g162 ( .A(n_134), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_155), .Y(n_163) );
INVx1_ASAP7_75t_SL g164 ( .A(n_145), .Y(n_164) );
AO22x1_ASAP7_75t_L g165 ( .A1(n_134), .A2(n_120), .B1(n_123), .B2(n_86), .Y(n_165) );
INVx1_ASAP7_75t_SL g166 ( .A(n_145), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_156), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_131), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_132), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_139), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_134), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_134), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_136), .B(n_121), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_134), .Y(n_174) );
AND3x1_ASAP7_75t_SL g175 ( .A(n_150), .B(n_120), .C(n_128), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_136), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_143), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_143), .B(n_121), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_144), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_135), .Y(n_180) );
OR2x2_ASAP7_75t_L g181 ( .A(n_137), .B(n_118), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_143), .A2(n_130), .B1(n_128), .B2(n_127), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_135), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_136), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_141), .B(n_108), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_143), .B(n_130), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_143), .B(n_127), .Y(n_187) );
HB1xp67_ASAP7_75t_SL g188 ( .A(n_143), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_146), .B(n_110), .Y(n_189) );
INVxp67_ASAP7_75t_SL g190 ( .A(n_147), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_159), .B(n_140), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_160), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_160), .Y(n_193) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_164), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_160), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_176), .Y(n_196) );
INVxp67_ASAP7_75t_SL g197 ( .A(n_188), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_171), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_164), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_163), .Y(n_200) );
OAI22xp5_ASAP7_75t_SL g201 ( .A1(n_175), .A2(n_110), .B1(n_140), .B2(n_138), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_171), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_189), .A2(n_111), .B(n_125), .C(n_154), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_166), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_163), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_159), .B(n_138), .Y(n_206) );
INVxp67_ASAP7_75t_L g207 ( .A(n_159), .Y(n_207) );
AOI221xp5_ASAP7_75t_L g208 ( .A1(n_158), .A2(n_113), .B1(n_114), .B2(n_122), .C(n_125), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_167), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_175), .A2(n_149), .B1(n_154), .B2(n_113), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_159), .B(n_149), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_158), .B(n_142), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_166), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_188), .A2(n_148), .B1(n_122), .B2(n_114), .Y(n_214) );
INVx5_ASAP7_75t_L g215 ( .A(n_157), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_171), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_158), .B(n_149), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_185), .A2(n_109), .B(n_112), .C(n_123), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_172), .B(n_149), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_161), .Y(n_220) );
BUFx12f_ASAP7_75t_L g221 ( .A(n_159), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_181), .A2(n_117), .B(n_109), .C(n_112), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_176), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_215), .Y(n_224) );
OAI22xp33_ASAP7_75t_L g225 ( .A1(n_199), .A2(n_182), .B1(n_181), .B2(n_178), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_200), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_217), .B(n_172), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_199), .A2(n_182), .B1(n_190), .B2(n_178), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_201), .A2(n_185), .B1(n_149), .B2(n_173), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_192), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_200), .Y(n_231) );
OAI21x1_ASAP7_75t_L g232 ( .A1(n_205), .A2(n_126), .B(n_180), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_192), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_208), .B(n_181), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_215), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_201), .A2(n_165), .B1(n_149), .B2(n_190), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_204), .A2(n_165), .B1(n_168), .B2(n_169), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_215), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_204), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_221), .A2(n_179), .B1(n_168), .B2(n_169), .Y(n_240) );
CKINVDCx9p33_ASAP7_75t_R g241 ( .A(n_213), .Y(n_241) );
NOR2xp33_ASAP7_75t_SL g242 ( .A(n_221), .B(n_172), .Y(n_242) );
AO21x1_ASAP7_75t_L g243 ( .A1(n_205), .A2(n_209), .B(n_192), .Y(n_243) );
AOI221xp5_ASAP7_75t_L g244 ( .A1(n_207), .A2(n_179), .B1(n_170), .B2(n_167), .C(n_187), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_220), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_217), .B(n_219), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_212), .B(n_186), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_213), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_234), .A2(n_191), .B1(n_212), .B2(n_194), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_226), .Y(n_250) );
AOI22xp33_ASAP7_75t_SL g251 ( .A1(n_239), .A2(n_209), .B1(n_214), .B2(n_220), .Y(n_251) );
AOI21xp33_ASAP7_75t_L g252 ( .A1(n_225), .A2(n_222), .B(n_210), .Y(n_252) );
OAI21xp33_ASAP7_75t_L g253 ( .A1(n_236), .A2(n_218), .B(n_210), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_228), .A2(n_220), .B1(n_193), .B2(n_195), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_239), .A2(n_193), .B1(n_195), .B2(n_211), .Y(n_255) );
OAI211xp5_ASAP7_75t_SL g256 ( .A1(n_229), .A2(n_203), .B(n_89), .C(n_90), .Y(n_256) );
AOI22xp33_ASAP7_75t_SL g257 ( .A1(n_248), .A2(n_174), .B1(n_177), .B2(n_219), .Y(n_257) );
OAI22xp33_ASAP7_75t_L g258 ( .A1(n_248), .A2(n_206), .B1(n_177), .B2(n_174), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_230), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_240), .A2(n_170), .B1(n_196), .B2(n_223), .Y(n_260) );
AND2x2_ASAP7_75t_SL g261 ( .A(n_242), .B(n_162), .Y(n_261) );
OAI211xp5_ASAP7_75t_L g262 ( .A1(n_237), .A2(n_109), .B(n_112), .C(n_107), .Y(n_262) );
AOI22xp33_ASAP7_75t_SL g263 ( .A1(n_241), .A2(n_174), .B1(n_177), .B2(n_219), .Y(n_263) );
OAI33xp33_ASAP7_75t_L g264 ( .A1(n_226), .A2(n_231), .A3(n_96), .B1(n_106), .B2(n_105), .B3(n_104), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_230), .A2(n_186), .B(n_187), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_244), .A2(n_223), .B1(n_196), .B2(n_219), .Y(n_266) );
OAI221xp5_ASAP7_75t_L g267 ( .A1(n_247), .A2(n_231), .B1(n_223), .B2(n_196), .C(n_233), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_233), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_245), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_250), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_259), .Y(n_271) );
OAI33xp33_ASAP7_75t_L g272 ( .A1(n_255), .A2(n_104), .A3(n_90), .B1(n_92), .B2(n_98), .B3(n_106), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_254), .A2(n_243), .B(n_232), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_254), .A2(n_245), .B1(n_247), .B2(n_227), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_252), .A2(n_232), .B(n_197), .Y(n_275) );
AOI222xp33_ASAP7_75t_L g276 ( .A1(n_249), .A2(n_246), .B1(n_89), .B2(n_105), .C1(n_92), .C2(n_103), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_259), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_269), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_268), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_267), .A2(n_227), .B1(n_162), .B2(n_246), .Y(n_280) );
AOI31xp33_ASAP7_75t_L g281 ( .A1(n_251), .A2(n_243), .A3(n_238), .B(n_235), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_250), .B(n_224), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_268), .B(n_246), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_261), .A2(n_266), .B1(n_260), .B2(n_263), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_269), .Y(n_285) );
AO21x2_ASAP7_75t_L g286 ( .A1(n_253), .A2(n_103), .B(n_133), .Y(n_286) );
OAI211xp5_ASAP7_75t_SL g287 ( .A1(n_253), .A2(n_262), .B(n_257), .C(n_258), .Y(n_287) );
INVxp67_ASAP7_75t_L g288 ( .A(n_264), .Y(n_288) );
OAI22xp33_ASAP7_75t_L g289 ( .A1(n_261), .A2(n_238), .B1(n_235), .B2(n_224), .Y(n_289) );
OAI31xp33_ASAP7_75t_L g290 ( .A1(n_256), .A2(n_227), .A3(n_223), .B(n_196), .Y(n_290) );
AOI22xp33_ASAP7_75t_SL g291 ( .A1(n_261), .A2(n_224), .B1(n_126), .B2(n_115), .Y(n_291) );
INVx4_ASAP7_75t_L g292 ( .A(n_282), .Y(n_292) );
INVxp67_ASAP7_75t_SL g293 ( .A(n_279), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_271), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_270), .B(n_126), .Y(n_295) );
NAND4xp25_ASAP7_75t_L g296 ( .A(n_276), .B(n_265), .C(n_8), .D(n_9), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_271), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_271), .Y(n_298) );
XNOR2xp5_ASAP7_75t_L g299 ( .A(n_284), .B(n_7), .Y(n_299) );
NOR2x1_ASAP7_75t_R g300 ( .A(n_282), .B(n_224), .Y(n_300) );
OAI21xp5_ASAP7_75t_L g301 ( .A1(n_288), .A2(n_126), .B(n_161), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_277), .B(n_126), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_270), .B(n_115), .Y(n_303) );
OAI31xp33_ASAP7_75t_L g304 ( .A1(n_280), .A2(n_161), .A3(n_176), .B(n_184), .Y(n_304) );
AOI21xp33_ASAP7_75t_SL g305 ( .A1(n_281), .A2(n_9), .B(n_10), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_277), .B(n_115), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_285), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_285), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_277), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_276), .A2(n_224), .B1(n_115), .B2(n_216), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_287), .A2(n_216), .B1(n_202), .B2(n_198), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_278), .B(n_10), .Y(n_312) );
NAND3xp33_ASAP7_75t_L g313 ( .A(n_281), .B(n_291), .C(n_290), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_283), .B(n_11), .Y(n_314) );
NAND3xp33_ASAP7_75t_SL g315 ( .A(n_290), .B(n_100), .C(n_12), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_280), .A2(n_216), .B1(n_202), .B2(n_198), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_278), .B(n_11), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_278), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_273), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_282), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_273), .Y(n_321) );
OAI31xp33_ASAP7_75t_L g322 ( .A1(n_274), .A2(n_176), .A3(n_184), .B(n_14), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_282), .B(n_12), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_293), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_320), .Y(n_325) );
NOR3xp33_ASAP7_75t_SL g326 ( .A(n_299), .B(n_272), .C(n_289), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_309), .B(n_283), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_299), .A2(n_275), .B1(n_135), .B2(n_152), .C(n_133), .Y(n_328) );
NAND3xp33_ASAP7_75t_L g329 ( .A(n_305), .B(n_275), .C(n_135), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_293), .B(n_286), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_309), .B(n_286), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_294), .B(n_286), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_292), .B(n_286), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_317), .B(n_13), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_307), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_317), .B(n_13), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_307), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_294), .B(n_14), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_308), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_294), .B(n_15), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_308), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_318), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_317), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_318), .B(n_16), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_297), .B(n_16), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_297), .B(n_17), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_297), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_323), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_298), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_323), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_298), .B(n_18), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_323), .B(n_18), .Y(n_352) );
OAI33xp33_ASAP7_75t_L g353 ( .A1(n_296), .A2(n_152), .A3(n_24), .B1(n_27), .B2(n_28), .B3(n_30), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_298), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_320), .B(n_21), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_300), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_312), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_306), .Y(n_358) );
BUFx3_ASAP7_75t_L g359 ( .A(n_320), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_292), .B(n_135), .Y(n_360) );
NAND3xp33_ASAP7_75t_L g361 ( .A(n_305), .B(n_216), .C(n_202), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_292), .B(n_31), .Y(n_362) );
AOI31xp33_ASAP7_75t_L g363 ( .A1(n_300), .A2(n_32), .A3(n_34), .B(n_37), .Y(n_363) );
AOI21xp33_ASAP7_75t_SL g364 ( .A1(n_313), .A2(n_38), .B(n_41), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_296), .B(n_45), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_314), .B(n_46), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_292), .B(n_49), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_303), .B(n_50), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_303), .Y(n_369) );
OAI21x1_ASAP7_75t_SL g370 ( .A1(n_324), .A2(n_310), .B(n_316), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_352), .B(n_315), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_327), .B(n_322), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_327), .B(n_322), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_348), .B(n_321), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_335), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_335), .B(n_306), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_337), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_353), .A2(n_313), .B(n_315), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_337), .B(n_306), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_347), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_339), .B(n_295), .Y(n_381) );
NAND4xp25_ASAP7_75t_L g382 ( .A(n_365), .B(n_304), .C(n_310), .D(n_311), .Y(n_382) );
NOR2x1p5_ASAP7_75t_L g383 ( .A(n_329), .B(n_321), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_350), .B(n_321), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_347), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g386 ( .A(n_367), .B(n_295), .Y(n_386) );
INVx1_ASAP7_75t_SL g387 ( .A(n_325), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_341), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_341), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_358), .B(n_319), .Y(n_390) );
NAND2xp5_ASAP7_75t_R g391 ( .A(n_362), .B(n_302), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_358), .B(n_319), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_343), .B(n_319), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_349), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_342), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_325), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_357), .B(n_302), .Y(n_397) );
INVx1_ASAP7_75t_SL g398 ( .A(n_359), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_342), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_354), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_354), .B(n_302), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_369), .B(n_301), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_344), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_344), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_345), .Y(n_405) );
INVx3_ASAP7_75t_L g406 ( .A(n_333), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_338), .B(n_51), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_359), .B(n_54), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_331), .B(n_332), .Y(n_409) );
NAND4xp25_ASAP7_75t_L g410 ( .A(n_328), .B(n_176), .C(n_184), .D(n_183), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_345), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_338), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_331), .B(n_56), .Y(n_413) );
NAND2xp33_ASAP7_75t_SL g414 ( .A(n_367), .B(n_216), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_340), .B(n_58), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_340), .B(n_59), .Y(n_416) );
INVx2_ASAP7_75t_SL g417 ( .A(n_360), .Y(n_417) );
O2A1O1Ixp33_ASAP7_75t_L g418 ( .A1(n_378), .A2(n_363), .B(n_326), .C(n_364), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_375), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_409), .B(n_351), .Y(n_420) );
NOR2x1p5_ASAP7_75t_L g421 ( .A(n_406), .B(n_361), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_409), .B(n_333), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_377), .Y(n_423) );
INVxp67_ASAP7_75t_L g424 ( .A(n_400), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_403), .B(n_404), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_387), .Y(n_426) );
AND2x2_ASAP7_75t_SL g427 ( .A(n_391), .B(n_362), .Y(n_427) );
NOR3xp33_ASAP7_75t_SL g428 ( .A(n_371), .B(n_334), .C(n_336), .Y(n_428) );
XNOR2xp5_ASAP7_75t_L g429 ( .A(n_396), .B(n_356), .Y(n_429) );
NAND3xp33_ASAP7_75t_L g430 ( .A(n_371), .B(n_330), .C(n_351), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_388), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_380), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_414), .A2(n_355), .B(n_346), .C(n_333), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_389), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_398), .B(n_332), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_405), .B(n_346), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_380), .Y(n_437) );
INVx2_ASAP7_75t_SL g438 ( .A(n_417), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_395), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_399), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_406), .B(n_355), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_417), .B(n_360), .Y(n_442) );
XOR2x2_ASAP7_75t_L g443 ( .A(n_386), .B(n_366), .Y(n_443) );
NOR2x1_ASAP7_75t_L g444 ( .A(n_383), .B(n_368), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_400), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_394), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_394), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_385), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_376), .Y(n_449) );
INVxp67_ASAP7_75t_SL g450 ( .A(n_385), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_379), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_411), .B(n_60), .Y(n_452) );
XOR2x2_ASAP7_75t_L g453 ( .A(n_386), .B(n_62), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_372), .B(n_63), .Y(n_454) );
XOR2xp5_ASAP7_75t_L g455 ( .A(n_373), .B(n_66), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_382), .B(n_68), .Y(n_456) );
INVx1_ASAP7_75t_SL g457 ( .A(n_408), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_406), .B(n_71), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_412), .A2(n_198), .B1(n_202), .B2(n_184), .Y(n_459) );
OAI211xp5_ASAP7_75t_L g460 ( .A1(n_410), .A2(n_215), .B(n_157), .C(n_198), .Y(n_460) );
AOI221x1_ASAP7_75t_L g461 ( .A1(n_370), .A2(n_180), .B1(n_183), .B2(n_184), .C(n_215), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_374), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_392), .Y(n_463) );
AOI31xp33_ASAP7_75t_SL g464 ( .A1(n_415), .A2(n_157), .A3(n_215), .B(n_397), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_401), .B(n_157), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_374), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_384), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_384), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_413), .Y(n_469) );
INVxp33_ASAP7_75t_L g470 ( .A(n_413), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_393), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_381), .Y(n_472) );
XNOR2xp5_ASAP7_75t_L g473 ( .A(n_401), .B(n_157), .Y(n_473) );
OAI21xp5_ASAP7_75t_SL g474 ( .A1(n_407), .A2(n_157), .B(n_416), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_402), .A2(n_371), .B1(n_299), .B2(n_372), .Y(n_475) );
AOI311xp33_ASAP7_75t_L g476 ( .A1(n_390), .A2(n_371), .A3(n_120), .B(n_378), .C(n_94), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_390), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_409), .B(n_403), .Y(n_478) );
XNOR2x1_ASAP7_75t_L g479 ( .A(n_386), .B(n_299), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_375), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_472), .B(n_451), .Y(n_481) );
INVxp33_ASAP7_75t_L g482 ( .A(n_453), .Y(n_482) );
AOI211xp5_ASAP7_75t_L g483 ( .A1(n_418), .A2(n_464), .B(n_456), .C(n_429), .Y(n_483) );
AOI221xp5_ASAP7_75t_SL g484 ( .A1(n_456), .A2(n_425), .B1(n_478), .B2(n_469), .C(n_424), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_445), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_479), .A2(n_475), .B1(n_427), .B2(n_453), .Y(n_486) );
AOI22x1_ASAP7_75t_L g487 ( .A1(n_455), .A2(n_421), .B1(n_426), .B2(n_438), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_427), .A2(n_479), .B1(n_470), .B2(n_433), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g489 ( .A1(n_428), .A2(n_449), .B1(n_424), .B2(n_430), .C(n_471), .Y(n_489) );
INVxp67_ASAP7_75t_SL g490 ( .A(n_450), .Y(n_490) );
OAI32xp33_ASAP7_75t_L g491 ( .A1(n_470), .A2(n_457), .A3(n_420), .B1(n_442), .B2(n_466), .Y(n_491) );
OAI21xp33_ASAP7_75t_SL g492 ( .A1(n_444), .A2(n_450), .B(n_422), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_419), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_433), .A2(n_428), .B1(n_462), .B2(n_468), .Y(n_494) );
OAI221xp5_ASAP7_75t_SL g495 ( .A1(n_474), .A2(n_460), .B1(n_454), .B2(n_436), .C(n_473), .Y(n_495) );
OAI221xp5_ASAP7_75t_L g496 ( .A1(n_476), .A2(n_443), .B1(n_454), .B2(n_434), .C(n_480), .Y(n_496) );
OAI211xp5_ASAP7_75t_L g497 ( .A1(n_486), .A2(n_461), .B(n_458), .C(n_452), .Y(n_497) );
OAI211xp5_ASAP7_75t_L g498 ( .A1(n_487), .A2(n_458), .B(n_459), .C(n_465), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_488), .A2(n_441), .B1(n_465), .B2(n_435), .Y(n_499) );
AOI221xp5_ASAP7_75t_L g500 ( .A1(n_489), .A2(n_447), .B1(n_446), .B2(n_439), .C(n_440), .Y(n_500) );
XNOR2xp5_ASAP7_75t_L g501 ( .A(n_482), .B(n_473), .Y(n_501) );
OA22x2_ASAP7_75t_L g502 ( .A1(n_494), .A2(n_477), .B1(n_467), .B2(n_463), .Y(n_502) );
AO22x1_ASAP7_75t_L g503 ( .A1(n_490), .A2(n_463), .B1(n_423), .B2(n_431), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_484), .A2(n_432), .B1(n_437), .B2(n_448), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_504), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_503), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_502), .Y(n_507) );
NAND3xp33_ASAP7_75t_SL g508 ( .A(n_498), .B(n_483), .C(n_496), .Y(n_508) );
NOR3x1_ASAP7_75t_L g509 ( .A(n_508), .B(n_497), .C(n_501), .Y(n_509) );
NOR3xp33_ASAP7_75t_L g510 ( .A(n_508), .B(n_500), .C(n_492), .Y(n_510) );
AOI22x1_ASAP7_75t_L g511 ( .A1(n_507), .A2(n_485), .B1(n_499), .B2(n_493), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_511), .Y(n_512) );
XNOR2xp5_ASAP7_75t_L g513 ( .A(n_510), .B(n_505), .Y(n_513) );
OR3x1_ASAP7_75t_L g514 ( .A(n_512), .B(n_509), .C(n_506), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_514), .Y(n_515) );
AOI22x1_ASAP7_75t_L g516 ( .A1(n_515), .A2(n_513), .B1(n_491), .B2(n_495), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_516), .A2(n_513), .B(n_481), .Y(n_517) );
endmodule