module real_jpeg_9879_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_343, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_342, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_343;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_342;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_0),
.A2(n_23),
.B1(n_32),
.B2(n_33),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_0),
.A2(n_23),
.B1(n_71),
.B2(n_73),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_0),
.A2(n_23),
.B1(n_53),
.B2(n_54),
.Y(n_269)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_3),
.A2(n_71),
.B1(n_73),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_3),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_3),
.A2(n_53),
.B1(n_54),
.B2(n_112),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_112),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_112),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_4),
.A2(n_71),
.B1(n_73),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_4),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_160),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_160),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_160),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_5),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_5),
.B(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_5),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_5),
.A2(n_133),
.B(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_5),
.A2(n_123),
.B1(n_159),
.B2(n_175),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

BUFx6f_ASAP7_75t_SL g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_10),
.A2(n_35),
.B1(n_53),
.B2(n_54),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_10),
.A2(n_35),
.B1(n_71),
.B2(n_73),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_11),
.A2(n_53),
.B1(n_54),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_11),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_11),
.A2(n_71),
.B1(n_73),
.B2(n_107),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_107),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_107),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_12),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_12),
.A2(n_71),
.B1(n_73),
.B2(n_95),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_95),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_95),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_13),
.A2(n_61),
.B1(n_71),
.B2(n_73),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_13),
.A2(n_53),
.B1(n_54),
.B2(n_61),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_61),
.Y(n_262)
);

A2O1A1O1Ixp25_ASAP7_75t_L g91 ( 
.A1(n_14),
.A2(n_54),
.B(n_66),
.C(n_92),
.D(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_14),
.B(n_54),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_14),
.B(n_52),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_14),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_14),
.A2(n_113),
.B(n_115),
.Y(n_135)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_14),
.A2(n_32),
.B(n_48),
.C(n_149),
.D(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_14),
.B(n_32),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_14),
.B(n_36),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g189 ( 
.A1(n_14),
.A2(n_29),
.B(n_33),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_130),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_16),
.A2(n_24),
.B1(n_25),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_16),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_16),
.A2(n_63),
.B1(n_71),
.B2(n_73),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_16),
.A2(n_53),
.B1(n_54),
.B2(n_63),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_63),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_40),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_38),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_21),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_21),
.B(n_42),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B1(n_34),
.B2(n_36),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_22),
.A2(n_26),
.B1(n_36),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_28),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_24),
.A2(n_28),
.B(n_130),
.C(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_34),
.B(n_36),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_26),
.A2(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_26),
.B(n_209),
.Y(n_218)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_27),
.A2(n_31),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_27),
.A2(n_31),
.B1(n_217),
.B2(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_27),
.A2(n_208),
.B(n_246),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_27),
.A2(n_31),
.B1(n_60),
.B2(n_290),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_31),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_31),
.A2(n_218),
.B(n_290),
.Y(n_289)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_49),
.B(n_51),
.C(n_52),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_49),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_36),
.B(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_81),
.B(n_340),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_76),
.C(n_78),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_43),
.A2(n_44),
.B1(n_335),
.B2(n_337),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_58),
.C(n_64),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_45),
.A2(n_46),
.B1(n_64),
.B2(n_315),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_47),
.A2(n_56),
.B1(n_169),
.B2(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_47),
.A2(n_203),
.B(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_47),
.A2(n_55),
.B1(n_56),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_52),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_48),
.B(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_48),
.A2(n_52),
.B1(n_243),
.B2(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_48),
.A2(n_52),
.B1(n_262),
.B2(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_50),
.B(n_53),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_51),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_52),
.Y(n_56)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_67),
.B(n_69),
.C(n_70),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_67),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_54),
.A2(n_149),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_56),
.B(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_56),
.A2(n_169),
.B(n_170),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_56),
.A2(n_170),
.B(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_58),
.A2(n_59),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_62),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_64),
.A2(n_313),
.B1(n_315),
.B2(n_316),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_64),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_74),
.B(n_75),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_65),
.A2(n_74),
.B1(n_106),
.B2(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_65),
.A2(n_147),
.B(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_65),
.A2(n_74),
.B1(n_200),
.B2(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_65),
.A2(n_74),
.B1(n_228),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_65),
.A2(n_74),
.B1(n_237),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_66),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_66),
.A2(n_70),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_73),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_67),
.B(n_73),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_71),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_70),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_71),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_114),
.Y(n_113)
);

BUFx24_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_73),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_106),
.B(n_108),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_74),
.B(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_74),
.A2(n_108),
.B(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_75),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_76),
.A2(n_78),
.B1(n_79),
.B2(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_76),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_333),
.B(n_339),
.Y(n_81)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_306),
.A3(n_326),
.B1(n_331),
.B2(n_332),
.C(n_342),
.Y(n_82)
);

AOI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_254),
.A3(n_294),
.B1(n_300),
.B2(n_305),
.C(n_343),
.Y(n_83)
);

NOR3xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_211),
.C(n_250),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_182),
.B(n_210),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_163),
.B(n_181),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_141),
.B(n_162),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_118),
.B(n_140),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_100),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_90),
.B(n_100),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_91),
.A2(n_96),
.B1(n_97),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_91),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_93),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_110),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_105),
.C(n_110),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_113),
.B(n_115),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_117),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_113),
.A2(n_114),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_113),
.A2(n_114),
.B1(n_193),
.B2(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_113),
.A2(n_114),
.B1(n_226),
.B2(n_235),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_113),
.A2(n_114),
.B(n_235),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_122),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_130),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_127),
.B(n_139),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_125),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_120),
.B(n_125),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_134),
.B(n_138),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_129),
.B(n_131),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_143),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_154),
.B2(n_161),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_148),
.B1(n_152),
.B2(n_153),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_146),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_148),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_153),
.C(n_161),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_150),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_151),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_158),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_164),
.B(n_165),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_177),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_178),
.C(n_179),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_172),
.B2(n_176),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_173),
.C(n_174),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_172),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_175),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_183),
.B(n_184),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_197),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_186),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_186),
.B(n_196),
.C(n_197),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_191),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_194),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_205),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_201),
.B1(n_202),
.B2(n_204),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_199),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_204),
.C(n_205),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g301 ( 
.A1(n_212),
.A2(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_230),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_213),
.B(n_230),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_224),
.C(n_229),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_223),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_219),
.B1(n_220),
.B2(n_222),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_216),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_222),
.C(n_223),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_229),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_227),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_248),
.B2(n_249),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_233),
.B(n_238),
.C(n_249),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_236),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_244),
.C(n_247),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_241),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_248),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_251),
.B(n_252),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_272),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_255),
.B(n_272),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_265),
.C(n_271),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_256),
.A2(n_257),
.B1(n_265),
.B2(n_299),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_261),
.C(n_263),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_265),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_270),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_267),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_266),
.A2(n_285),
.B(n_289),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_268),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_268),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_269),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_292),
.B2(n_293),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_283),
.B2(n_284),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_275),
.B(n_284),
.C(n_293),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_280),
.B(n_282),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_280),
.Y(n_282)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_281),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_282),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_282),
.A2(n_308),
.B1(n_317),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_291),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_287),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_292),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_295),
.A2(n_301),
.B(n_304),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_296),
.B(n_297),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_319),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_319),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_317),
.C(n_318),
.Y(n_307)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_309),
.A2(n_310),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_315),
.C(n_316),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_321),
.C(n_325),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_313),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_329),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_325),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_327),
.B(n_328),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_338),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_338),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_335),
.Y(n_337)
);


endmodule