module fake_ibex_395_n_1015 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1015);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1015;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_328;
wire n_372;
wire n_293;
wire n_341;
wire n_418;
wire n_256;
wire n_193;
wire n_510;
wire n_845;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_412;
wire n_357;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_317;
wire n_375;
wire n_340;
wire n_280;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_400;
wire n_306;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_980;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_560;
wire n_429;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_1004;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_837;
wire n_797;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_894;
wire n_803;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_951;
wire n_272;
wire n_881;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_320;
wire n_285;
wire n_247;
wire n_379;
wire n_288;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_440;
wire n_268;
wire n_858;
wire n_385;
wire n_342;
wire n_233;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_866;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_1005;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_921;
wire n_912;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_947;
wire n_559;
wire n_425;

BUFx3_ASAP7_75t_L g184 ( 
.A(n_18),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_92),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_53),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_50),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_86),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_93),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_53),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_29),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_79),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_75),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_91),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_98),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_16),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_89),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_21),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_23),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_105),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_22),
.Y(n_204)
);

BUFx2_ASAP7_75t_SL g205 ( 
.A(n_168),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_4),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_100),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_116),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_81),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_10),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_146),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_66),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_125),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_162),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_131),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_121),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_26),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_80),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_133),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_95),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_65),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_2),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_102),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_51),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_77),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_129),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_157),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_36),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_83),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_85),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_36),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_114),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_25),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_44),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_111),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_33),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_19),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_45),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_120),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_97),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_182),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_171),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_1),
.Y(n_245)
);

NOR2xp67_ASAP7_75t_L g246 ( 
.A(n_154),
.B(n_12),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_135),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_172),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_90),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_117),
.Y(n_250)
);

NOR2xp67_ASAP7_75t_L g251 ( 
.A(n_27),
.B(n_158),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_124),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_143),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_21),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_128),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_138),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_150),
.B(n_166),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_180),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_60),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_159),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_107),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_96),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_113),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_38),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_7),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_29),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_144),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_165),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_109),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_82),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_141),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_153),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_38),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_156),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_15),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_48),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_58),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_183),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_22),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_58),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_134),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_20),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_32),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_47),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_177),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_142),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_39),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_88),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_71),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_118),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_72),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_110),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_155),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_136),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_149),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_119),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_51),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_147),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_1),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_6),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_68),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_18),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_163),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_181),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_76),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_164),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_123),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_130),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_7),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_145),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_62),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_104),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_132),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_126),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_37),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_178),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_152),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_17),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_26),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_54),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_35),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_30),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_55),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_69),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_151),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_137),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_108),
.B(n_115),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_70),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_78),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_189),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_245),
.Y(n_331)
);

AND2x2_ASAP7_75t_SL g332 ( 
.A(n_196),
.B(n_59),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_189),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_217),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_271),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_295),
.Y(n_336)
);

INVx5_ASAP7_75t_L g337 ( 
.A(n_222),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_217),
.Y(n_338)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_222),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_232),
.Y(n_340)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_222),
.Y(n_341)
);

OAI22x1_ASAP7_75t_L g342 ( 
.A1(n_200),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_342)
);

BUFx12f_ASAP7_75t_L g343 ( 
.A(n_269),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_329),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_289),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_289),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_184),
.Y(n_347)
);

CKINVDCx11_ASAP7_75t_R g348 ( 
.A(n_206),
.Y(n_348)
);

NOR2x1_ASAP7_75t_L g349 ( 
.A(n_184),
.B(n_61),
.Y(n_349)
);

INVx6_ASAP7_75t_L g350 ( 
.A(n_222),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_198),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_249),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_290),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_249),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_225),
.Y(n_355)
);

AND2x4_ASAP7_75t_L g356 ( 
.A(n_225),
.B(n_5),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_247),
.B(n_8),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

OAI22x1_ASAP7_75t_SL g359 ( 
.A1(n_206),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_359)
);

INVx5_ASAP7_75t_L g360 ( 
.A(n_249),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_279),
.Y(n_361)
);

OAI21x1_ASAP7_75t_L g362 ( 
.A1(n_304),
.A2(n_94),
.B(n_179),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_275),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_363)
);

BUFx8_ASAP7_75t_L g364 ( 
.A(n_279),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_304),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_305),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_283),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_201),
.A2(n_218),
.B1(n_223),
.B2(n_204),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_236),
.Y(n_369)
);

BUFx8_ASAP7_75t_SL g370 ( 
.A(n_233),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_239),
.B(n_11),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_186),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_211),
.B(n_13),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_188),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_305),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_249),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_272),
.Y(n_377)
);

OA21x2_ASAP7_75t_L g378 ( 
.A1(n_187),
.A2(n_99),
.B(n_176),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_264),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_272),
.Y(n_380)
);

OAI22x1_ASAP7_75t_SL g381 ( 
.A1(n_233),
.A2(n_254),
.B1(n_265),
.B2(n_240),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_220),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_273),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_276),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_277),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_385)
);

OA21x2_ASAP7_75t_L g386 ( 
.A1(n_193),
.A2(n_101),
.B(n_175),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_272),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_220),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_264),
.Y(n_389)
);

CKINVDCx11_ASAP7_75t_R g390 ( 
.A(n_240),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_191),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_255),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_190),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_190),
.A2(n_14),
.B1(n_19),
.B2(n_20),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_255),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_282),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_299),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_194),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_302),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_309),
.B(n_23),
.Y(n_400)
);

CKINVDCx11_ASAP7_75t_R g401 ( 
.A(n_254),
.Y(n_401)
);

OAI21x1_ASAP7_75t_L g402 ( 
.A1(n_195),
.A2(n_103),
.B(n_174),
.Y(n_402)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_185),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_199),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_202),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_203),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_319),
.B(n_24),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_321),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_214),
.B(n_231),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_192),
.B(n_28),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_264),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_210),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_297),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_234),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_269),
.B(n_63),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_243),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_260),
.B(n_28),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_262),
.B(n_30),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_297),
.B(n_31),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_212),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_229),
.B(n_34),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_267),
.B(n_40),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_281),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_235),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_335),
.B(n_403),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_330),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_347),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_335),
.B(n_308),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_352),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_356),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_354),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_336),
.B(n_238),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_356),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_356),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_364),
.B(n_372),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_354),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g437 ( 
.A1(n_400),
.A2(n_318),
.B1(n_284),
.B2(n_323),
.Y(n_437)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_391),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_333),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_374),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_334),
.Y(n_441)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_373),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_424),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_400),
.A2(n_318),
.B1(n_315),
.B2(n_320),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_332),
.B(n_197),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_376),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_373),
.Y(n_447)
);

NAND2xp33_ASAP7_75t_SL g448 ( 
.A(n_417),
.B(n_212),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_400),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_343),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_397),
.B(n_322),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_377),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_419),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_377),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_412),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_377),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_371),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_332),
.B(n_207),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_412),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_417),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_397),
.B(n_291),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_417),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_362),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_398),
.B(n_208),
.Y(n_464)
);

NAND2xp33_ASAP7_75t_L g465 ( 
.A(n_357),
.B(n_257),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_338),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_349),
.B(n_327),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_369),
.B(n_293),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_422),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_380),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_422),
.B(n_209),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_380),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_418),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_382),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_387),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_340),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_389),
.Y(n_477)
);

NOR2x1p5_ASAP7_75t_L g478 ( 
.A(n_343),
.B(n_265),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_389),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_340),
.Y(n_480)
);

NAND2xp33_ASAP7_75t_L g481 ( 
.A(n_398),
.B(n_215),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_383),
.B(n_216),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_345),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_384),
.B(n_224),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_396),
.B(n_227),
.Y(n_485)
);

INVxp33_ASAP7_75t_L g486 ( 
.A(n_410),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_399),
.B(n_408),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_404),
.B(n_228),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_346),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_405),
.B(n_406),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_405),
.B(n_230),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_346),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_353),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_353),
.Y(n_494)
);

NOR2x1p5_ASAP7_75t_L g495 ( 
.A(n_393),
.B(n_266),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_358),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_358),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_365),
.Y(n_498)
);

NAND3xp33_ASAP7_75t_L g499 ( 
.A(n_368),
.B(n_316),
.C(n_313),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_414),
.B(n_241),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_365),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_416),
.B(n_317),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_421),
.Y(n_503)
);

NOR3xp33_ASAP7_75t_L g504 ( 
.A(n_385),
.B(n_287),
.C(n_325),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_416),
.B(n_242),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_423),
.B(n_244),
.Y(n_506)
);

INVxp33_ASAP7_75t_L g507 ( 
.A(n_370),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_366),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_366),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_341),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_375),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_375),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_388),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_361),
.B(n_326),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_351),
.Y(n_515)
);

NOR3xp33_ASAP7_75t_L g516 ( 
.A(n_394),
.B(n_328),
.C(n_237),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_392),
.B(n_248),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_407),
.A2(n_392),
.B1(n_395),
.B2(n_355),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_395),
.B(n_250),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_350),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_331),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_344),
.A2(n_285),
.B1(n_263),
.B2(n_296),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_350),
.Y(n_523)
);

AO21x2_ASAP7_75t_L g524 ( 
.A1(n_402),
.A2(n_251),
.B(n_246),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_367),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_350),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_379),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_411),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_413),
.B(n_252),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_415),
.B(n_253),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_337),
.Y(n_531)
);

OR2x2_ASAP7_75t_SL g532 ( 
.A(n_381),
.B(n_266),
.Y(n_532)
);

NAND3xp33_ASAP7_75t_L g533 ( 
.A(n_363),
.B(n_258),
.C(n_256),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_337),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_443),
.Y(n_535)
);

OAI221xp5_ASAP7_75t_L g536 ( 
.A1(n_504),
.A2(n_448),
.B1(n_440),
.B2(n_516),
.C(n_453),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_425),
.B(n_331),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_428),
.B(n_393),
.Y(n_538)
);

NOR3xp33_ASAP7_75t_L g539 ( 
.A(n_522),
.B(n_390),
.C(n_348),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_L g540 ( 
.A(n_460),
.B(n_259),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_463),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_427),
.B(n_449),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_451),
.B(n_261),
.Y(n_543)
);

BUFx6f_ASAP7_75t_SL g544 ( 
.A(n_455),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_433),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_433),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_461),
.B(n_274),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_433),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_426),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_438),
.B(n_226),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_426),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_465),
.A2(n_386),
.B(n_378),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_459),
.B(n_278),
.Y(n_553)
);

BUFx5_ASAP7_75t_L g554 ( 
.A(n_463),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_457),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_442),
.Y(n_556)
);

BUFx6f_ASAP7_75t_SL g557 ( 
.A(n_507),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_439),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_438),
.B(n_268),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_442),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_473),
.B(n_288),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_441),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_462),
.B(n_294),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_469),
.B(n_298),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_462),
.B(n_301),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_432),
.B(n_270),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_441),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_462),
.B(n_303),
.Y(n_568)
);

AND2x6_ASAP7_75t_L g569 ( 
.A(n_447),
.B(n_430),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_450),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_447),
.B(n_310),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_434),
.B(n_311),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_445),
.A2(n_342),
.B1(n_213),
.B2(n_219),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_518),
.B(n_314),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_480),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_458),
.A2(n_285),
.B1(n_213),
.B2(n_219),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_437),
.B(n_292),
.Y(n_577)
);

INVx8_ASAP7_75t_L g578 ( 
.A(n_480),
.Y(n_578)
);

NOR2x1p5_ASAP7_75t_L g579 ( 
.A(n_533),
.B(n_348),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_466),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_503),
.B(n_378),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_450),
.B(n_420),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_483),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_L g584 ( 
.A(n_444),
.B(n_306),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_499),
.B(n_390),
.Y(n_585)
);

BUFx6f_ASAP7_75t_SL g586 ( 
.A(n_507),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_483),
.Y(n_587)
);

OAI22xp33_ASAP7_75t_L g588 ( 
.A1(n_486),
.A2(n_280),
.B1(n_300),
.B2(n_221),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_489),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_467),
.B(n_378),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_464),
.B(n_324),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_511),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_471),
.B(n_205),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_467),
.B(n_386),
.Y(n_594)
);

NOR3xp33_ASAP7_75t_L g595 ( 
.A(n_448),
.B(n_401),
.C(n_359),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_491),
.B(n_221),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_495),
.B(n_401),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_500),
.B(n_386),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_505),
.B(n_263),
.Y(n_599)
);

NOR2xp67_ASAP7_75t_L g600 ( 
.A(n_435),
.B(n_337),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_482),
.B(n_286),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_506),
.B(n_286),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_487),
.B(n_280),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_478),
.B(n_41),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_489),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_492),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_468),
.B(n_296),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_484),
.B(n_307),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_492),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_493),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_485),
.B(n_312),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_513),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_488),
.B(n_300),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_474),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_481),
.A2(n_360),
.B1(n_339),
.B2(n_44),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_517),
.B(n_519),
.Y(n_616)
);

CKINVDCx14_ASAP7_75t_R g617 ( 
.A(n_532),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_515),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_525),
.B(n_42),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_530),
.B(n_64),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_514),
.B(n_67),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_493),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_524),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_494),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_502),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_496),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_496),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_598),
.A2(n_524),
.B(n_490),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_535),
.B(n_497),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_605),
.B(n_498),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_542),
.B(n_498),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_536),
.A2(n_501),
.B1(n_508),
.B2(n_509),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_578),
.Y(n_633)
);

O2A1O1Ixp33_ASAP7_75t_L g634 ( 
.A1(n_607),
.A2(n_509),
.B(n_508),
.C(n_501),
.Y(n_634)
);

NAND3xp33_ASAP7_75t_SL g635 ( 
.A(n_595),
.B(n_529),
.C(n_476),
.Y(n_635)
);

NAND2x1p5_ASAP7_75t_L g636 ( 
.A(n_560),
.B(n_626),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_623),
.A2(n_512),
.B1(n_528),
.B2(n_527),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_542),
.B(n_528),
.Y(n_638)
);

O2A1O1Ixp33_ASAP7_75t_L g639 ( 
.A1(n_607),
.A2(n_527),
.B(n_534),
.C(n_531),
.Y(n_639)
);

CKINVDCx10_ASAP7_75t_R g640 ( 
.A(n_557),
.Y(n_640)
);

A2O1A1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_581),
.A2(n_526),
.B(n_523),
.C(n_520),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_545),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_603),
.B(n_43),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_555),
.B(n_46),
.Y(n_644)
);

A2O1A1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_581),
.A2(n_526),
.B(n_523),
.C(n_520),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_541),
.Y(n_646)
);

NOR3xp33_ASAP7_75t_L g647 ( 
.A(n_588),
.B(n_539),
.C(n_599),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_570),
.B(n_510),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_625),
.B(n_48),
.Y(n_649)
);

A2O1A1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_546),
.A2(n_548),
.B(n_551),
.C(n_549),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_556),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_543),
.B(n_49),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_543),
.B(n_50),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_600),
.B(n_52),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_626),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_550),
.B(n_52),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_618),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_578),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_563),
.A2(n_429),
.B(n_431),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_563),
.A2(n_472),
.B(n_436),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_578),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_565),
.A2(n_568),
.B(n_571),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_565),
.A2(n_472),
.B(n_436),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_559),
.B(n_56),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_554),
.B(n_456),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_619),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_566),
.B(n_57),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_568),
.A2(n_571),
.B(n_572),
.Y(n_668)
);

BUFx4f_ASAP7_75t_L g669 ( 
.A(n_604),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_602),
.A2(n_576),
.B1(n_627),
.B2(n_624),
.Y(n_670)
);

NOR3xp33_ASAP7_75t_L g671 ( 
.A(n_537),
.B(n_596),
.C(n_608),
.Y(n_671)
);

O2A1O1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_584),
.A2(n_577),
.B(n_585),
.C(n_611),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_544),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_538),
.B(n_57),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_582),
.B(n_73),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_569),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_591),
.B(n_74),
.Y(n_677)
);

OAI21xp33_ASAP7_75t_L g678 ( 
.A1(n_573),
.A2(n_613),
.B(n_601),
.Y(n_678)
);

BUFx2_ASAP7_75t_SL g679 ( 
.A(n_544),
.Y(n_679)
);

BUFx10_ASAP7_75t_L g680 ( 
.A(n_557),
.Y(n_680)
);

OR2x6_ASAP7_75t_L g681 ( 
.A(n_597),
.B(n_477),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_558),
.A2(n_479),
.B1(n_477),
.B2(n_475),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_575),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_575),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_553),
.B(n_84),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_562),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_567),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_580),
.Y(n_688)
);

O2A1O1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_574),
.A2(n_610),
.B(n_622),
.C(n_609),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_561),
.B(n_87),
.Y(n_690)
);

O2A1O1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_583),
.A2(n_589),
.B(n_587),
.C(n_606),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_592),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_593),
.A2(n_540),
.B1(n_616),
.B2(n_547),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_579),
.B(n_106),
.Y(n_694)
);

NOR2xp67_ASAP7_75t_L g695 ( 
.A(n_615),
.B(n_112),
.Y(n_695)
);

CKINVDCx6p67_ASAP7_75t_R g696 ( 
.A(n_586),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_621),
.A2(n_454),
.B(n_452),
.C(n_446),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_564),
.B(n_122),
.Y(n_698)
);

BUFx2_ASAP7_75t_SL g699 ( 
.A(n_586),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_631),
.A2(n_630),
.B1(n_632),
.B2(n_686),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_629),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_687),
.B(n_612),
.Y(n_702)
);

AOI21xp33_ASAP7_75t_SL g703 ( 
.A1(n_647),
.A2(n_617),
.B(n_620),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_688),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_680),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_696),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_657),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_633),
.B(n_614),
.Y(n_708)
);

AO31x2_ASAP7_75t_L g709 ( 
.A1(n_641),
.A2(n_470),
.A3(n_139),
.B(n_140),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_666),
.B(n_127),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_678),
.A2(n_670),
.B1(n_671),
.B2(n_643),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_661),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_679),
.B(n_148),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_661),
.Y(n_714)
);

NAND2x1p5_ASAP7_75t_L g715 ( 
.A(n_633),
.B(n_167),
.Y(n_715)
);

OAI21xp5_ASAP7_75t_L g716 ( 
.A1(n_650),
.A2(n_691),
.B(n_634),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_669),
.B(n_681),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_675),
.B(n_638),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_642),
.Y(n_719)
);

OAI21x1_ASAP7_75t_L g720 ( 
.A1(n_659),
.A2(n_660),
.B(n_663),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_644),
.Y(n_721)
);

NOR2x1_ASAP7_75t_R g722 ( 
.A(n_699),
.B(n_640),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_680),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_697),
.A2(n_639),
.B(n_677),
.Y(n_724)
);

A2O1A1Ixp33_ASAP7_75t_L g725 ( 
.A1(n_674),
.A2(n_672),
.B(n_652),
.C(n_653),
.Y(n_725)
);

OAI21xp5_ASAP7_75t_SL g726 ( 
.A1(n_649),
.A2(n_693),
.B(n_694),
.Y(n_726)
);

AOI221xp5_ASAP7_75t_L g727 ( 
.A1(n_635),
.A2(n_669),
.B1(n_673),
.B2(n_637),
.C(n_667),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_654),
.Y(n_728)
);

AOI21x1_ASAP7_75t_L g729 ( 
.A1(n_695),
.A2(n_664),
.B(n_656),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_654),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_681),
.B(n_658),
.Y(n_731)
);

AO21x1_ASAP7_75t_L g732 ( 
.A1(n_637),
.A2(n_685),
.B(n_698),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_658),
.B(n_655),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_636),
.Y(n_734)
);

AO31x2_ASAP7_75t_L g735 ( 
.A1(n_682),
.A2(n_690),
.A3(n_683),
.B(n_684),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_655),
.B(n_676),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_681),
.B(n_648),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_651),
.Y(n_738)
);

AO22x2_ASAP7_75t_L g739 ( 
.A1(n_646),
.A2(n_522),
.B1(n_647),
.B2(n_445),
.Y(n_739)
);

INVx4_ASAP7_75t_L g740 ( 
.A(n_692),
.Y(n_740)
);

OAI21xp5_ASAP7_75t_L g741 ( 
.A1(n_628),
.A2(n_552),
.B(n_662),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_629),
.B(n_451),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_629),
.B(n_451),
.Y(n_743)
);

AOI221xp5_ASAP7_75t_L g744 ( 
.A1(n_647),
.A2(n_536),
.B1(n_516),
.B2(n_678),
.C(n_504),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_629),
.B(n_451),
.Y(n_745)
);

A2O1A1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_668),
.A2(n_662),
.B(n_689),
.C(n_634),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_629),
.B(n_535),
.Y(n_747)
);

AO31x2_ASAP7_75t_L g748 ( 
.A1(n_641),
.A2(n_645),
.A3(n_628),
.B(n_552),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_629),
.B(n_451),
.Y(n_749)
);

AOI31xp67_ASAP7_75t_L g750 ( 
.A1(n_665),
.A2(n_598),
.A3(n_590),
.B(n_594),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_629),
.B(n_451),
.Y(n_751)
);

NOR3xp33_ASAP7_75t_L g752 ( 
.A(n_678),
.B(n_521),
.C(n_647),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_629),
.B(n_451),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_629),
.B(n_451),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_628),
.A2(n_552),
.B(n_662),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_629),
.B(n_451),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_629),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_629),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_629),
.Y(n_759)
);

AO31x2_ASAP7_75t_L g760 ( 
.A1(n_641),
.A2(n_645),
.A3(n_628),
.B(n_552),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_629),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_629),
.B(n_451),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_L g763 ( 
.A1(n_631),
.A2(n_630),
.B1(n_332),
.B2(n_632),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_631),
.A2(n_630),
.B1(n_332),
.B2(n_632),
.Y(n_764)
);

OAI22x1_ASAP7_75t_L g765 ( 
.A1(n_654),
.A2(n_393),
.B1(n_535),
.B2(n_495),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_631),
.A2(n_630),
.B1(n_332),
.B2(n_632),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_629),
.B(n_535),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_628),
.A2(n_552),
.B(n_662),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_686),
.B(n_687),
.Y(n_769)
);

OAI21xp5_ASAP7_75t_L g770 ( 
.A1(n_628),
.A2(n_552),
.B(n_662),
.Y(n_770)
);

AO31x2_ASAP7_75t_L g771 ( 
.A1(n_641),
.A2(n_645),
.A3(n_628),
.B(n_552),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_629),
.B(n_451),
.Y(n_772)
);

AO31x2_ASAP7_75t_L g773 ( 
.A1(n_641),
.A2(n_645),
.A3(n_628),
.B(n_552),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_647),
.A2(n_678),
.B1(n_670),
.B2(n_671),
.Y(n_774)
);

AND3x4_ASAP7_75t_L g775 ( 
.A(n_647),
.B(n_595),
.C(n_539),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_629),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_661),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_629),
.B(n_451),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_633),
.B(n_629),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_629),
.Y(n_780)
);

AO31x2_ASAP7_75t_L g781 ( 
.A1(n_641),
.A2(n_645),
.A3(n_628),
.B(n_552),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_628),
.A2(n_552),
.B(n_662),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_628),
.A2(n_552),
.B(n_662),
.Y(n_783)
);

BUFx12f_ASAP7_75t_L g784 ( 
.A(n_680),
.Y(n_784)
);

A2O1A1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_668),
.A2(n_662),
.B(n_689),
.C(n_634),
.Y(n_785)
);

NOR3xp33_ASAP7_75t_L g786 ( 
.A(n_678),
.B(n_521),
.C(n_647),
.Y(n_786)
);

OAI22x1_ASAP7_75t_L g787 ( 
.A1(n_654),
.A2(n_393),
.B1(n_535),
.B2(n_495),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_629),
.B(n_535),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_696),
.Y(n_789)
);

BUFx12f_ASAP7_75t_L g790 ( 
.A(n_784),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_779),
.B(n_731),
.Y(n_791)
);

BUFx12f_ASAP7_75t_L g792 ( 
.A(n_705),
.Y(n_792)
);

AOI332xp33_ASAP7_75t_L g793 ( 
.A1(n_757),
.A2(n_759),
.A3(n_776),
.B1(n_761),
.B2(n_788),
.B3(n_767),
.C1(n_747),
.C2(n_774),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_742),
.B(n_743),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_707),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_718),
.A2(n_725),
.B(n_774),
.Y(n_796)
);

BUFx2_ASAP7_75t_SL g797 ( 
.A(n_706),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_704),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_712),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_701),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_719),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_769),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_789),
.Y(n_803)
);

AO21x2_ASAP7_75t_L g804 ( 
.A1(n_741),
.A2(n_768),
.B(n_755),
.Y(n_804)
);

OAI21x1_ASAP7_75t_L g805 ( 
.A1(n_741),
.A2(n_770),
.B(n_768),
.Y(n_805)
);

AO21x2_ASAP7_75t_L g806 ( 
.A1(n_770),
.A2(n_783),
.B(n_782),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_769),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_SL g808 ( 
.A1(n_700),
.A2(n_763),
.B(n_764),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_720),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_758),
.B(n_780),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_745),
.B(n_749),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_746),
.A2(n_785),
.B(n_724),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_SL g813 ( 
.A(n_722),
.B(n_723),
.Y(n_813)
);

OAI21x1_ASAP7_75t_SL g814 ( 
.A1(n_700),
.A2(n_766),
.B(n_764),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_714),
.Y(n_815)
);

AOI21xp33_ASAP7_75t_L g816 ( 
.A1(n_726),
.A2(n_787),
.B(n_765),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_702),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_SL g818 ( 
.A1(n_739),
.A2(n_730),
.B1(n_717),
.B2(n_715),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_722),
.Y(n_819)
);

BUFx4f_ASAP7_75t_SL g820 ( 
.A(n_708),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_702),
.Y(n_821)
);

NAND2x1p5_ASAP7_75t_L g822 ( 
.A(n_740),
.B(n_734),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_751),
.B(n_753),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_740),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_SL g825 ( 
.A1(n_739),
.A2(n_728),
.B1(n_713),
.B2(n_721),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_711),
.A2(n_716),
.B(n_744),
.C(n_726),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_748),
.Y(n_827)
);

INVx1_ASAP7_75t_SL g828 ( 
.A(n_737),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_748),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_754),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_738),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_756),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_762),
.Y(n_833)
);

OAI211xp5_ASAP7_75t_L g834 ( 
.A1(n_727),
.A2(n_786),
.B(n_752),
.C(n_703),
.Y(n_834)
);

OAI21x1_ASAP7_75t_SL g835 ( 
.A1(n_729),
.A2(n_732),
.B(n_710),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_772),
.Y(n_836)
);

OAI21x1_ASAP7_75t_L g837 ( 
.A1(n_736),
.A2(n_733),
.B(n_773),
.Y(n_837)
);

OA21x2_ASAP7_75t_L g838 ( 
.A1(n_748),
.A2(n_771),
.B(n_773),
.Y(n_838)
);

INVxp67_ASAP7_75t_SL g839 ( 
.A(n_778),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_775),
.Y(n_840)
);

OAI21x1_ASAP7_75t_L g841 ( 
.A1(n_760),
.A2(n_781),
.B(n_771),
.Y(n_841)
);

AO21x2_ASAP7_75t_L g842 ( 
.A1(n_771),
.A2(n_781),
.B(n_709),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_735),
.A2(n_535),
.B1(n_393),
.B2(n_763),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_757),
.B(n_759),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_747),
.B(n_678),
.Y(n_845)
);

AOI221xp5_ASAP7_75t_L g846 ( 
.A1(n_763),
.A2(n_536),
.B1(n_766),
.B2(n_764),
.C(n_744),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_747),
.B(n_678),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_SL g848 ( 
.A1(n_763),
.A2(n_764),
.B1(n_766),
.B2(n_393),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_757),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_757),
.Y(n_850)
);

O2A1O1Ixp33_ASAP7_75t_SL g851 ( 
.A1(n_746),
.A2(n_785),
.B(n_725),
.C(n_764),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_777),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_750),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_706),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_747),
.Y(n_855)
);

NAND2xp33_ASAP7_75t_SL g856 ( 
.A(n_763),
.B(n_764),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_809),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_802),
.B(n_807),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_820),
.Y(n_859)
);

CKINVDCx11_ASAP7_75t_R g860 ( 
.A(n_790),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_817),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_790),
.Y(n_862)
);

AO21x2_ASAP7_75t_L g863 ( 
.A1(n_812),
.A2(n_814),
.B(n_835),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_846),
.B(n_826),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_810),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_820),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_826),
.B(n_796),
.Y(n_867)
);

CKINVDCx16_ASAP7_75t_R g868 ( 
.A(n_813),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_848),
.A2(n_808),
.B1(n_843),
.B2(n_821),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_856),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_805),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_852),
.B(n_837),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_798),
.B(n_801),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_804),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_800),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_804),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_806),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_806),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_856),
.B(n_839),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_828),
.B(n_845),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_819),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_853),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_799),
.Y(n_883)
);

A2O1A1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_834),
.A2(n_816),
.B(n_793),
.C(n_823),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_795),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_827),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_799),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_840),
.B(n_855),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_815),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_824),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_829),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_792),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_851),
.B(n_845),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_847),
.B(n_791),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_886),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_874),
.B(n_876),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_872),
.B(n_863),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_870),
.B(n_838),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_891),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_870),
.B(n_838),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_877),
.B(n_841),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_880),
.B(n_841),
.Y(n_902)
);

AOI221xp5_ASAP7_75t_L g903 ( 
.A1(n_884),
.A2(n_823),
.B1(n_811),
.B2(n_847),
.C(n_830),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_878),
.B(n_842),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_868),
.B(n_818),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_880),
.B(n_849),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_867),
.B(n_825),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_873),
.B(n_850),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_867),
.B(n_864),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_873),
.B(n_831),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_861),
.B(n_894),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_890),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_857),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_864),
.B(n_836),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_861),
.B(n_844),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_858),
.B(n_885),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_910),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_898),
.B(n_871),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_898),
.B(n_900),
.Y(n_919)
);

AOI222xp33_ASAP7_75t_L g920 ( 
.A1(n_903),
.A2(n_840),
.B1(n_869),
.B2(n_832),
.C1(n_833),
.C2(n_811),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_902),
.B(n_899),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_899),
.Y(n_922)
);

OR2x2_ASAP7_75t_L g923 ( 
.A(n_902),
.B(n_879),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_895),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_900),
.B(n_871),
.Y(n_925)
);

INVxp67_ASAP7_75t_SL g926 ( 
.A(n_913),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_911),
.B(n_865),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_897),
.B(n_863),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_910),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_916),
.B(n_885),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_916),
.B(n_883),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_901),
.B(n_882),
.Y(n_932)
);

OR2x2_ASAP7_75t_L g933 ( 
.A(n_921),
.B(n_896),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_919),
.B(n_918),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_917),
.B(n_908),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_921),
.B(n_931),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_924),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_926),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_929),
.B(n_930),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_928),
.B(n_897),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_928),
.B(n_897),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_927),
.B(n_908),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_931),
.B(n_896),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_927),
.B(n_907),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_L g945 ( 
.A1(n_920),
.A2(n_840),
.B1(n_903),
.B2(n_869),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_SL g946 ( 
.A(n_922),
.B(n_868),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_932),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_919),
.B(n_904),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_944),
.B(n_918),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_938),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_937),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_936),
.B(n_923),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_938),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_934),
.B(n_928),
.Y(n_954)
);

NAND2x1p5_ASAP7_75t_L g955 ( 
.A(n_940),
.B(n_912),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_934),
.B(n_928),
.Y(n_956)
);

INVxp67_ASAP7_75t_SL g957 ( 
.A(n_947),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_937),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_948),
.B(n_925),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_948),
.B(n_925),
.Y(n_960)
);

OAI22xp33_ASAP7_75t_SL g961 ( 
.A1(n_957),
.A2(n_946),
.B1(n_905),
.B2(n_936),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_952),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_950),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_952),
.Y(n_964)
);

NAND3xp33_ASAP7_75t_L g965 ( 
.A(n_953),
.B(n_945),
.C(n_840),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_951),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_954),
.A2(n_909),
.B1(n_894),
.B2(n_907),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_954),
.B(n_940),
.Y(n_968)
);

NOR2x1_ASAP7_75t_L g969 ( 
.A(n_956),
.B(n_797),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_956),
.A2(n_941),
.B1(n_940),
.B2(n_939),
.Y(n_970)
);

OAI21xp33_ASAP7_75t_L g971 ( 
.A1(n_949),
.A2(n_943),
.B(n_933),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_951),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_958),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_963),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_971),
.B(n_959),
.Y(n_975)
);

AOI211xp5_ASAP7_75t_SL g976 ( 
.A1(n_961),
.A2(n_893),
.B(n_909),
.C(n_888),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_966),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_972),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_973),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_975),
.B(n_962),
.Y(n_980)
);

NAND4xp25_ASAP7_75t_L g981 ( 
.A(n_976),
.B(n_965),
.C(n_969),
.D(n_967),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_974),
.A2(n_963),
.B(n_970),
.Y(n_982)
);

OAI21xp33_ASAP7_75t_L g983 ( 
.A1(n_974),
.A2(n_967),
.B(n_964),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_978),
.A2(n_955),
.B1(n_968),
.B2(n_960),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_977),
.B(n_955),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_979),
.B(n_860),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_986),
.B(n_892),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_983),
.B(n_980),
.Y(n_988)
);

OAI221xp5_ASAP7_75t_L g989 ( 
.A1(n_981),
.A2(n_892),
.B1(n_977),
.B2(n_819),
.C(n_955),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_984),
.B(n_862),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_982),
.B(n_959),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_985),
.B(n_803),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_990),
.B(n_803),
.Y(n_993)
);

NOR2x1p5_ASAP7_75t_L g994 ( 
.A(n_988),
.B(n_854),
.Y(n_994)
);

NOR3xp33_ASAP7_75t_L g995 ( 
.A(n_989),
.B(n_854),
.C(n_881),
.Y(n_995)
);

NOR2x1_ASAP7_75t_L g996 ( 
.A(n_992),
.B(n_866),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_991),
.A2(n_875),
.B(n_859),
.C(n_889),
.Y(n_997)
);

NAND2x1p5_ASAP7_75t_L g998 ( 
.A(n_996),
.B(n_866),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_997),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_994),
.Y(n_1000)
);

NOR2x1_ASAP7_75t_L g1001 ( 
.A(n_993),
.B(n_987),
.Y(n_1001)
);

NOR2x1_ASAP7_75t_L g1002 ( 
.A(n_995),
.B(n_866),
.Y(n_1002)
);

NAND2x1p5_ASAP7_75t_L g1003 ( 
.A(n_1002),
.B(n_792),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_1001),
.B(n_941),
.Y(n_1004)
);

XOR2xp5_ASAP7_75t_L g1005 ( 
.A(n_1003),
.B(n_1000),
.Y(n_1005)
);

OR4x1_ASAP7_75t_L g1006 ( 
.A(n_1003),
.B(n_999),
.C(n_998),
.D(n_859),
.Y(n_1006)
);

INVxp67_ASAP7_75t_SL g1007 ( 
.A(n_1005),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_1006),
.A2(n_1004),
.B1(n_914),
.B2(n_887),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_1007),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_1009),
.A2(n_1008),
.B1(n_914),
.B2(n_915),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_1009),
.A2(n_794),
.B(n_883),
.Y(n_1011)
);

OA21x2_ASAP7_75t_L g1012 ( 
.A1(n_1011),
.A2(n_942),
.B(n_935),
.Y(n_1012)
);

BUFx24_ASAP7_75t_SL g1013 ( 
.A(n_1012),
.Y(n_1013)
);

AO21x2_ASAP7_75t_L g1014 ( 
.A1(n_1013),
.A2(n_1010),
.B(n_791),
.Y(n_1014)
);

AOI21xp33_ASAP7_75t_SL g1015 ( 
.A1(n_1014),
.A2(n_906),
.B(n_822),
.Y(n_1015)
);


endmodule