module fake_jpeg_10803_n_644 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_644);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_644;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_59),
.Y(n_143)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_28),
.B(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_63),
.B(n_68),
.Y(n_136)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_56),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_65),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_52),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_69),
.Y(n_148)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_71),
.Y(n_203)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_28),
.B(n_15),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_74),
.B(n_80),
.Y(n_140)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_75),
.Y(n_175)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_76),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_77),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_29),
.B(n_15),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g135 ( 
.A(n_81),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_82),
.B(n_86),
.Y(n_200)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_43),
.B(n_13),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_87),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_89),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_91),
.Y(n_177)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_94),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_96),
.Y(n_205)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_13),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_100),
.B(n_104),
.Y(n_202)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

BUFx10_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_42),
.B(n_12),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_105),
.Y(n_181)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_107),
.Y(n_184)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_34),
.Y(n_108)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_108),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_25),
.B(n_12),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_109),
.B(n_57),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_50),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_112),
.B(n_116),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_31),
.Y(n_113)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_57),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_25),
.B(n_12),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_17),
.Y(n_117)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_17),
.Y(n_118)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_36),
.Y(n_119)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_17),
.Y(n_120)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_36),
.Y(n_121)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_47),
.Y(n_122)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_17),
.Y(n_123)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_26),
.B(n_12),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_124),
.B(n_58),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_67),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_125),
.A2(n_132),
.B1(n_142),
.B2(n_158),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_68),
.B(n_26),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_129),
.B(n_137),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_131),
.B(n_190),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_71),
.A2(n_44),
.B1(n_51),
.B2(n_45),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_68),
.B(n_33),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_89),
.A2(n_44),
.B1(n_38),
.B2(n_51),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g257 ( 
.A1(n_139),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_66),
.A2(n_103),
.B1(n_77),
.B2(n_70),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_75),
.B(n_23),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_145),
.B(n_65),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_92),
.B(n_58),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_149),
.B(n_179),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_155),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_66),
.A2(n_23),
.B1(n_17),
.B2(n_22),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_77),
.A2(n_23),
.B1(n_22),
.B2(n_18),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_171),
.A2(n_180),
.B1(n_182),
.B2(n_204),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_73),
.A2(n_33),
.B1(n_22),
.B2(n_18),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_78),
.A2(n_18),
.B1(n_38),
.B2(n_53),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_59),
.Y(n_183)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_69),
.Y(n_185)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_76),
.Y(n_188)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_79),
.A2(n_23),
.B1(n_38),
.B2(n_53),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_192),
.A2(n_39),
.B1(n_32),
.B2(n_49),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_108),
.A2(n_21),
.B(n_54),
.C(n_53),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_197),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_84),
.B(n_21),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_81),
.A2(n_21),
.B1(n_54),
.B2(n_30),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_206),
.Y(n_281)
);

INVx4_ASAP7_75t_SL g208 ( 
.A(n_199),
.Y(n_208)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_208),
.Y(n_302)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_209),
.Y(n_299)
);

BUFx8_ASAP7_75t_L g211 ( 
.A(n_133),
.Y(n_211)
);

BUFx8_ASAP7_75t_L g292 ( 
.A(n_211),
.Y(n_292)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_146),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_212),
.Y(n_297)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_213),
.Y(n_309)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_214),
.Y(n_340)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_216),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_193),
.A2(n_103),
.B1(n_91),
.B2(n_87),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_217),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_133),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_218),
.B(n_260),
.Y(n_329)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_143),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_220),
.Y(n_301)
);

BUFx8_ASAP7_75t_L g221 ( 
.A(n_133),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_221),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_223),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_153),
.A2(n_95),
.B1(n_88),
.B2(n_122),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_224),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_199),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_225),
.B(n_236),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_226),
.Y(n_310)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_228),
.Y(n_290)
);

BUFx2_ASAP7_75t_SL g229 ( 
.A(n_177),
.Y(n_229)
);

INVx11_ASAP7_75t_L g338 ( 
.A(n_229),
.Y(n_338)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_231),
.Y(n_298)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_162),
.Y(n_232)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_232),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_141),
.Y(n_233)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_233),
.Y(n_312)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_134),
.Y(n_234)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_234),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_136),
.A2(n_106),
.B1(n_96),
.B2(n_105),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_235),
.A2(n_276),
.B1(n_40),
.B2(n_172),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_147),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_170),
.Y(n_238)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_238),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_141),
.Y(n_239)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_239),
.Y(n_322)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_240),
.Y(n_325)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_148),
.Y(n_241)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_241),
.Y(n_327)
);

BUFx2_ASAP7_75t_SL g242 ( 
.A(n_126),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_242),
.Y(n_323)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_165),
.Y(n_243)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_243),
.Y(n_334)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_160),
.Y(n_244)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_244),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g245 ( 
.A(n_155),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_245),
.Y(n_333)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_246),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_247),
.A2(n_253),
.B1(n_264),
.B2(n_265),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_145),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_248),
.B(n_249),
.Y(n_304)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_186),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_190),
.A2(n_121),
.B1(n_119),
.B2(n_114),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_251),
.A2(n_271),
.B1(n_279),
.B2(n_280),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_139),
.A2(n_90),
.B1(n_93),
.B2(n_110),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_252),
.A2(n_135),
.B1(n_171),
.B2(n_152),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g253 ( 
.A(n_175),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_138),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_254),
.B(n_256),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_136),
.B(n_94),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_255),
.B(n_261),
.C(n_263),
.Y(n_332)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_164),
.Y(n_256)
);

OA22x2_ASAP7_75t_L g288 ( 
.A1(n_257),
.A2(n_277),
.B1(n_35),
.B2(n_40),
.Y(n_288)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_178),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_258),
.B(n_259),
.Y(n_330)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_166),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_182),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_139),
.B(n_115),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_151),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_266),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_202),
.B(n_130),
.C(n_128),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_181),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_194),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_154),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_200),
.B(n_50),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_267),
.B(n_273),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_173),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_268),
.A2(n_270),
.B1(n_274),
.B2(n_278),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_202),
.B(n_118),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_269),
.B(n_0),
.C(n_1),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_159),
.A2(n_23),
.B1(n_54),
.B2(n_49),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_132),
.A2(n_113),
.B1(n_39),
.B2(n_35),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_180),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_156),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_200),
.B(n_50),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_142),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_125),
.A2(n_23),
.B1(n_39),
.B2(n_49),
.Y(n_276)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_191),
.Y(n_278)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_203),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_158),
.A2(n_201),
.B1(n_187),
.B2(n_157),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_283),
.A2(n_285),
.B1(n_295),
.B2(n_303),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_227),
.A2(n_219),
.B(n_261),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_284),
.A2(n_289),
.B(n_308),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_263),
.A2(n_150),
.B1(n_144),
.B2(n_152),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_287),
.B(n_4),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_288),
.B(n_315),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_261),
.A2(n_161),
.B(n_30),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_248),
.A2(n_140),
.B1(n_127),
.B2(n_150),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_237),
.A2(n_140),
.B1(n_144),
.B2(n_205),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_195),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_305),
.B(n_311),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_215),
.A2(n_205),
.B1(n_135),
.B2(n_157),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_307),
.A2(n_318),
.B1(n_213),
.B2(n_214),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_226),
.A2(n_40),
.B(n_32),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_269),
.B(n_172),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_226),
.A2(n_255),
.B(n_245),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_314),
.A2(n_324),
.B(n_207),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_L g318 ( 
.A1(n_277),
.A2(n_257),
.B1(n_235),
.B2(n_276),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_255),
.A2(n_50),
.B(n_57),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_207),
.A2(n_50),
.B1(n_1),
.B2(n_2),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_328),
.A2(n_315),
.B1(n_313),
.B2(n_302),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_250),
.B(n_0),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_335),
.C(n_336),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_272),
.B(n_0),
.Y(n_336)
);

AO22x1_ASAP7_75t_L g341 ( 
.A1(n_257),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_341),
.B(n_1),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_317),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_342),
.B(n_356),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_338),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_344),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_345),
.A2(n_354),
.B1(n_363),
.B2(n_366),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_346),
.Y(n_408)
);

NAND2xp33_ASAP7_75t_R g347 ( 
.A(n_305),
.B(n_311),
.Y(n_347)
);

OAI21xp33_ASAP7_75t_SL g407 ( 
.A1(n_347),
.A2(n_327),
.B(n_337),
.Y(n_407)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_325),
.Y(n_348)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_348),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_282),
.A2(n_257),
.B1(n_278),
.B2(n_212),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_349),
.A2(n_350),
.B(n_370),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_282),
.B(n_208),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_287),
.A2(n_223),
.B(n_268),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_351),
.A2(n_338),
.B(n_322),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_206),
.C(n_210),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_352),
.B(n_367),
.C(n_372),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_313),
.A2(n_228),
.B1(n_279),
.B2(n_232),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_325),
.Y(n_355)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_355),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_330),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_308),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_357),
.B(n_369),
.Y(n_422)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_301),
.Y(n_359)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_359),
.Y(n_406)
);

NOR3xp33_ASAP7_75t_SL g360 ( 
.A(n_329),
.B(n_284),
.C(n_341),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_360),
.B(n_378),
.Y(n_416)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_334),
.Y(n_362)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_362),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_318),
.A2(n_247),
.B1(n_264),
.B2(n_209),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_364),
.A2(n_375),
.B1(n_383),
.B2(n_385),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g394 ( 
.A(n_365),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_332),
.A2(n_265),
.B1(n_240),
.B2(n_243),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_310),
.B(n_222),
.C(n_230),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_296),
.B(n_244),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_368),
.B(n_323),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_304),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_303),
.A2(n_246),
.B1(n_220),
.B2(n_241),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_314),
.A2(n_289),
.B1(n_288),
.B2(n_307),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_371),
.A2(n_374),
.B1(n_382),
.B2(n_297),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_324),
.B(n_231),
.C(n_239),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_288),
.A2(n_233),
.B1(n_249),
.B2(n_221),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_285),
.A2(n_221),
.B1(n_211),
.B2(n_4),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_334),
.Y(n_376)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

O2A1O1Ixp33_ASAP7_75t_L g377 ( 
.A1(n_291),
.A2(n_211),
.B(n_3),
.C(n_4),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_377),
.A2(n_384),
.B(n_300),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_319),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_298),
.Y(n_379)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_379),
.Y(n_421)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_298),
.Y(n_380)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_380),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_333),
.B(n_1),
.C(n_4),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_381),
.B(n_321),
.C(n_286),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_341),
.A2(n_291),
.B1(n_326),
.B2(n_288),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_295),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_326),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_302),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_386),
.A2(n_387),
.B1(n_337),
.B2(n_327),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_335),
.A2(n_7),
.B1(n_10),
.B2(n_316),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_328),
.B(n_10),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_388),
.B(n_286),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_389),
.B(n_342),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_374),
.A2(n_290),
.B1(n_306),
.B2(n_293),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_391),
.A2(n_427),
.B1(n_429),
.B2(n_281),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_368),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_392),
.B(n_414),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_361),
.A2(n_339),
.B1(n_319),
.B2(n_290),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_395),
.A2(n_399),
.B1(n_403),
.B2(n_411),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_358),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_396),
.B(n_410),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_397),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_361),
.A2(n_364),
.B1(n_349),
.B2(n_357),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_352),
.B(n_336),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_400),
.B(n_281),
.C(n_309),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_358),
.A2(n_316),
.B1(n_320),
.B2(n_306),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_350),
.A2(n_294),
.B(n_293),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_404),
.A2(n_346),
.B(n_377),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_407),
.A2(n_412),
.B(n_351),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_358),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_350),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_352),
.B(n_331),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_415),
.B(n_428),
.C(n_400),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_417),
.B(n_419),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_386),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_418),
.B(n_354),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_370),
.A2(n_297),
.B1(n_301),
.B2(n_321),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_425),
.A2(n_366),
.B1(n_377),
.B2(n_376),
.Y(n_440)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_348),
.Y(n_426)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_426),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_358),
.A2(n_297),
.B1(n_301),
.B2(n_340),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_367),
.B(n_353),
.Y(n_428)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_430),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_429),
.A2(n_363),
.B1(n_375),
.B2(n_365),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_431),
.A2(n_446),
.B1(n_454),
.B2(n_463),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_433),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_398),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_434),
.B(n_435),
.Y(n_484)
);

OAI32xp33_ASAP7_75t_L g435 ( 
.A1(n_416),
.A2(n_373),
.A3(n_347),
.B1(n_371),
.B2(n_384),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_389),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_436),
.Y(n_483)
);

OAI32xp33_ASAP7_75t_L g437 ( 
.A1(n_416),
.A2(n_373),
.A3(n_360),
.B1(n_345),
.B2(n_343),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_437),
.B(n_443),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_367),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_438),
.B(n_441),
.C(n_457),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_395),
.A2(n_382),
.B1(n_378),
.B2(n_372),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_439),
.A2(n_466),
.B(n_424),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_440),
.A2(n_455),
.B1(n_458),
.B2(n_459),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_392),
.B(n_380),
.Y(n_442)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_442),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_445),
.B(n_465),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_396),
.A2(n_343),
.B1(n_383),
.B2(n_360),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_402),
.Y(n_447)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_447),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_379),
.Y(n_451)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_451),
.Y(n_501)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_402),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_453),
.B(n_456),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_410),
.A2(n_385),
.B1(n_387),
.B2(n_356),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_399),
.A2(n_388),
.B1(n_355),
.B2(n_362),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_405),
.Y(n_456)
);

MAJx2_ASAP7_75t_L g457 ( 
.A(n_409),
.B(n_353),
.C(n_381),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_SL g458 ( 
.A1(n_403),
.A2(n_344),
.B1(n_359),
.B2(n_322),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_401),
.A2(n_388),
.B1(n_381),
.B2(n_344),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_405),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_461),
.Y(n_496)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_413),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_394),
.B(n_388),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_464),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_412),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_413),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_408),
.A2(n_312),
.B(n_292),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_467),
.B(n_420),
.C(n_423),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_451),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_471),
.B(n_472),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_442),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_441),
.B(n_428),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_473),
.B(n_474),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_448),
.B(n_415),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_448),
.B(n_422),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_475),
.B(n_480),
.C(n_485),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_434),
.B(n_398),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_477),
.B(n_481),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_438),
.B(n_422),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g516 ( 
.A(n_479),
.B(n_482),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_407),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_449),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_457),
.B(n_419),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_437),
.B(n_417),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_435),
.B(n_419),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_493),
.C(n_498),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g489 ( 
.A(n_446),
.B(n_393),
.Y(n_489)
);

XOR2x2_ASAP7_75t_L g523 ( 
.A(n_489),
.B(n_431),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_439),
.A2(n_393),
.B1(n_390),
.B2(n_391),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_490),
.A2(n_492),
.B1(n_498),
.B2(n_469),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_450),
.B(n_390),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_432),
.A2(n_418),
.B1(n_394),
.B2(n_397),
.Y(n_495)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_495),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_445),
.B(n_426),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_497),
.B(n_423),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_432),
.B(n_404),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_499),
.B(n_444),
.C(n_465),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_502),
.A2(n_433),
.B(n_464),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_476),
.A2(n_440),
.B1(n_430),
.B2(n_459),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_505),
.A2(n_529),
.B1(n_530),
.B2(n_501),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_506),
.A2(n_526),
.B(n_292),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_491),
.Y(n_507)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_507),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_508),
.B(n_514),
.C(n_515),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_502),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_509),
.B(n_532),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_476),
.A2(n_452),
.B1(n_455),
.B2(n_443),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_510),
.A2(n_490),
.B1(n_469),
.B2(n_478),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_SL g512 ( 
.A(n_486),
.B(n_452),
.C(n_462),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_512),
.B(n_524),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_473),
.B(n_466),
.C(n_454),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_470),
.B(n_461),
.C(n_460),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_470),
.B(n_456),
.C(n_453),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_517),
.B(n_520),
.C(n_488),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_474),
.B(n_447),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_518),
.B(n_523),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_499),
.B(n_444),
.C(n_420),
.Y(n_520)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_468),
.Y(n_522)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_522),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_484),
.B(n_312),
.Y(n_524)
);

INVx11_ASAP7_75t_L g525 ( 
.A(n_483),
.Y(n_525)
);

CKINVDCx16_ASAP7_75t_R g539 ( 
.A(n_525),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_478),
.A2(n_486),
.B(n_500),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_527),
.A2(n_521),
.B1(n_514),
.B2(n_509),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_528),
.B(n_531),
.Y(n_551)
);

AOI22x1_ASAP7_75t_L g529 ( 
.A1(n_484),
.A2(n_425),
.B1(n_401),
.B2(n_411),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_487),
.A2(n_421),
.B1(n_424),
.B2(n_406),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_494),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_487),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_475),
.B(n_421),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_533),
.B(n_491),
.Y(n_555)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_534),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_538),
.A2(n_548),
.B1(n_556),
.B2(n_527),
.Y(n_565)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_540),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_511),
.B(n_483),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_541),
.B(n_508),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_542),
.B(n_543),
.C(n_547),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_515),
.B(n_485),
.C(n_479),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_507),
.B(n_501),
.Y(n_545)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_545),
.Y(n_571)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_513),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_546),
.B(n_559),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_517),
.B(n_480),
.C(n_482),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_523),
.A2(n_493),
.B1(n_500),
.B2(n_489),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_507),
.B(n_496),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_549),
.B(n_526),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_519),
.B(n_496),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_550),
.B(n_554),
.Y(n_569)
);

XNOR2x1_ASAP7_75t_L g554 ( 
.A(n_504),
.B(n_494),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_555),
.B(n_558),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_510),
.A2(n_406),
.B1(n_309),
.B2(n_340),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_557),
.A2(n_540),
.B(n_556),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_518),
.B(n_299),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_525),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_551),
.B(n_536),
.Y(n_560)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_560),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_561),
.B(n_563),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_565),
.B(n_548),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_535),
.B(n_520),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_566),
.B(n_568),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_537),
.B(n_519),
.C(n_503),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_536),
.A2(n_506),
.B(n_512),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_572),
.A2(n_573),
.B(n_575),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_555),
.B(n_533),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_552),
.B(n_504),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_557),
.A2(n_529),
.B(n_503),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_576),
.A2(n_580),
.B(n_558),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_544),
.B(n_529),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_577),
.B(n_578),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_545),
.B(n_549),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_535),
.B(n_516),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_579),
.B(n_553),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_561),
.Y(n_583)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_583),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_566),
.B(n_537),
.C(n_542),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_584),
.B(n_586),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_562),
.A2(n_552),
.B1(n_539),
.B2(n_550),
.Y(n_585)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_585),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_575),
.B(n_538),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_560),
.B(n_553),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_587),
.B(n_588),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_589),
.B(n_598),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_L g603 ( 
.A1(n_590),
.A2(n_578),
.B(n_570),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_564),
.B(n_543),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_591),
.B(n_593),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_577),
.B(n_547),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_565),
.B(n_516),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_594),
.B(n_595),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_568),
.B(n_554),
.C(n_299),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_580),
.B(n_292),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_596),
.A2(n_572),
.B(n_563),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_600),
.A2(n_603),
.B(n_608),
.Y(n_620)
);

FAx1_ASAP7_75t_SL g602 ( 
.A(n_592),
.B(n_579),
.CI(n_576),
.CON(n_602),
.SN(n_602)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_602),
.B(n_610),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_581),
.A2(n_570),
.B(n_571),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_584),
.B(n_562),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_597),
.B(n_567),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_611),
.B(n_612),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_582),
.B(n_567),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_SL g613 ( 
.A1(n_585),
.A2(n_571),
.B1(n_569),
.B2(n_573),
.Y(n_613)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_613),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_606),
.B(n_587),
.Y(n_614)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_614),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_599),
.B(n_589),
.Y(n_615)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_615),
.A2(n_602),
.B(n_609),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_SL g616 ( 
.A1(n_600),
.A2(n_595),
.B(n_590),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_616),
.B(n_621),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_605),
.A2(n_607),
.B(n_608),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_601),
.Y(n_622)
);

AO21x1_ASAP7_75t_L g626 ( 
.A1(n_622),
.A2(n_604),
.B(n_602),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_601),
.B(n_603),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_623),
.B(n_624),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_609),
.B(n_588),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_626),
.B(n_620),
.C(n_624),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_628),
.B(n_629),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_SL g629 ( 
.A1(n_618),
.A2(n_604),
.B(n_569),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_617),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_L g635 ( 
.A1(n_630),
.A2(n_631),
.B(n_620),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_SL g631 ( 
.A(n_619),
.B(n_598),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_SL g633 ( 
.A1(n_625),
.A2(n_632),
.B(n_627),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_633),
.B(n_635),
.Y(n_638)
);

NAND2x1_ASAP7_75t_SL g637 ( 
.A(n_636),
.B(n_627),
.Y(n_637)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_637),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_634),
.A2(n_622),
.B1(n_574),
.B2(n_292),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_639),
.B(n_574),
.C(n_10),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_641),
.A2(n_638),
.B(n_637),
.Y(n_642)
);

XNOR2xp5_ASAP7_75t_L g643 ( 
.A(n_642),
.B(n_640),
.Y(n_643)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_643),
.B(n_10),
.Y(n_644)
);


endmodule