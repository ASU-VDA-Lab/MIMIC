module fake_jpeg_18374_n_322 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_322);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

CKINVDCx6p67_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_5),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_33),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_34),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_35),
.B(n_16),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_26),
.A2(n_21),
.B1(n_17),
.B2(n_18),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_28),
.B1(n_16),
.B2(n_11),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_32),
.B(n_34),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_20),
.B(n_13),
.Y(n_74)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_29),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_55),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_37),
.B1(n_16),
.B2(n_14),
.Y(n_72)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_29),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_59),
.Y(n_63)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_24),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_37),
.Y(n_75)
);

AO22x2_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_28),
.B1(n_41),
.B2(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_72),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_42),
.C(n_44),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_70),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_28),
.B1(n_36),
.B2(n_41),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_60),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_41),
.B1(n_40),
.B2(n_27),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_40),
.B1(n_27),
.B2(n_37),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_44),
.C(n_31),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_74),
.B(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_54),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_30),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_99),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_54),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_62),
.B1(n_48),
.B2(n_50),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_95),
.Y(n_106)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_24),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_11),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_74),
.B1(n_30),
.B2(n_75),
.Y(n_102)
);

BUFx10_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_102),
.A2(n_105),
.B(n_112),
.Y(n_141)
);

AO22x1_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_62),
.B1(n_67),
.B2(n_69),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_109),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_108),
.A2(n_119),
.B1(n_98),
.B2(n_29),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_65),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_110),
.B(n_113),
.Y(n_162)
);

XOR2x2_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_62),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_99),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_68),
.B1(n_21),
.B2(n_48),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_71),
.B(n_52),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_125),
.B(n_127),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_68),
.B1(n_71),
.B2(n_60),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_82),
.A2(n_55),
.B1(n_21),
.B2(n_17),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_124),
.B1(n_128),
.B2(n_18),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_31),
.C(n_24),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_96),
.C(n_90),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_55),
.B1(n_21),
.B2(n_17),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_31),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_83),
.A2(n_14),
.B(n_12),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_92),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_136),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_87),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_131),
.B(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_90),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_135),
.B(n_139),
.Y(n_194)
);

AOI32xp33_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_96),
.A3(n_97),
.B1(n_85),
.B2(n_99),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_159),
.C(n_164),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_143),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_111),
.B(n_96),
.Y(n_139)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_98),
.B(n_88),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_151),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_94),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_144),
.B(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_146),
.Y(n_176)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_155),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_101),
.B(n_94),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_160),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_115),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_125),
.B1(n_124),
.B2(n_121),
.Y(n_180)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_112),
.A2(n_98),
.B1(n_19),
.B2(n_18),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_158),
.A2(n_127),
.B1(n_108),
.B2(n_129),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_98),
.C(n_24),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_104),
.B(n_33),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_149),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_104),
.B(n_13),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_165),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_24),
.C(n_33),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_47),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_167),
.B(n_174),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_160),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_158),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_146),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_120),
.Y(n_175)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_113),
.Y(n_177)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

NOR2x1_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_107),
.Y(n_178)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_179),
.A2(n_19),
.B1(n_12),
.B2(n_16),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_180),
.A2(n_135),
.B1(n_142),
.B2(n_143),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_154),
.A2(n_116),
.B1(n_102),
.B2(n_128),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_186),
.A2(n_187),
.B(n_142),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_154),
.A2(n_102),
.B1(n_33),
.B2(n_30),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_102),
.Y(n_189)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_162),
.C(n_141),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_164),
.C(n_155),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_138),
.B(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_195),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_198),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_141),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_205),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_207),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_212),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_209),
.B1(n_219),
.B2(n_178),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_157),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_186),
.A2(n_130),
.B1(n_147),
.B2(n_153),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_168),
.A2(n_147),
.B(n_47),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_220),
.B(n_184),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_20),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_169),
.B(n_23),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_217),
.C(n_169),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_216),
.A2(n_180),
.B1(n_167),
.B2(n_174),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_24),
.C(n_38),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_173),
.A2(n_19),
.B1(n_11),
.B2(n_14),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_170),
.A2(n_47),
.B(n_13),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_23),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_223),
.A2(n_219),
.B1(n_12),
.B2(n_11),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_196),
.B(n_188),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_224),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_190),
.C(n_195),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_230),
.C(n_235),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_185),
.Y(n_226)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_229),
.A2(n_232),
.B1(n_209),
.B2(n_204),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_183),
.C(n_185),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_202),
.A2(n_191),
.B1(n_181),
.B2(n_187),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_171),
.Y(n_233)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_198),
.A2(n_194),
.B(n_213),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_210),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_183),
.C(n_194),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_179),
.C(n_191),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_238),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_184),
.C(n_193),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_206),
.A2(n_9),
.B(n_10),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_242),
.A2(n_20),
.B(n_14),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_199),
.B(n_38),
.C(n_25),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_38),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_251),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_215),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_252),
.Y(n_264)
);

NOR3xp33_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_218),
.C(n_216),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_258),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_241),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_254),
.B(n_261),
.Y(n_273)
);

OAI321xp33_ASAP7_75t_L g256 ( 
.A1(n_234),
.A2(n_23),
.A3(n_25),
.B1(n_8),
.B2(n_10),
.C(n_4),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_223),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_262),
.C(n_221),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_238),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_12),
.Y(n_262)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_248),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_246),
.A2(n_245),
.B(n_260),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_267),
.A2(n_270),
.B(n_271),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_225),
.C(n_228),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_269),
.C(n_274),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_236),
.C(n_235),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_250),
.A2(n_231),
.B(n_227),
.Y(n_270)
);

NOR2xp67_ASAP7_75t_SL g271 ( 
.A(n_257),
.B(n_232),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_227),
.C(n_243),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_229),
.C(n_25),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_277),
.C(n_0),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_23),
.C(n_1),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_289),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_249),
.Y(n_280)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_280),
.Y(n_301)
);

OA21x2_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_247),
.B(n_254),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_4),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_253),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_6),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_276),
.B(n_252),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_290),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_286),
.B(n_287),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

AOI21x1_ASAP7_75t_L g288 ( 
.A1(n_263),
.A2(n_265),
.B(n_6),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_10),
.Y(n_298)
);

NOR2xp67_ASAP7_75t_SL g289 ( 
.A(n_265),
.B(n_6),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_268),
.B(n_6),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_0),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_287),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_292),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_294),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_279),
.A2(n_4),
.B(n_9),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_297),
.A2(n_302),
.B1(n_7),
.B2(n_1),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_7),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_282),
.A2(n_4),
.B(n_8),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_305),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_282),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_284),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_0),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_7),
.Y(n_308)
);

O2A1O1Ixp33_ASAP7_75t_SL g312 ( 
.A1(n_309),
.A2(n_295),
.B(n_300),
.C(n_2),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_SL g314 ( 
.A1(n_311),
.A2(n_300),
.B(n_1),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_315),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_314),
.B(n_307),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_310),
.B(n_313),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_303),
.Y(n_319)
);

AOI31xp33_ASAP7_75t_SL g320 ( 
.A1(n_319),
.A2(n_316),
.A3(n_311),
.B(n_2),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_0),
.B(n_1),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_3),
.B(n_307),
.Y(n_322)
);


endmodule