module fake_jpeg_12626_n_176 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_9),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_4),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_3),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_37),
.B(n_40),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_4),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_58),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_5),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_54),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_7),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_57),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_8),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_16),
.B(n_24),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_16),
.B(n_22),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_61),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_63),
.Y(n_71)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_10),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_11),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_13),
.B(n_11),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_35),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_91),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_13),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_92),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_94),
.B1(n_81),
.B2(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_80),
.B(n_85),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_42),
.A2(n_25),
.B1(n_34),
.B2(n_23),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g83 ( 
.A1(n_37),
.A2(n_25),
.B(n_34),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_20),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_46),
.A2(n_51),
.B1(n_41),
.B2(n_49),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_96),
.B(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_20),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_75),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_40),
.A2(n_35),
.B1(n_58),
.B2(n_53),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_64),
.B1(n_60),
.B2(n_61),
.Y(n_96)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_88),
.B(n_83),
.C(n_84),
.Y(n_102)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_115),
.A3(n_121),
.B1(n_112),
.B2(n_111),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_96),
.B(n_71),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_117),
.C(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_112),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_109),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_70),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_98),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

AOI32xp33_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_96),
.A3(n_97),
.B1(n_90),
.B2(n_86),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_108),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_67),
.Y(n_113)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_79),
.Y(n_114)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_77),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_73),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_78),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_116),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_72),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_136),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_117),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_129),
.B1(n_124),
.B2(n_131),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_103),
.C(n_121),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_101),
.C(n_107),
.Y(n_147)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_135),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_106),
.B1(n_104),
.B2(n_102),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_122),
.B1(n_117),
.B2(n_110),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_115),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_139),
.B(n_141),
.Y(n_150)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_140),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_137),
.B(n_100),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_143),
.B(n_145),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_110),
.B1(n_113),
.B2(n_99),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_148),
.B1(n_127),
.B2(n_123),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_138),
.B(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_139),
.B1(n_145),
.B2(n_147),
.Y(n_160)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_149),
.Y(n_159)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_132),
.B(n_142),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_160),
.Y(n_164)
);

NOR2xp67_ASAP7_75t_R g161 ( 
.A(n_156),
.B(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_151),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_150),
.A2(n_148),
.B1(n_142),
.B2(n_138),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_162),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_167),
.B(n_160),
.Y(n_169)
);

OAI31xp33_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_166),
.A3(n_141),
.B(n_158),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_169),
.B(n_170),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_159),
.B(n_151),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_146),
.B(n_157),
.Y(n_173)
);

OAI321xp33_ASAP7_75t_L g175 ( 
.A1(n_173),
.A2(n_174),
.A3(n_153),
.B1(n_154),
.B2(n_140),
.C(n_128),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_164),
.C(n_134),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_125),
.Y(n_176)
);


endmodule