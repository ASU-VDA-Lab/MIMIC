module fake_jpeg_26222_n_143 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx10_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_35),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_0),
.C(n_1),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_30),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g38 ( 
.A(n_18),
.B(n_22),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_20),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_22),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_32),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_52),
.B1(n_16),
.B2(n_17),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_49),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_29),
.B1(n_23),
.B2(n_25),
.Y(n_45)
);

AO21x1_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_52),
.B(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_17),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_34),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_65),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_62),
.Y(n_78)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_60),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_39),
.B1(n_31),
.B2(n_27),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_67),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_31),
.B1(n_39),
.B2(n_24),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_69),
.B1(n_43),
.B2(n_15),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_70),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_39),
.B1(n_25),
.B2(n_21),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

FAx1_ASAP7_75t_SL g71 ( 
.A(n_65),
.B(n_40),
.CI(n_52),
.CON(n_71),
.SN(n_71)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_83),
.B1(n_61),
.B2(n_49),
.Y(n_91)
);

OAI32xp33_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_47),
.A3(n_21),
.B1(n_20),
.B2(n_36),
.Y(n_83)
);

XNOR2x2_ASAP7_75t_SL g84 ( 
.A(n_56),
.B(n_47),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_84),
.B(n_36),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_71),
.B1(n_46),
.B2(n_20),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_61),
.C(n_67),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_100),
.C(n_78),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_96),
.B(n_99),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_36),
.B(n_57),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_78),
.B(n_74),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_97),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_82),
.B(n_79),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_36),
.B(n_46),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_67),
.C(n_57),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_100),
.C(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_78),
.B(n_84),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_106),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_81),
.B(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_83),
.Y(n_109)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_0),
.B(n_2),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_111),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_101),
.C(n_92),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_91),
.B1(n_96),
.B2(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_112),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_108),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_120),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_123),
.A2(n_126),
.B(n_127),
.Y(n_130)
);

OA21x2_ASAP7_75t_SL g124 ( 
.A1(n_113),
.A2(n_107),
.B(n_105),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_114),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_118),
.A2(n_109),
.B(n_103),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_103),
.B(n_109),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_89),
.C(n_9),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_129),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_7),
.C(n_12),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_118),
.B(n_119),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_121),
.B(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_125),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_7),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_137),
.C(n_138),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_116),
.B1(n_13),
.B2(n_11),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_130),
.B(n_116),
.Y(n_139)
);

NOR2xp67_ASAP7_75t_SL g141 ( 
.A(n_139),
.B(n_140),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_10),
.C(n_5),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_6),
.Y(n_143)
);


endmodule