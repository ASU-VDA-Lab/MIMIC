module fake_jpeg_794_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_43;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

AOI21xp33_ASAP7_75t_L g7 ( 
.A1(n_3),
.A2(n_6),
.B(n_4),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_SL g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_2),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_10),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_18),
.Y(n_24)
);

AND2x2_ASAP7_75t_SL g17 ( 
.A(n_11),
.B(n_1),
.Y(n_17)
);

NOR3xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_21),
.C(n_22),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_8),
.Y(n_18)
);

INVxp67_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_9),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_14),
.B1(n_13),
.B2(n_7),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_28),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_19),
.B(n_16),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_23),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVxp33_ASAP7_75t_SL g37 ( 
.A(n_32),
.Y(n_37)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_25),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_41),
.B(n_42),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_38),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_38),
.C(n_37),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);


endmodule