module fake_jpeg_8524_n_295 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_37),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_0),
.C(n_1),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_21),
.C(n_24),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_44),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_57),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_18),
.B1(n_25),
.B2(n_31),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_58),
.B1(n_21),
.B2(n_22),
.Y(n_83)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_18),
.B1(n_25),
.B2(n_29),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_52),
.A2(n_47),
.B1(n_22),
.B2(n_57),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_12),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_54),
.B(n_66),
.Y(n_85)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_18),
.B1(n_25),
.B2(n_31),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_18),
.B1(n_31),
.B2(n_29),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_59),
.A2(n_65),
.B1(n_28),
.B2(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_60),
.B(n_0),
.Y(n_103)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_64),
.Y(n_102)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_31),
.B1(n_29),
.B2(n_26),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_23),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_21),
.Y(n_68)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_84),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_19),
.B1(n_35),
.B2(n_29),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_71),
.A2(n_74),
.B1(n_83),
.B2(n_64),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_26),
.B1(n_19),
.B2(n_33),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_72),
.A2(n_89),
.B1(n_90),
.B2(n_101),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_82),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_26),
.B1(n_36),
.B2(n_40),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_22),
.B(n_26),
.C(n_33),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_SL g111 ( 
.A(n_75),
.B(n_95),
.C(n_27),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_78),
.B(n_79),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_40),
.B1(n_36),
.B2(n_33),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_81),
.A2(n_56),
.B1(n_46),
.B2(n_67),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_66),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_36),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_97),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_37),
.C(n_34),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_37),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_47),
.A2(n_23),
.B1(n_32),
.B2(n_28),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_98),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_27),
.B1(n_30),
.B2(n_46),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_17),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_49),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_100),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_58),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_32),
.B1(n_28),
.B2(n_30),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_27),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_116),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_124),
.B1(n_83),
.B2(n_80),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_121),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_114),
.B(n_129),
.Y(n_162)
);

AO21x2_ASAP7_75t_L g115 ( 
.A1(n_74),
.A2(n_50),
.B(n_51),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_115),
.A2(n_119),
.B1(n_97),
.B2(n_74),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g116 ( 
.A(n_77),
.Y(n_116)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_32),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_77),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_102),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_115),
.B1(n_100),
.B2(n_89),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_30),
.B1(n_27),
.B2(n_20),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_1),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_69),
.B(n_46),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_118),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_139),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_128),
.A2(n_87),
.B(n_79),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_135),
.A2(n_55),
.B(n_127),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_137),
.A2(n_140),
.B1(n_156),
.B2(n_30),
.Y(n_186)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_138),
.B(n_143),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_103),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_85),
.B(n_82),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_161),
.B(n_34),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_142),
.B(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_88),
.B1(n_78),
.B2(n_85),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_153),
.B1(n_160),
.B2(n_126),
.Y(n_168)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_95),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_155),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_110),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_154),
.Y(n_181)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_125),
.B(n_95),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_74),
.B1(n_102),
.B2(n_71),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_112),
.B(n_86),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_91),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_86),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_98),
.B1(n_71),
.B2(n_81),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_111),
.A2(n_71),
.B(n_34),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_133),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_172),
.C(n_188),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_166),
.B(n_20),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_168),
.A2(n_170),
.B1(n_185),
.B2(n_192),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_105),
.B1(n_129),
.B2(n_122),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_114),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_177),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_176),
.B(n_178),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_132),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g178 ( 
.A1(n_151),
.A2(n_120),
.B(n_127),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_184),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_131),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_131),
.Y(n_183)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_135),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_152),
.A2(n_110),
.B1(n_20),
.B2(n_17),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_167),
.B1(n_181),
.B2(n_179),
.Y(n_214)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_189),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_141),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_190),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_20),
.B1(n_17),
.B2(n_30),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_188),
.B(n_148),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_180),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_155),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_199),
.C(n_201),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_195),
.B(n_165),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_151),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_161),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_151),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_204),
.C(n_216),
.Y(n_231)
);

OAI22x1_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_137),
.B1(n_156),
.B2(n_160),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_203),
.A2(n_210),
.B(n_175),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_140),
.Y(n_204)
);

AOI322xp5_ASAP7_75t_L g209 ( 
.A1(n_170),
.A2(n_147),
.A3(n_138),
.B1(n_142),
.B2(n_143),
.C1(n_136),
.C2(n_157),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_191),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_34),
.B(n_2),
.Y(n_210)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_214),
.A2(n_215),
.B1(n_8),
.B2(n_15),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_168),
.A2(n_20),
.B1(n_17),
.B2(n_3),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_163),
.B(n_182),
.C(n_189),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_163),
.C(n_177),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_218),
.B(n_223),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_173),
.Y(n_219)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_204),
.Y(n_249)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_227),
.Y(n_246)
);

XOR2x2_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_191),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_236),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_165),
.B1(n_185),
.B2(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_187),
.Y(n_226)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_232),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_229),
.B(n_233),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_210),
.B(n_200),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_215),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_205),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_214),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_211),
.B(n_175),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_234),
.B(n_227),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_197),
.B1(n_9),
.B2(n_16),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_8),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_194),
.C(n_199),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_238),
.C(n_239),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_193),
.C(n_201),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_202),
.C(n_208),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_224),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_249),
.B(n_220),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_207),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_1),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_217),
.B(n_198),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_198),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_223),
.B1(n_222),
.B2(n_235),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_255),
.B1(n_257),
.B2(n_264),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_246),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_259),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_240),
.A2(n_229),
.B1(n_225),
.B2(n_230),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_265),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_243),
.A2(n_218),
.B1(n_219),
.B2(n_217),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_16),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_262),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_247),
.A2(n_245),
.B(n_241),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_236),
.C(n_2),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_242),
.C(n_249),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_241),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_250),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_268),
.C(n_275),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_263),
.A2(n_238),
.B(n_237),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_7),
.B(n_13),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_242),
.C(n_10),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_268),
.C(n_272),
.Y(n_283)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_274),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_8),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_275),
.B(n_257),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_277),
.B(n_280),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_273),
.A2(n_255),
.B(n_259),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_266),
.B(n_253),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_256),
.C(n_10),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_281),
.A2(n_282),
.B(n_283),
.Y(n_288)
);

AOI21x1_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_270),
.B(n_271),
.Y(n_284)
);

NAND2xp33_ASAP7_75t_SL g290 ( 
.A(n_284),
.B(n_285),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_279),
.A2(n_272),
.B1(n_7),
.B2(n_5),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_14),
.B1(n_5),
.B2(n_6),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_286),
.C(n_13),
.Y(n_291)
);

NOR4xp25_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_5),
.C(n_6),
.D(n_11),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_289),
.A2(n_13),
.B(n_14),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_291),
.A2(n_3),
.B1(n_4),
.B2(n_290),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_292),
.B(n_293),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_4),
.Y(n_295)
);


endmodule