module fake_jpeg_20799_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

INVx8_ASAP7_75t_SL g10 ( 
.A(n_1),
.Y(n_10)
);

INVx13_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_11),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_9),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_13),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_25),
.B1(n_24),
.B2(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_41),
.Y(n_44)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

OAI21x1_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_21),
.B(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_39),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_23),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_16),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_41),
.C(n_34),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_34),
.C(n_25),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_53),
.C(n_55),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_42),
.C(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_56),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_23),
.C(n_20),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_15),
.C(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_14),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_44),
.B1(n_49),
.B2(n_16),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_61),
.B1(n_12),
.B2(n_4),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_15),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_44),
.B1(n_14),
.B2(n_9),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_46),
.B1(n_19),
.B2(n_12),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_64),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_67),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_58),
.B(n_6),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_40),
.Y(n_69)
);

OAI321xp33_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_68),
.A3(n_39),
.B1(n_8),
.B2(n_2),
.C(n_33),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_70),
.Y(n_72)
);


endmodule