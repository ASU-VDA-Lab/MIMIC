module real_aes_14805_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_905;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_919;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_656;
wire n_153;
wire n_316;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx2_ASAP7_75t_SL g681 ( .A(n_0), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_1), .Y(n_570) );
INVx1_ASAP7_75t_L g143 ( .A(n_2), .Y(n_143) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_2), .A2(n_46), .B(n_145), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_3), .B(n_256), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_4), .B(n_252), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_5), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_6), .B(n_211), .Y(n_210) );
NAND2xp33_ASAP7_75t_L g235 ( .A(n_7), .B(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g661 ( .A(n_8), .B(n_239), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_9), .A2(n_89), .B1(n_912), .B2(n_913), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_9), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_10), .B(n_270), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_11), .B(n_159), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_12), .B(n_184), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_13), .Y(n_140) );
BUFx3_ASAP7_75t_L g161 ( .A(n_14), .Y(n_161) );
INVx1_ASAP7_75t_L g178 ( .A(n_14), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_15), .B(n_238), .Y(n_638) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_16), .A2(n_192), .B(n_193), .C(n_195), .Y(n_191) );
BUFx10_ASAP7_75t_L g542 ( .A(n_17), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_18), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_19), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_20), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_21), .B(n_258), .Y(n_315) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_22), .A2(n_175), .B(n_179), .C(n_182), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_23), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g696 ( .A(n_24), .B(n_280), .C(n_694), .Y(n_696) );
AND2x2_ASAP7_75t_L g248 ( .A(n_25), .B(n_247), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_26), .B(n_211), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_27), .B(n_238), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g166 ( .A1(n_28), .A2(n_70), .B1(n_162), .B2(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g151 ( .A(n_29), .Y(n_151) );
INVx1_ASAP7_75t_L g215 ( .A(n_30), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_31), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_32), .B(n_162), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_33), .B(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g112 ( .A(n_34), .Y(n_112) );
AND3x2_ASAP7_75t_L g919 ( .A(n_34), .B(n_104), .C(n_547), .Y(n_919) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_35), .B(n_176), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_36), .B(n_192), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_37), .B(n_238), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_38), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_39), .B(n_200), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_40), .Y(n_194) );
AND2x4_ASAP7_75t_L g150 ( .A(n_41), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_42), .B(n_238), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_43), .B(n_247), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_44), .B(n_238), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g158 ( .A1(n_45), .A2(n_83), .B1(n_159), .B2(n_162), .Y(n_158) );
INVx1_ASAP7_75t_L g142 ( .A(n_46), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g655 ( .A(n_47), .Y(n_655) );
A2O1A1Ixp33_ASAP7_75t_L g679 ( .A1(n_48), .A2(n_656), .B(n_680), .C(n_682), .Y(n_679) );
INVx1_ASAP7_75t_L g145 ( .A(n_49), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_50), .B(n_238), .Y(n_575) );
AND2x4_ASAP7_75t_L g109 ( .A(n_51), .B(n_110), .Y(n_109) );
OAI22xp33_ASAP7_75t_L g129 ( .A1(n_52), .A2(n_97), .B1(n_130), .B2(n_131), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_52), .Y(n_131) );
INVx3_ASAP7_75t_L g622 ( .A(n_53), .Y(n_622) );
NOR2xp67_ASAP7_75t_L g105 ( .A(n_54), .B(n_72), .Y(n_105) );
AND2x2_ASAP7_75t_L g322 ( .A(n_55), .B(n_239), .Y(n_322) );
INVx1_ASAP7_75t_L g110 ( .A(n_56), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_57), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_58), .B(n_598), .Y(n_603) );
NAND2x1_ASAP7_75t_L g285 ( .A(n_59), .B(n_192), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_60), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g634 ( .A(n_61), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_62), .B(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_63), .B(n_268), .Y(n_267) );
AND3x2_ASAP7_75t_L g103 ( .A(n_64), .B(n_104), .C(n_106), .Y(n_103) );
INVx2_ASAP7_75t_L g122 ( .A(n_64), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_65), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_66), .B(n_159), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_67), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_68), .B(n_280), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_69), .B(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_71), .B(n_176), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_73), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_74), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_75), .B(n_270), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g916 ( .A(n_76), .Y(n_916) );
NAND2xp33_ASAP7_75t_SL g208 ( .A(n_77), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_78), .B(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g674 ( .A(n_79), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_80), .B(n_203), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g657 ( .A(n_81), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_82), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g155 ( .A(n_84), .Y(n_155) );
BUFx3_ASAP7_75t_L g184 ( .A(n_84), .Y(n_184) );
INVx1_ASAP7_75t_L g206 ( .A(n_84), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_85), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_86), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_87), .B(n_159), .Y(n_568) );
INVx1_ASAP7_75t_L g620 ( .A(n_88), .Y(n_620) );
INVx1_ASAP7_75t_L g913 ( .A(n_89), .Y(n_913) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_90), .B(n_268), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_91), .B(n_239), .Y(n_588) );
NAND2xp33_ASAP7_75t_L g229 ( .A(n_92), .B(n_230), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g921 ( .A(n_93), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_94), .B(n_602), .Y(n_601) );
CKINVDCx5p33_ASAP7_75t_R g616 ( .A(n_95), .Y(n_616) );
INVx1_ASAP7_75t_L g612 ( .A(n_96), .Y(n_612) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_97), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g651 ( .A(n_98), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_99), .B(n_200), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_100), .B(n_598), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_113), .B(n_920), .Y(n_101) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
BUFx6f_ASAP7_75t_L g923 ( .A(n_103), .Y(n_923) );
AND2x2_ASAP7_75t_L g546 ( .A(n_104), .B(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_105), .B(n_112), .Y(n_123) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_111), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g554 ( .A(n_111), .Y(n_554) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_124), .Y(n_113) );
NOR2xp67_ASAP7_75t_L g125 ( .A(n_114), .B(n_126), .Y(n_125) );
NOR2xp67_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g537 ( .A(n_119), .Y(n_537) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NOR2x1p5_ASAP7_75t_L g120 ( .A(n_121), .B(n_123), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g547 ( .A(n_122), .Y(n_547) );
OAI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_538), .B(n_543), .Y(n_124) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_536), .Y(n_127) );
XNOR2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_132), .Y(n_128) );
AOI22x1_ASAP7_75t_L g550 ( .A1(n_132), .A2(n_551), .B1(n_555), .B2(n_909), .Y(n_550) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_440), .Y(n_132) );
NOR3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_349), .C(n_413), .Y(n_133) );
OAI221xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_241), .B1(n_288), .B2(n_299), .C(n_304), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_169), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g361 ( .A(n_137), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g376 ( .A(n_137), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g449 ( .A(n_137), .B(n_196), .Y(n_449) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g296 ( .A(n_138), .Y(n_296) );
INVx1_ASAP7_75t_L g328 ( .A(n_138), .Y(n_328) );
AND2x2_ASAP7_75t_L g347 ( .A(n_138), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g374 ( .A(n_138), .B(n_364), .Y(n_374) );
INVxp67_ASAP7_75t_L g389 ( .A(n_138), .Y(n_389) );
AND2x2_ASAP7_75t_L g412 ( .A(n_138), .B(n_223), .Y(n_412) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_138), .Y(n_439) );
OR2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_146), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_141), .B(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g189 ( .A(n_141), .Y(n_189) );
AO21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_144), .Y(n_141) );
AOI21x1_ASAP7_75t_L g157 ( .A1(n_142), .A2(n_143), .B(n_144), .Y(n_157) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_158), .B1(n_164), .B2(n_166), .Y(n_146) );
NAND3xp33_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .C(n_156), .Y(n_147) );
NAND3xp33_ASAP7_75t_L g164 ( .A(n_148), .B(n_156), .C(n_165), .Y(n_164) );
BUFx2_ASAP7_75t_L g660 ( .A(n_148), .Y(n_660) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OAI21xp33_ASAP7_75t_L g683 ( .A1(n_149), .A2(n_189), .B(n_678), .Y(n_683) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g187 ( .A(n_150), .Y(n_187) );
BUFx6f_ASAP7_75t_SL g221 ( .A(n_150), .Y(n_221) );
INVx1_ASAP7_75t_L g312 ( .A(n_150), .Y(n_312) );
INVx3_ASAP7_75t_L g614 ( .A(n_150), .Y(n_614) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_153), .B(n_614), .Y(n_617) );
NOR3xp33_ASAP7_75t_L g621 ( .A(n_153), .B(n_614), .C(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g195 ( .A(n_154), .Y(n_195) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx3_ASAP7_75t_L g165 ( .A(n_155), .Y(n_165) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_156), .Y(n_608) );
NOR2xp33_ASAP7_75t_SL g623 ( .A(n_156), .B(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g211 ( .A(n_160), .Y(n_211) );
INVx2_ASAP7_75t_L g234 ( .A(n_160), .Y(n_234) );
INVx2_ASAP7_75t_L g258 ( .A(n_160), .Y(n_258) );
INVx2_ASAP7_75t_L g572 ( .A(n_160), .Y(n_572) );
INVx3_ASAP7_75t_L g648 ( .A(n_160), .Y(n_648) );
INVx3_ASAP7_75t_L g673 ( .A(n_160), .Y(n_673) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g163 ( .A(n_161), .Y(n_163) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_161), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_162), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g236 ( .A(n_163), .Y(n_236) );
INVx1_ASAP7_75t_L g280 ( .A(n_163), .Y(n_280) );
O2A1O1Ixp5_ASAP7_75t_L g282 ( .A1(n_165), .A2(n_283), .B(n_284), .C(n_285), .Y(n_282) );
INVx2_ASAP7_75t_L g316 ( .A(n_165), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_165), .A2(n_582), .B(n_583), .Y(n_581) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g203 ( .A(n_168), .Y(n_203) );
INVx2_ASAP7_75t_L g228 ( .A(n_168), .Y(n_228) );
INVx2_ASAP7_75t_L g320 ( .A(n_168), .Y(n_320) );
OAI21xp33_ASAP7_75t_L g417 ( .A1(n_169), .A2(n_418), .B(n_422), .Y(n_417) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_196), .Y(n_169) );
AND2x2_ASAP7_75t_L g519 ( .A(n_170), .B(n_412), .Y(n_519) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
BUFx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g292 ( .A(n_172), .Y(n_292) );
INVx1_ASAP7_75t_L g330 ( .A(n_172), .Y(n_330) );
AND2x2_ASAP7_75t_L g358 ( .A(n_172), .B(n_295), .Y(n_358) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_172), .Y(n_387) );
NAND2x1p5_ASAP7_75t_L g172 ( .A(n_173), .B(n_190), .Y(n_172) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_173), .B(n_190), .Y(n_348) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_185), .B(n_188), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_175), .A2(n_598), .B1(n_619), .B2(n_621), .Y(n_618) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_176), .B(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g587 ( .A(n_176), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_176), .B(n_612), .Y(n_611) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx3_ASAP7_75t_L g181 ( .A(n_177), .Y(n_181) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_178), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
INVx2_ASAP7_75t_L g192 ( .A(n_181), .Y(n_192) );
INVx2_ASAP7_75t_L g252 ( .A(n_181), .Y(n_252) );
INVx2_ASAP7_75t_L g268 ( .A(n_181), .Y(n_268) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_181), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_182), .A2(n_233), .B(n_235), .Y(n_232) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_183), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g212 ( .A(n_184), .Y(n_212) );
INVx1_ASAP7_75t_L g231 ( .A(n_184), .Y(n_231) );
AOI211x1_ASAP7_75t_L g249 ( .A1(n_184), .A2(n_248), .B(n_250), .C(n_254), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_184), .B(n_614), .Y(n_613) );
NOR3xp33_ASAP7_75t_L g619 ( .A(n_184), .B(n_614), .C(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g190 ( .A(n_185), .B(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g605 ( .A(n_186), .Y(n_605) );
INVx2_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g286 ( .A(n_187), .Y(n_286) );
INVx1_ASAP7_75t_L g574 ( .A(n_187), .Y(n_574) );
INVxp67_ASAP7_75t_L g659 ( .A(n_189), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_195), .A2(n_597), .B(n_599), .Y(n_596) );
INVx1_ASAP7_75t_L g658 ( .A(n_195), .Y(n_658) );
AND2x2_ASAP7_75t_L g346 ( .A(n_196), .B(n_347), .Y(n_346) );
INVx3_ASAP7_75t_L g535 ( .A(n_196), .Y(n_535) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_222), .Y(n_196) );
INVx2_ASAP7_75t_L g295 ( .A(n_197), .Y(n_295) );
AND2x2_ASAP7_75t_L g329 ( .A(n_197), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g340 ( .A(n_197), .Y(n_340) );
OR2x2_ASAP7_75t_L g378 ( .A(n_197), .B(n_348), .Y(n_378) );
AND2x2_ASAP7_75t_L g390 ( .A(n_197), .B(n_348), .Y(n_390) );
AND2x2_ASAP7_75t_L g460 ( .A(n_197), .B(n_223), .Y(n_460) );
AO31x2_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_207), .A3(n_213), .B(n_218), .Y(n_197) );
AO21x1_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_202), .B(n_204), .Y(n_198) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g209 ( .A(n_201), .Y(n_209) );
INVx1_ASAP7_75t_L g230 ( .A(n_201), .Y(n_230) );
INVx2_ASAP7_75t_L g256 ( .A(n_201), .Y(n_256) );
INVx2_ASAP7_75t_L g284 ( .A(n_203), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_204), .A2(n_255), .B(n_257), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_204), .A2(n_267), .B(n_269), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_204), .A2(n_279), .B(n_281), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_204), .A2(n_567), .B(n_568), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_204), .A2(n_585), .B(n_586), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_204), .A2(n_636), .B(n_637), .Y(n_635) );
BUFx10_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g694 ( .A(n_205), .Y(n_694) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
BUFx3_ASAP7_75t_L g652 ( .A(n_206), .Y(n_652) );
AO21x1_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_210), .B(n_212), .Y(n_207) );
INVx2_ASAP7_75t_L g270 ( .A(n_209), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_212), .A2(n_264), .B(n_265), .Y(n_263) );
O2A1O1Ixp5_ASAP7_75t_L g569 ( .A1(n_212), .A2(n_570), .B(n_571), .C(n_573), .Y(n_569) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_214), .A2(n_219), .B(n_221), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
INVxp33_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
BUFx2_ASAP7_75t_L g220 ( .A(n_217), .Y(n_220) );
INVx1_ASAP7_75t_L g240 ( .A(n_217), .Y(n_240) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_217), .Y(n_247) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
BUFx3_ASAP7_75t_L g224 ( .A(n_220), .Y(n_224) );
OAI21x1_ASAP7_75t_L g225 ( .A1(n_221), .A2(n_226), .B(n_232), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_221), .A2(n_246), .B(n_248), .Y(n_245) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_221), .A2(n_263), .B(n_266), .Y(n_262) );
OAI21x1_ASAP7_75t_L g580 ( .A1(n_221), .A2(n_581), .B(n_584), .Y(n_580) );
OAI21x1_ASAP7_75t_L g628 ( .A1(n_221), .A2(n_629), .B(n_635), .Y(n_628) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g298 ( .A(n_223), .Y(n_298) );
INVx1_ASAP7_75t_L g364 ( .A(n_223), .Y(n_364) );
AND2x2_ASAP7_75t_L g386 ( .A(n_223), .B(n_296), .Y(n_386) );
AND2x2_ASAP7_75t_L g469 ( .A(n_223), .B(n_363), .Y(n_469) );
OAI21x1_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_237), .Y(n_223) );
OAI21x1_ASAP7_75t_L g564 ( .A1(n_224), .A2(n_565), .B(n_575), .Y(n_564) );
OAI21x1_ASAP7_75t_L g627 ( .A1(n_224), .A2(n_628), .B(n_638), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_229), .B(n_231), .Y(n_226) );
INVx2_ASAP7_75t_L g598 ( .A(n_228), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_228), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g602 ( .A(n_230), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_231), .A2(n_319), .B(n_321), .Y(n_318) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_238), .Y(n_687) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_259), .Y(n_241) );
AND2x2_ASAP7_75t_L g392 ( .A(n_242), .B(n_383), .Y(n_392) );
OR2x2_ASAP7_75t_L g408 ( .A(n_242), .B(n_343), .Y(n_408) );
INVx2_ASAP7_75t_L g420 ( .A(n_242), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_242), .B(n_356), .Y(n_423) );
AND2x2_ASAP7_75t_L g520 ( .A(n_242), .B(n_435), .Y(n_520) );
BUFx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g300 ( .A(n_243), .B(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g430 ( .A(n_243), .B(n_335), .Y(n_430) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g323 ( .A(n_244), .B(n_261), .Y(n_323) );
INVx2_ASAP7_75t_L g354 ( .A(n_244), .Y(n_354) );
BUFx2_ASAP7_75t_L g381 ( .A(n_244), .Y(n_381) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_244), .Y(n_398) );
INVx1_ASAP7_75t_L g405 ( .A(n_244), .Y(n_405) );
AND2x2_ASAP7_75t_L g464 ( .A(n_244), .B(n_407), .Y(n_464) );
INVx1_ASAP7_75t_L g525 ( .A(n_244), .Y(n_525) );
OR2x6_ASAP7_75t_L g244 ( .A(n_245), .B(n_249), .Y(n_244) );
INVxp67_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_247), .Y(n_272) );
NOR2xp67_ASAP7_75t_SL g311 ( .A(n_247), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g732 ( .A(n_247), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_253), .Y(n_250) );
INVx2_ASAP7_75t_L g656 ( .A(n_256), .Y(n_656) );
INVxp67_ASAP7_75t_L g630 ( .A(n_258), .Y(n_630) );
INVxp67_ASAP7_75t_L g654 ( .A(n_258), .Y(n_654) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_274), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_260), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g334 ( .A(n_261), .B(n_335), .Y(n_334) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_271), .B(n_273), .Y(n_261) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_262), .A2(n_271), .B(n_273), .Y(n_303) );
INVx2_ASAP7_75t_L g650 ( .A(n_268), .Y(n_650) );
OAI21x1_ASAP7_75t_L g276 ( .A1(n_271), .A2(n_277), .B(n_287), .Y(n_276) );
OAI21x1_ASAP7_75t_L g579 ( .A1(n_271), .A2(n_580), .B(n_588), .Y(n_579) );
OAI21x1_ASAP7_75t_L g716 ( .A1(n_271), .A2(n_645), .B(n_717), .Y(n_716) );
OAI21x1_ASAP7_75t_L g722 ( .A1(n_271), .A2(n_580), .B(n_588), .Y(n_722) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2x1_ASAP7_75t_SL g604 ( .A(n_272), .B(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g490 ( .A(n_274), .Y(n_490) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g407 ( .A(n_275), .Y(n_407) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g333 ( .A(n_276), .Y(n_333) );
INVx1_ASAP7_75t_L g370 ( .A(n_276), .Y(n_370) );
OAI21xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_282), .B(n_286), .Y(n_277) );
OAI211xp5_ASAP7_75t_L g413 ( .A1(n_288), .A2(n_414), .B(n_417), .C(n_424), .Y(n_413) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2x1p5_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_292), .Y(n_337) );
AND2x2_ASAP7_75t_L g456 ( .A(n_292), .B(n_386), .Y(n_456) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
AND2x2_ASAP7_75t_L g366 ( .A(n_294), .B(n_362), .Y(n_366) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g427 ( .A(n_295), .Y(n_427) );
INVx2_ASAP7_75t_L g400 ( .A(n_297), .Y(n_400) );
BUFx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_298), .B(n_340), .Y(n_339) );
INVxp67_ASAP7_75t_SL g502 ( .A(n_298), .Y(n_502) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g356 ( .A(n_301), .B(n_333), .Y(n_356) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g369 ( .A(n_302), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g383 ( .A(n_302), .B(n_309), .Y(n_383) );
AND2x2_ASAP7_75t_L g506 ( .A(n_302), .B(n_333), .Y(n_506) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g344 ( .A(n_303), .B(n_309), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_324), .B1(n_331), .B2(n_336), .C(n_341), .Y(n_304) );
AOI222xp33_ASAP7_75t_L g498 ( .A1(n_305), .A2(n_436), .B1(n_499), .B2(n_504), .C1(n_507), .C2(n_508), .Y(n_498) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2x1_ASAP7_75t_L g306 ( .A(n_307), .B(n_323), .Y(n_306) );
INVx4_ASAP7_75t_R g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_308), .B(n_399), .Y(n_416) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g335 ( .A(n_309), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_309), .B(n_333), .Y(n_343) );
AND2x4_ASAP7_75t_L g404 ( .A(n_309), .B(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_317), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_311), .A2(n_318), .B(n_322), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B(n_316), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_316), .A2(n_601), .B(n_603), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_320), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g359 ( .A(n_323), .Y(n_359) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_329), .Y(n_325) );
NAND3xp33_ASAP7_75t_L g511 ( .A(n_326), .B(n_512), .C(n_515), .Y(n_511) );
OR2x2_ASAP7_75t_L g527 ( .A(n_326), .B(n_515), .Y(n_527) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI21xp33_ASAP7_75t_L g472 ( .A1(n_327), .A2(n_397), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g461 ( .A(n_328), .B(n_348), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_329), .B(n_412), .Y(n_432) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
OR2x2_ASAP7_75t_L g475 ( .A(n_332), .B(n_344), .Y(n_475) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g453 ( .A(n_334), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_334), .B(n_380), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_334), .B(n_464), .Y(n_463) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_334), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_334), .B(n_490), .Y(n_518) );
AND2x4_ASAP7_75t_SL g353 ( .A(n_335), .B(n_354), .Y(n_353) );
NOR2x1p5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
BUFx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g411 ( .A(n_340), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_340), .B(n_502), .Y(n_501) );
AOI21xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_344), .B(n_345), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx4_ASAP7_75t_L g435 ( .A(n_344), .Y(n_435) );
NOR2x1_ASAP7_75t_L g532 ( .A(n_344), .B(n_524), .Y(n_532) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g467 ( .A(n_347), .B(n_460), .Y(n_467) );
INVx2_ASAP7_75t_L g363 ( .A(n_348), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_350), .B(n_393), .Y(n_349) );
NOR3xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_371), .C(n_384), .Y(n_350) );
OAI322xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_355), .A3(n_357), .B1(n_359), .B2(n_360), .C1(n_365), .C2(n_367), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g491 ( .A(n_353), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_355), .A2(n_466), .B1(n_468), .B2(n_470), .Y(n_465) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_356), .B(n_404), .Y(n_509) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_SL g373 ( .A(n_358), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g454 ( .A(n_358), .B(n_412), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_358), .B(n_389), .Y(n_530) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g486 ( .A(n_361), .B(n_427), .Y(n_486) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI322xp5_ASAP7_75t_L g424 ( .A1(n_367), .A2(n_404), .A3(n_425), .B1(n_428), .B2(n_431), .C1(n_433), .C2(n_436), .Y(n_424) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp33_ASAP7_75t_L g429 ( .A(n_368), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g421 ( .A(n_369), .Y(n_421) );
OR2x2_ASAP7_75t_L g444 ( .A(n_369), .B(n_430), .Y(n_444) );
BUFx2_ASAP7_75t_L g399 ( .A(n_370), .Y(n_399) );
AOI21xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_375), .B(n_379), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_372), .A2(n_402), .B1(n_408), .B2(n_409), .Y(n_401) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g494 ( .A(n_374), .Y(n_494) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g397 ( .A(n_378), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g437 ( .A(n_378), .B(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g477 ( .A(n_378), .B(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g493 ( .A(n_378), .B(n_494), .Y(n_493) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_381), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g452 ( .A(n_381), .Y(n_452) );
OR2x2_ASAP7_75t_L g470 ( .A(n_382), .B(n_406), .Y(n_470) );
OR2x2_ASAP7_75t_L g496 ( .A(n_382), .B(n_490), .Y(n_496) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI21xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_388), .B(n_391), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_386), .B(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx2_ASAP7_75t_L g515 ( .A(n_390), .Y(n_515) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_400), .B(n_401), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_399), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_404), .B(n_506), .Y(n_505) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_405), .Y(n_481) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g524 ( .A(n_407), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_409), .B(n_493), .Y(n_492) );
INVx2_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx1_ASAP7_75t_L g447 ( .A(n_411), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_412), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g478 ( .A(n_412), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_414), .B(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g497 ( .A(n_420), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_420), .B(n_435), .C(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g534 ( .A(n_438), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NOR3xp33_ASAP7_75t_SL g440 ( .A(n_441), .B(n_482), .C(n_510), .Y(n_440) );
NAND3xp33_ASAP7_75t_SL g441 ( .A(n_442), .B(n_455), .C(n_471), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_445), .B1(n_450), .B2(n_454), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_449), .A2(n_517), .B1(n_519), .B2(n_520), .Y(n_516) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B1(n_459), .B2(n_462), .C(n_465), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g473 ( .A(n_459), .Y(n_473) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
INVx2_ASAP7_75t_L g503 ( .A(n_461), .Y(n_503) );
INVxp67_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVxp33_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g531 ( .A(n_470), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_474), .B1(n_476), .B2(n_479), .Y(n_471) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OAI211xp5_ASAP7_75t_SL g482 ( .A1(n_483), .A2(n_485), .B(n_487), .C(n_498), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_486), .A2(n_488), .B1(n_492), .B2(n_495), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g514 ( .A(n_490), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .Y(n_500) );
INVxp67_ASAP7_75t_SL g507 ( .A(n_501), .Y(n_507) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVxp67_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
NAND4xp25_ASAP7_75t_L g510 ( .A(n_511), .B(n_516), .C(n_521), .D(n_528), .Y(n_510) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_526), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVxp67_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_531), .B1(n_532), .B2(n_533), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx12f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OR2x6_ASAP7_75t_L g545 ( .A(n_541), .B(n_546), .Y(n_545) );
INVx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_542), .B(n_919), .Y(n_918) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_548), .B(n_915), .Y(n_543) );
CKINVDCx6p67_ASAP7_75t_R g544 ( .A(n_545), .Y(n_544) );
OAI22xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .B1(n_911), .B2(n_914), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx8_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
CKINVDCx10_ASAP7_75t_R g910 ( .A(n_553), .Y(n_910) );
BUFx6f_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_835), .Y(n_555) );
NOR3xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_770), .C(n_796), .Y(n_556) );
NAND4xp25_ASAP7_75t_SL g557 ( .A(n_558), .B(n_639), .C(n_726), .D(n_750), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_576), .Y(n_558) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g898 ( .A(n_560), .Y(n_898) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_561), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g641 ( .A(n_562), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g803 ( .A(n_562), .B(n_712), .Y(n_803) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g709 ( .A(n_563), .B(n_710), .Y(n_709) );
INVx3_ASAP7_75t_L g718 ( .A(n_563), .Y(n_718) );
AND2x2_ASAP7_75t_L g827 ( .A(n_563), .B(n_716), .Y(n_827) );
INVx2_ASAP7_75t_L g874 ( .A(n_563), .Y(n_874) );
INVx3_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OAI21xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_569), .B(n_574), .Y(n_565) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OAI21x1_ASAP7_75t_L g688 ( .A1(n_574), .A2(n_689), .B(n_692), .Y(n_688) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_589), .Y(n_576) );
OR2x2_ASAP7_75t_L g843 ( .A(n_577), .B(n_668), .Y(n_843) );
AND2x2_ASAP7_75t_L g855 ( .A(n_577), .B(n_856), .Y(n_855) );
BUFx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g740 ( .A(n_578), .Y(n_740) );
AND2x2_ASAP7_75t_L g794 ( .A(n_578), .B(n_723), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_578), .B(n_812), .Y(n_811) );
AND2x4_ASAP7_75t_L g897 ( .A(n_578), .B(n_779), .Y(n_897) );
AND2x2_ASAP7_75t_L g904 ( .A(n_578), .B(n_591), .Y(n_904) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
HB1xp67_ASAP7_75t_L g891 ( .A(n_579), .Y(n_891) );
INVxp67_ASAP7_75t_L g695 ( .A(n_587), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g837 ( .A1(n_589), .A2(n_783), .B(n_838), .C(n_839), .Y(n_837) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_606), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_590), .B(n_808), .Y(n_819) );
OR2x2_ASAP7_75t_L g834 ( .A(n_590), .B(n_811), .Y(n_834) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_590), .Y(n_846) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx2_ASAP7_75t_L g782 ( .A(n_591), .Y(n_782) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g667 ( .A(n_592), .Y(n_667) );
BUFx2_ASAP7_75t_L g700 ( .A(n_592), .Y(n_700) );
OR2x2_ASAP7_75t_L g724 ( .A(n_592), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g729 ( .A(n_592), .B(n_730), .Y(n_729) );
AND2x4_ASAP7_75t_L g829 ( .A(n_592), .B(n_749), .Y(n_829) );
INVx1_ASAP7_75t_L g886 ( .A(n_592), .Y(n_886) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2x1_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
OAI21x1_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_600), .B(n_604), .Y(n_595) );
AND2x2_ASAP7_75t_L g701 ( .A(n_606), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g795 ( .A(n_606), .B(n_788), .Y(n_795) );
AND2x2_ASAP7_75t_L g826 ( .A(n_606), .B(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g860 ( .A(n_606), .Y(n_860) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_625), .Y(n_606) );
INVx1_ASAP7_75t_L g710 ( .A(n_607), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_607), .B(n_872), .Y(n_871) );
AO21x1_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B(n_623), .Y(n_607) );
AO21x2_ASAP7_75t_L g714 ( .A1(n_608), .A2(n_609), .B(n_623), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_618), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_613), .B1(n_615), .B2(n_617), .Y(n_610) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx3_ASAP7_75t_L g664 ( .A(n_626), .Y(n_664) );
AND2x2_ASAP7_75t_L g737 ( .A(n_626), .B(n_714), .Y(n_737) );
INVx1_ASAP7_75t_L g746 ( .A(n_626), .Y(n_746) );
INVx1_ASAP7_75t_L g752 ( .A(n_626), .Y(n_752) );
AND2x2_ASAP7_75t_L g764 ( .A(n_626), .B(n_713), .Y(n_764) );
AND2x2_ASAP7_75t_L g799 ( .A(n_626), .B(n_716), .Y(n_799) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_626), .Y(n_818) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B(n_632), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_665), .B1(n_698), .B2(n_701), .C(n_705), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_662), .Y(n_640) );
AND2x2_ASAP7_75t_L g751 ( .A(n_641), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g768 ( .A(n_643), .B(n_718), .Y(n_768) );
OR2x2_ASAP7_75t_L g785 ( .A(n_643), .B(n_664), .Y(n_785) );
AO31x2_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_659), .A3(n_660), .B(n_661), .Y(n_643) );
AO31x2_ASAP7_75t_L g704 ( .A1(n_644), .A2(n_659), .A3(n_660), .B(n_661), .Y(n_704) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI22x1_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_652), .B1(n_653), .B2(n_658), .Y(n_645) );
OAI22x1_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B1(n_650), .B2(n_651), .Y(n_646) );
INVxp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g682 ( .A(n_652), .Y(n_682) );
AOI21x1_ASAP7_75t_L g689 ( .A1(n_652), .A2(n_690), .B(n_691), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_653) );
AOI21x1_ASAP7_75t_SL g671 ( .A1(n_658), .A2(n_672), .B(n_675), .Y(n_671) );
INVx1_ASAP7_75t_L g717 ( .A(n_661), .Y(n_717) );
BUFx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g833 ( .A(n_663), .B(n_815), .Y(n_833) );
NOR2xp67_ASAP7_75t_L g873 ( .A(n_663), .B(n_874), .Y(n_873) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI22xp33_ASAP7_75t_L g762 ( .A1(n_666), .A2(n_763), .B1(n_765), .B2(n_769), .Y(n_762) );
OR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_667), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g754 ( .A(n_667), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_667), .B(n_758), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_667), .B(n_791), .Y(n_790) );
NOR2xp67_ASAP7_75t_R g857 ( .A(n_667), .B(n_858), .Y(n_857) );
OR2x2_ASAP7_75t_L g699 ( .A(n_668), .B(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g739 ( .A(n_668), .B(n_740), .Y(n_739) );
OR2x6_ASAP7_75t_L g668 ( .A(n_669), .B(n_684), .Y(n_668) );
INVx2_ASAP7_75t_L g779 ( .A(n_669), .Y(n_779) );
OR2x2_ASAP7_75t_SL g809 ( .A(n_669), .B(n_730), .Y(n_809) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g723 ( .A(n_670), .Y(n_723) );
OAI21x1_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_677), .B(n_683), .Y(n_670) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
AND2x2_ASAP7_75t_L g757 ( .A(n_684), .B(n_722), .Y(n_757) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVxp67_ASAP7_75t_SL g725 ( .A(n_685), .Y(n_725) );
INVx2_ASAP7_75t_L g749 ( .A(n_685), .Y(n_749) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI21x1_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_688), .B(n_697), .Y(n_686) );
OA21x2_ASAP7_75t_L g730 ( .A1(n_688), .A2(n_697), .B(n_731), .Y(n_730) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_695), .B(n_696), .Y(n_692) );
OAI21xp5_ASAP7_75t_L g887 ( .A1(n_698), .A2(n_888), .B(n_892), .Y(n_887) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g832 ( .A(n_700), .B(n_794), .Y(n_832) );
OR2x2_ASAP7_75t_L g862 ( .A(n_700), .B(n_748), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_700), .B(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OR2x2_ASAP7_75t_L g734 ( .A(n_703), .B(n_735), .Y(n_734) );
OR2x2_ASAP7_75t_L g744 ( .A(n_703), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g838 ( .A(n_703), .Y(n_838) );
BUFx3_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g708 ( .A(n_704), .Y(n_708) );
AOI21xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_711), .B(n_719), .Y(n_705) );
OAI22xp33_ASAP7_75t_L g741 ( .A1(n_706), .A2(n_742), .B1(n_744), .B2(n_747), .Y(n_741) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
AND2x2_ASAP7_75t_L g736 ( .A(n_708), .B(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_708), .B(n_764), .Y(n_763) );
OR2x6_ASAP7_75t_L g773 ( .A(n_708), .B(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g788 ( .A(n_708), .Y(n_788) );
INVx1_ASAP7_75t_L g774 ( .A(n_709), .Y(n_774) );
INVx1_ASAP7_75t_L g815 ( .A(n_709), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_715), .Y(n_711) );
INVx1_ASAP7_75t_L g849 ( .A(n_712), .Y(n_849) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_713), .B(n_718), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_713), .B(n_746), .Y(n_745) );
BUFx2_ASAP7_75t_L g824 ( .A(n_713), .Y(n_824) );
INVx3_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_715), .B(n_817), .Y(n_816) );
AND2x2_ASAP7_75t_L g823 ( .A(n_715), .B(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g861 ( .A(n_715), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_715), .B(n_737), .Y(n_863) );
AND2x2_ASAP7_75t_L g900 ( .A(n_715), .B(n_901), .Y(n_900) );
AND2x4_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .Y(n_715) );
INVx1_ASAP7_75t_L g872 ( .A(n_716), .Y(n_872) );
OR2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_724), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_721), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g851 ( .A(n_721), .B(n_782), .Y(n_851) );
INVx1_ASAP7_75t_L g867 ( .A(n_721), .Y(n_867) );
AOI322xp5_ASAP7_75t_L g899 ( .A1(n_721), .A2(n_900), .A3(n_902), .B1(n_904), .B2(n_905), .C1(n_907), .C2(n_908), .Y(n_899) );
AND2x4_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
AND2x4_ASAP7_75t_L g778 ( .A(n_722), .B(n_779), .Y(n_778) );
AND2x4_ASAP7_75t_L g828 ( .A(n_722), .B(n_829), .Y(n_828) );
OR2x2_ASAP7_75t_L g840 ( .A(n_722), .B(n_809), .Y(n_840) );
AND2x2_ASAP7_75t_L g743 ( .A(n_723), .B(n_730), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_723), .B(n_749), .Y(n_748) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_723), .Y(n_758) );
INVx1_ASAP7_75t_L g792 ( .A(n_723), .Y(n_792) );
INVx2_ASAP7_75t_L g903 ( .A(n_724), .Y(n_903) );
AOI221xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_733), .B1(n_736), .B2(n_738), .C(n_741), .Y(n_726) );
OR2x2_ASAP7_75t_L g889 ( .A(n_728), .B(n_890), .Y(n_889) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g793 ( .A(n_729), .B(n_794), .Y(n_793) );
AND2x2_ASAP7_75t_L g896 ( .A(n_729), .B(n_897), .Y(n_896) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g784 ( .A(n_735), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g800 ( .A(n_735), .Y(n_800) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_737), .Y(n_761) );
AND2x2_ASAP7_75t_L g892 ( .A(n_737), .B(n_827), .Y(n_892) );
AOI22xp5_ASAP7_75t_L g894 ( .A1(n_738), .A2(n_775), .B1(n_895), .B2(n_896), .Y(n_894) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_L g747 ( .A(n_740), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g805 ( .A(n_742), .Y(n_805) );
INVxp67_ASAP7_75t_SL g901 ( .A(n_745), .Y(n_901) );
INVx2_ASAP7_75t_L g755 ( .A(n_748), .Y(n_755) );
INVx1_ASAP7_75t_L g812 ( .A(n_749), .Y(n_812) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_749), .Y(n_856) );
AOI221xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_753), .B1(n_756), .B2(n_759), .C(n_762), .Y(n_750) );
INVx2_ASAP7_75t_L g767 ( .A(n_752), .Y(n_767) );
AND2x4_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_754), .B(n_778), .Y(n_777) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_755), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_756), .B(n_782), .Y(n_781) );
AND2x2_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
AND2x2_ASAP7_75t_L g791 ( .A(n_757), .B(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g865 ( .A(n_761), .Y(n_865) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_764), .B(n_788), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_764), .B(n_788), .Y(n_906) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_766), .B(n_849), .Y(n_848) );
NOR2x1p5_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
INVx1_ASAP7_75t_L g775 ( .A(n_767), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g770 ( .A(n_771), .B(n_786), .Y(n_770) );
AOI32xp33_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_775), .A3(n_776), .B1(n_780), .B2(n_783), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g907 ( .A(n_773), .Y(n_907) );
INVxp67_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g882 ( .A(n_779), .Y(n_882) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx2_ASAP7_75t_SL g804 ( .A(n_785), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_789), .B1(n_793), .B2(n_795), .Y(n_786) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g858 ( .A(n_792), .Y(n_858) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_794), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_794), .B(n_829), .Y(n_866) );
INVx1_ASAP7_75t_L g883 ( .A(n_795), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_820), .Y(n_796) );
AOI221xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_801), .B1(n_802), .B2(n_805), .C(n_806), .Y(n_797) );
AND2x4_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g814 ( .A(n_799), .Y(n_814) );
AND2x4_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_813), .B1(n_816), .B2(n_819), .Y(n_806) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_810), .Y(n_807) );
AND2x2_ASAP7_75t_L g908 ( .A(n_808), .B(n_904), .Y(n_908) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
OR2x2_ASAP7_75t_L g884 ( .A(n_809), .B(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OR2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
OR2x2_ASAP7_75t_L g876 ( .A(n_817), .B(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
AOI21xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_828), .B(n_830), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_825), .Y(n_821) );
OAI22xp33_ASAP7_75t_L g830 ( .A1(n_822), .A2(n_831), .B1(n_833), .B2(n_834), .Y(n_830) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_SL g852 ( .A(n_833), .Y(n_852) );
NOR3xp33_ASAP7_75t_L g835 ( .A(n_836), .B(n_875), .C(n_893), .Y(n_835) );
NAND3xp33_ASAP7_75t_SL g836 ( .A(n_837), .B(n_841), .C(n_850), .Y(n_836) );
INVx3_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OAI31xp33_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_844), .A3(n_845), .B(n_847), .Y(n_841) );
INVx2_ASAP7_75t_SL g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx2_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g895 ( .A(n_849), .Y(n_895) );
AOI211xp5_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_852), .B(n_853), .C(n_864), .Y(n_850) );
OAI22xp33_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_859), .B1(n_862), .B2(n_863), .Y(n_853) );
NOR2xp33_ASAP7_75t_SL g854 ( .A(n_855), .B(n_857), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_855), .B(n_880), .Y(n_879) );
OR2x2_ASAP7_75t_L g859 ( .A(n_860), .B(n_861), .Y(n_859) );
OAI22xp33_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_866), .B1(n_867), .B2(n_868), .Y(n_864) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_870), .B(n_873), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_870), .B(n_878), .Y(n_877) );
INVx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g878 ( .A(n_874), .Y(n_878) );
OAI221xp5_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_879), .B1(n_883), .B2(n_884), .C(n_887), .Y(n_875) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
OAI21xp5_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_898), .B(n_899), .Y(n_893) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_SL g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g914 ( .A(n_911), .Y(n_914) );
NOR2xp33_ASAP7_75t_L g915 ( .A(n_916), .B(n_917), .Y(n_915) );
BUFx3_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_921), .B(n_922), .Y(n_920) );
BUFx4f_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
endmodule