module fake_jpeg_28583_n_348 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_348);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_12),
.B(n_17),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_22),
.B(n_9),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_57),
.Y(n_87)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_22),
.A2(n_9),
.B1(n_17),
.B2(n_16),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_80),
.Y(n_103)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_21),
.B(n_9),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_34),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_82),
.Y(n_105)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_29),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_37),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_109),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_29),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_36),
.B1(n_25),
.B2(n_44),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_99),
.A2(n_100),
.B1(n_76),
.B2(n_67),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_51),
.B1(n_25),
.B2(n_44),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_27),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_37),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_79),
.A2(n_44),
.B1(n_46),
.B2(n_41),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_56),
.B1(n_62),
.B2(n_61),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_124),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_87),
.B(n_27),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_127),
.Y(n_158)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_73),
.B1(n_65),
.B2(n_72),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_110),
.B(n_105),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_130),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_34),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_146),
.C(n_40),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_133),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.Y(n_161)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_134),
.Y(n_172)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_136),
.Y(n_169)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_20),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_140),
.Y(n_165)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_143),
.Y(n_176)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

BUFx2_ASAP7_75t_SL g173 ( 
.A(n_142),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_20),
.Y(n_143)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_112),
.B(n_76),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_153),
.Y(n_162)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_111),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_32),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_152),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_84),
.B(n_32),
.Y(n_152)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_89),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_154),
.A2(n_155),
.B1(n_120),
.B2(n_88),
.Y(n_170)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_146),
.B1(n_142),
.B2(n_120),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_110),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_139),
.Y(n_177)
);

OAI22x1_ASAP7_75t_SL g168 ( 
.A1(n_133),
.A2(n_100),
.B1(n_99),
.B2(n_119),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_168),
.A2(n_144),
.B1(n_91),
.B2(n_95),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_174),
.B(n_132),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_182),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_168),
.A2(n_155),
.B1(n_130),
.B2(n_129),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_188),
.B1(n_190),
.B2(n_193),
.Y(n_197)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_180),
.A2(n_184),
.B1(n_186),
.B2(n_164),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_173),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_172),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_143),
.Y(n_182)
);

NOR2x1_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_125),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_191),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_163),
.A2(n_153),
.B1(n_149),
.B2(n_150),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_91),
.B1(n_88),
.B2(n_95),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_163),
.A2(n_146),
.B(n_134),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_166),
.C(n_174),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_154),
.B1(n_138),
.B2(n_137),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_128),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_189),
.B(n_165),
.Y(n_199)
);

NOR2x1_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_148),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_169),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_159),
.A2(n_136),
.B1(n_111),
.B2(n_122),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_176),
.B1(n_165),
.B2(n_97),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_195),
.A2(n_180),
.B1(n_185),
.B2(n_192),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_183),
.B(n_178),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_199),
.Y(n_215)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_156),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_201),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_157),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_209),
.B(n_192),
.C(n_187),
.D(n_158),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_158),
.B1(n_167),
.B2(n_164),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_204),
.A2(n_207),
.B1(n_190),
.B2(n_189),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_157),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_206),
.B(n_208),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_189),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_191),
.C(n_192),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_218),
.C(n_199),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_184),
.Y(n_211)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_217),
.Y(n_225)
);

OAI32xp33_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_183),
.A3(n_187),
.B1(n_190),
.B2(n_189),
.Y(n_216)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_188),
.B1(n_183),
.B2(n_170),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_197),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_225),
.B1(n_228),
.B2(n_207),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_205),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_237),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_222),
.B(n_201),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_233),
.B(n_198),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_206),
.Y(n_234)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_196),
.C(n_209),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_238),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_203),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_211),
.Y(n_239)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_227),
.B(n_202),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_247),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_218),
.C(n_217),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_242),
.C(n_243),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_214),
.C(n_203),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_212),
.C(n_213),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_224),
.B1(n_197),
.B2(n_216),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_246),
.A2(n_250),
.B1(n_252),
.B2(n_239),
.Y(n_260)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_175),
.B1(n_172),
.B2(n_160),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_223),
.C(n_221),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_172),
.C(n_160),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_211),
.B1(n_219),
.B2(n_220),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_219),
.B1(n_195),
.B2(n_204),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_181),
.B1(n_193),
.B2(n_159),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_167),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_230),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_256),
.B(n_31),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_231),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_266),
.C(n_268),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_236),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_263),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_264),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_243),
.A2(n_230),
.B(n_229),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_261),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_245),
.B(n_229),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_262),
.B(n_15),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_159),
.B(n_175),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_84),
.B(n_1),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_265),
.A2(n_250),
.B1(n_97),
.B2(n_89),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_241),
.A2(n_162),
.B1(n_175),
.B2(n_44),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_254),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_173),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_160),
.C(n_171),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_270),
.C(n_271),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_171),
.C(n_117),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_162),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_171),
.C(n_122),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_115),
.C(n_121),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_283),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_278),
.A2(n_38),
.B1(n_35),
.B2(n_3),
.Y(n_303)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_273),
.Y(n_279)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_286),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_258),
.A2(n_41),
.B(n_26),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_289),
.B(n_269),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_271),
.A2(n_17),
.B(n_19),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_285),
.A2(n_26),
.B(n_41),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_257),
.A2(n_20),
.B1(n_26),
.B2(n_46),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_16),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_287),
.B(n_288),
.Y(n_295)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_272),
.Y(n_288)
);

MAJx2_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_282),
.C(n_276),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_291),
.B(n_11),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_283),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_299),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_257),
.B(n_270),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_302),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_288),
.A2(n_268),
.B1(n_46),
.B2(n_115),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_301),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_281),
.A2(n_40),
.B1(n_38),
.B2(n_35),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_303),
.B(n_287),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_279),
.A2(n_10),
.B1(n_19),
.B2(n_3),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_305),
.A2(n_11),
.B1(n_19),
.B2(n_4),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_277),
.C(n_276),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_307),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_277),
.C(n_274),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_310),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_274),
.C(n_275),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_314),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_278),
.C(n_289),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_293),
.B(n_285),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_315),
.B(n_297),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_317),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_290),
.Y(n_317)
);

OAI21x1_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_301),
.B(n_298),
.Y(n_318)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_318),
.Y(n_335)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_315),
.A2(n_292),
.B(n_10),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_13),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_308),
.B(n_8),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_324),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_312),
.B(n_8),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_313),
.A2(n_13),
.B1(n_15),
.B2(n_6),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_327),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_13),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_321),
.Y(n_330)
);

OAI21x1_ASAP7_75t_L g339 ( 
.A1(n_330),
.A2(n_334),
.B(n_7),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_331),
.Y(n_340)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_328),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_329),
.A2(n_326),
.B(n_319),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_336),
.A2(n_337),
.B(n_338),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_322),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_330),
.A2(n_6),
.B(n_7),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_339),
.Y(n_341)
);

AOI321xp33_ASAP7_75t_L g342 ( 
.A1(n_340),
.A2(n_333),
.A3(n_332),
.B1(n_7),
.B2(n_15),
.C(n_31),
.Y(n_342)
);

A2O1A1Ixp33_ASAP7_75t_SL g345 ( 
.A1(n_342),
.A2(n_0),
.B(n_2),
.C(n_31),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_31),
.C(n_28),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_344),
.A2(n_345),
.B1(n_341),
.B2(n_2),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_0),
.B(n_28),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_28),
.Y(n_348)
);


endmodule