module fake_netlist_5_1378_n_1138 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_1138);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1138;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_785;
wire n_316;
wire n_855;
wire n_389;
wire n_843;
wire n_194;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_146;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_1055;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_916;
wire n_885;
wire n_1081;
wire n_452;
wire n_397;
wire n_525;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_155;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_983;
wire n_725;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_629;
wire n_590;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_1120;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_864;
wire n_443;
wire n_173;
wire n_859;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_604;
wire n_433;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_947;
wire n_936;
wire n_373;
wire n_147;
wire n_820;
wire n_757;
wire n_1090;
wire n_307;
wire n_633;
wire n_530;
wire n_439;
wire n_150;
wire n_1024;
wire n_1063;
wire n_556;
wire n_1107;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_186;
wire n_1124;
wire n_537;
wire n_902;
wire n_587;
wire n_191;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_171;
wire n_153;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_519;
wire n_406;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_1016;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_390;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_167;
wire n_976;
wire n_1096;
wire n_1095;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_570;
wire n_457;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_156;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_157;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_223;
wire n_1114;
wire n_1129;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_995;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_882;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_181;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_178;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_681;
wire n_584;
wire n_591;
wire n_922;
wire n_145;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_974;
wire n_395;
wire n_164;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_432;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_928;
wire n_445;
wire n_829;
wire n_749;
wire n_1064;
wire n_144;
wire n_858;
wire n_446;
wire n_923;
wire n_772;
wire n_691;
wire n_1134;
wire n_881;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_866;
wire n_573;
wire n_197;
wire n_969;
wire n_1069;
wire n_236;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_149;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_151;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_466;
wire n_239;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_846;
wire n_586;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_170;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_161;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_774;
wire n_365;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_176;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_182;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_679;
wire n_710;
wire n_795;
wire n_695;
wire n_832;
wire n_180;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_879;
wire n_421;
wire n_1072;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_202;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_1038;
wire n_409;
wire n_797;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_159;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_200;
wire n_1032;
wire n_1056;
wire n_162;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_806;
wire n_438;
wire n_713;
wire n_1011;
wire n_1123;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_348;
wire n_1029;
wire n_166;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

INVxp33_ASAP7_75t_SL g144 ( 
.A(n_134),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_113),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_70),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_60),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_26),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_8),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_32),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_66),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_65),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_98),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_58),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_124),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_48),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_115),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_7),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_74),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_24),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_72),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_69),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_15),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_125),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_126),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_101),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_89),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_14),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_122),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_9),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_35),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_108),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_121),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_128),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_137),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_135),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_45),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_55),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_140),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_102),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_100),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_132),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_59),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_106),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_111),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_1),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_146),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_153),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_180),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_148),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_152),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_154),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_155),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_163),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_171),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_172),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_151),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_174),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_176),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_183),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_183),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_145),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_185),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_149),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_186),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_188),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_150),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_203),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_202),
.Y(n_234)
);

INVxp67_ASAP7_75t_SL g235 ( 
.A(n_215),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_205),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_222),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_206),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_207),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_210),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_201),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_204),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_211),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_212),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_214),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_217),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_222),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_219),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_221),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_220),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_208),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_144),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_225),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_227),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_204),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_209),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_203),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_202),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_202),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_215),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_222),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_222),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_222),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_215),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_234),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

INVxp33_ASAP7_75t_SL g280 ( 
.A(n_256),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_239),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_241),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_239),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_253),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_237),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_246),
.Y(n_289)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_265),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_258),
.Y(n_291)
);

INVxp33_ASAP7_75t_SL g292 ( 
.A(n_238),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_264),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_230),
.Y(n_295)
);

BUFx2_ASAP7_75t_SL g296 ( 
.A(n_248),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_233),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_236),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_240),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_243),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_273),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_266),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_270),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_270),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_266),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_235),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_255),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_253),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_274),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_268),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_255),
.Y(n_314)
);

INVxp33_ASAP7_75t_SL g315 ( 
.A(n_259),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_274),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_245),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_232),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_232),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_267),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_283),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_278),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_299),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_280),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_283),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_282),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_280),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_285),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_289),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_286),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_305),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_293),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_286),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_307),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_318),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_319),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_315),
.B(n_242),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_300),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_317),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_296),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_311),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_288),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_306),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_309),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_295),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_281),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_311),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_297),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_298),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_312),
.Y(n_354)
);

BUFx2_ASAP7_75t_SL g355 ( 
.A(n_316),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_301),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_292),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_316),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_290),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_290),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_313),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_287),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_302),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_308),
.Y(n_364)
);

BUFx12f_ASAP7_75t_L g365 ( 
.A(n_322),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_315),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_346),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_350),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_337),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_323),
.B(n_284),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_340),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_342),
.Y(n_373)
);

INVx5_ASAP7_75t_L g374 ( 
.A(n_354),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_341),
.B(n_249),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_349),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_347),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_352),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_356),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_325),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_327),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_332),
.B(n_329),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_330),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_333),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_334),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_336),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_324),
.Y(n_389)
);

AND2x6_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_169),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_343),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_364),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_362),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_362),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_326),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_363),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_250),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_342),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_363),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_359),
.B(n_284),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_357),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_326),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_360),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_328),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_328),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_360),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_358),
.Y(n_407)
);

OAI22x1_ASAP7_75t_SL g408 ( 
.A1(n_358),
.A2(n_276),
.B1(n_275),
.B2(n_251),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_335),
.Y(n_409)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_355),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_331),
.B(n_252),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_335),
.B(n_284),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_345),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_345),
.B(n_231),
.Y(n_414)
);

OA21x2_ASAP7_75t_L g415 ( 
.A1(n_351),
.A2(n_304),
.B(n_303),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_351),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_338),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_337),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_348),
.B(n_254),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_341),
.B(n_257),
.Y(n_420)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_337),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_348),
.B(n_260),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_348),
.B(n_261),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_325),
.B(n_231),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_322),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_348),
.B(n_263),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_337),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_348),
.B(n_269),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_325),
.B(n_271),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_338),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_337),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_323),
.B(n_284),
.Y(n_432)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_337),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_348),
.B(n_310),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_338),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_338),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_338),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_337),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_338),
.Y(n_439)
);

INVx5_ASAP7_75t_L g440 ( 
.A(n_354),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g441 ( 
.A1(n_338),
.A2(n_314),
.B(n_187),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_338),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_338),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_338),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_338),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_338),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_350),
.Y(n_447)
);

NOR2x1_ASAP7_75t_L g448 ( 
.A(n_341),
.B(n_166),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_348),
.B(n_157),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_323),
.B(n_158),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_350),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_337),
.Y(n_452)
);

OAI21x1_ASAP7_75t_L g453 ( 
.A1(n_441),
.A2(n_187),
.B(n_169),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_376),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_376),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_386),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_378),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_378),
.Y(n_458)
);

NAND2x1_ASAP7_75t_L g459 ( 
.A(n_379),
.B(n_160),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_451),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_375),
.A2(n_276),
.B1(n_275),
.B2(n_420),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_380),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_380),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_375),
.B(n_147),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_420),
.A2(n_184),
.B1(n_199),
.B2(n_159),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_368),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_447),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_386),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_384),
.B(n_147),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_383),
.B(n_162),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_383),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_381),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_385),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_387),
.Y(n_474)
);

INVx6_ASAP7_75t_L g475 ( 
.A(n_386),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_384),
.B(n_164),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_367),
.B(n_159),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_417),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_373),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_435),
.B(n_445),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_435),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_412),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_367),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_418),
.B(n_167),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_371),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_367),
.B(n_377),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_372),
.Y(n_488)
);

BUFx12f_ASAP7_75t_L g489 ( 
.A(n_374),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_418),
.B(n_175),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_430),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_436),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_437),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_367),
.B(n_161),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_427),
.B(n_177),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_377),
.B(n_161),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_480),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_481),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_R g499 ( 
.A(n_480),
.B(n_373),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_489),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_474),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_474),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_489),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_479),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_460),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_466),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_481),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_464),
.B(n_377),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_456),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_479),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_472),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_461),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_467),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_486),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_483),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_483),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_486),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_488),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_465),
.B(n_366),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_469),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_482),
.Y(n_521)
);

NOR2xp67_ASAP7_75t_L g522 ( 
.A(n_478),
.B(n_398),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_494),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_488),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_484),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_456),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_496),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_476),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_491),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_484),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_476),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_491),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_475),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_484),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_484),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_475),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_492),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_492),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_SL g539 ( 
.A(n_499),
.B(n_484),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_509),
.Y(n_540)
);

NOR2x1p5_ASAP7_75t_L g541 ( 
.A(n_497),
.B(n_425),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_509),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_508),
.B(n_522),
.Y(n_543)
);

OR2x6_ASAP7_75t_L g544 ( 
.A(n_508),
.B(n_487),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_519),
.B(n_419),
.Y(n_545)
);

BUFx4f_ASAP7_75t_L g546 ( 
.A(n_509),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_501),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_501),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_518),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_502),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_509),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_502),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_520),
.B(n_416),
.Y(n_553)
);

NAND3xp33_ASAP7_75t_L g554 ( 
.A(n_523),
.B(n_448),
.C(n_397),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_530),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_504),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_526),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_527),
.B(n_397),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_528),
.B(n_429),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_532),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_506),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_534),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_538),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_535),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_504),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_520),
.B(n_531),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_498),
.B(n_429),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_526),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_510),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_514),
.Y(n_570)
);

BUFx10_ASAP7_75t_L g571 ( 
.A(n_513),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_533),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_510),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_521),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_517),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_511),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_524),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_529),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_537),
.Y(n_579)
);

AND3x1_ASAP7_75t_L g580 ( 
.A(n_512),
.B(n_394),
.C(n_393),
.Y(n_580)
);

INVxp33_ASAP7_75t_L g581 ( 
.A(n_507),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_505),
.B(n_413),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_526),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_515),
.A2(n_470),
.B1(n_413),
.B2(n_415),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_526),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_525),
.Y(n_586)
);

OAI22xp33_ASAP7_75t_L g587 ( 
.A1(n_516),
.A2(n_493),
.B1(n_374),
.B2(n_440),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_525),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_536),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_500),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_525),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_503),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_518),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_518),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_533),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_519),
.B(n_412),
.Y(n_596)
);

AND3x1_ASAP7_75t_L g597 ( 
.A(n_519),
.B(n_394),
.C(n_393),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_518),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_533),
.B(n_412),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_519),
.B(n_413),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_509),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_501),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_506),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_519),
.B(n_415),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_506),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_501),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_518),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_519),
.A2(n_470),
.B1(n_415),
.B2(n_450),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_518),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_508),
.B(n_422),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_518),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_501),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_530),
.Y(n_613)
);

CKINVDCx14_ASAP7_75t_R g614 ( 
.A(n_499),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_519),
.B(n_396),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_533),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_509),
.Y(n_617)
);

INVxp67_ASAP7_75t_R g618 ( 
.A(n_499),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_518),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_554),
.B(n_389),
.Y(n_620)
);

OR2x6_ASAP7_75t_L g621 ( 
.A(n_544),
.B(n_456),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_573),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_614),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_558),
.B(n_389),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_604),
.B(n_545),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_545),
.B(n_455),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_568),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_574),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_572),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_570),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_594),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_596),
.B(n_470),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_572),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_575),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_577),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_555),
.B(n_468),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_578),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_600),
.B(n_389),
.Y(n_638)
);

BUFx2_ASAP7_75t_L g639 ( 
.A(n_595),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_615),
.B(n_395),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_568),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_579),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_549),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_555),
.B(n_468),
.Y(n_644)
);

INVx3_ASAP7_75t_R g645 ( 
.A(n_605),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_600),
.B(n_455),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_560),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_599),
.B(n_450),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_547),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_544),
.B(n_457),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_603),
.B(n_409),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_559),
.B(n_409),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_544),
.B(n_457),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_548),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_597),
.B(n_389),
.Y(n_655)
);

INVx8_ASAP7_75t_L g656 ( 
.A(n_542),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_563),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_595),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_616),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_593),
.B(n_458),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_598),
.Y(n_661)
);

NAND2x1p5_ASAP7_75t_L g662 ( 
.A(n_543),
.B(n_456),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_607),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_542),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_609),
.B(n_458),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_550),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_542),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_546),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_611),
.B(n_402),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_616),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_562),
.Y(n_671)
);

INVx6_ASAP7_75t_L g672 ( 
.A(n_571),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_550),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_552),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_561),
.B(n_411),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_619),
.B(n_462),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_571),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_599),
.B(n_450),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_556),
.Y(n_679)
);

AO22x2_ASAP7_75t_L g680 ( 
.A1(n_610),
.A2(n_399),
.B1(n_396),
.B2(n_406),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_540),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_580),
.B(n_391),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_542),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_546),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_610),
.B(n_462),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_556),
.B(n_463),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_565),
.B(n_463),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_540),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_565),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_569),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_587),
.B(n_391),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_614),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_562),
.B(n_468),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_602),
.Y(n_694)
);

BUFx4f_ASAP7_75t_L g695 ( 
.A(n_592),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_564),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_602),
.Y(n_697)
);

AND2x6_ASAP7_75t_L g698 ( 
.A(n_586),
.B(n_456),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_681),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_658),
.B(n_587),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_625),
.B(n_631),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_620),
.A2(n_633),
.B1(n_639),
.B2(n_629),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_658),
.B(n_374),
.Y(n_703)
);

NOR2x1_ASAP7_75t_L g704 ( 
.A(n_638),
.B(n_543),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_634),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_630),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_672),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_635),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_637),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_643),
.B(n_589),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_624),
.A2(n_553),
.B1(n_584),
.B2(n_608),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_632),
.A2(n_553),
.B1(n_584),
.B2(n_608),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_643),
.B(n_582),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_672),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_642),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_658),
.B(n_374),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_625),
.B(n_606),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_647),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_671),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_631),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_621),
.B(n_564),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_656),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_657),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_661),
.Y(n_724)
);

AND3x4_ASAP7_75t_L g725 ( 
.A(n_670),
.B(n_401),
.C(n_425),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_659),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_646),
.B(n_567),
.Y(n_727)
);

AO21x2_ASAP7_75t_L g728 ( 
.A1(n_655),
.A2(n_453),
.B(n_441),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_648),
.A2(n_566),
.B1(n_582),
.B2(n_165),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_623),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_649),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_651),
.B(n_576),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_640),
.B(n_566),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_621),
.B(n_613),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_663),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_663),
.B(n_581),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_650),
.Y(n_737)
);

CKINVDCx8_ASAP7_75t_R g738 ( 
.A(n_692),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_626),
.B(n_612),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_650),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_621),
.B(n_613),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_654),
.Y(n_742)
);

NAND3xp33_ASAP7_75t_SL g743 ( 
.A(n_682),
.B(n_426),
.C(n_423),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_653),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_653),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_690),
.B(n_612),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_669),
.Y(n_747)
);

AO22x2_ASAP7_75t_L g748 ( 
.A1(n_691),
.A2(n_588),
.B1(n_585),
.B2(n_583),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_666),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_659),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_694),
.B(n_697),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_659),
.B(n_592),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_652),
.B(n_407),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_681),
.Y(n_754)
);

BUFx2_ASAP7_75t_L g755 ( 
.A(n_695),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_673),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_675),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_681),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_674),
.Y(n_759)
);

AND2x6_ASAP7_75t_L g760 ( 
.A(n_668),
.B(n_540),
.Y(n_760)
);

AND2x2_ASAP7_75t_SL g761 ( 
.A(n_695),
.B(n_398),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_660),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_718),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_752),
.B(n_592),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_757),
.B(n_677),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_737),
.B(n_680),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_714),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_740),
.B(n_680),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_732),
.B(n_645),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_705),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_704),
.B(n_696),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_704),
.B(n_696),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_738),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_711),
.B(n_685),
.C(n_192),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_753),
.B(n_592),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_743),
.A2(n_700),
.B1(n_711),
.B2(n_712),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_744),
.B(n_622),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_745),
.B(n_628),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_720),
.B(n_665),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_720),
.B(n_676),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_761),
.B(n_391),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_701),
.B(n_676),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_733),
.B(n_407),
.Y(n_783)
);

O2A1O1Ixp5_ASAP7_75t_L g784 ( 
.A1(n_703),
.A2(n_539),
.B(n_644),
.C(n_636),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_712),
.A2(n_678),
.B1(n_407),
.B2(n_590),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_747),
.B(n_407),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_713),
.B(n_636),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_709),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_707),
.B(n_391),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_701),
.B(n_662),
.Y(n_790)
);

NOR2xp67_ASAP7_75t_L g791 ( 
.A(n_735),
.B(n_627),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_723),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_724),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_736),
.B(n_727),
.Y(n_794)
);

AOI221xp5_ASAP7_75t_L g795 ( 
.A1(n_702),
.A2(n_168),
.B1(n_200),
.B2(n_189),
.C(n_191),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_721),
.B(n_644),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_716),
.A2(n_428),
.B(n_662),
.C(n_449),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_719),
.B(n_693),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_762),
.B(n_679),
.Y(n_799)
);

NOR2xp67_ASAP7_75t_L g800 ( 
.A(n_726),
.B(n_627),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_706),
.B(n_689),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_721),
.B(n_693),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_729),
.A2(n_539),
.B(n_165),
.C(n_196),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_708),
.B(n_715),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_750),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_725),
.B(n_408),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_710),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_717),
.A2(n_405),
.B(n_156),
.C(n_668),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_729),
.B(n_440),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_731),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_748),
.A2(n_656),
.B(n_664),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_751),
.B(n_686),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_751),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_734),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_734),
.B(n_398),
.Y(n_815)
);

AND2x6_ASAP7_75t_SL g816 ( 
.A(n_730),
.B(n_414),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_742),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_739),
.B(n_687),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_741),
.B(n_440),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_741),
.A2(n_684),
.B1(n_410),
.B2(n_541),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_749),
.B(n_687),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_756),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_755),
.B(n_440),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_759),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_748),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_746),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_722),
.B(n_403),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_722),
.B(n_403),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_699),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_699),
.Y(n_830)
);

OR2x6_ASAP7_75t_L g831 ( 
.A(n_754),
.B(n_656),
.Y(n_831)
);

INVx4_ASAP7_75t_L g832 ( 
.A(n_754),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_770),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_793),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_831),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_814),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_825),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_807),
.B(n_754),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_798),
.B(n_764),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_787),
.B(n_758),
.Y(n_840)
);

AND2x2_ASAP7_75t_SL g841 ( 
.A(n_776),
.B(n_684),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_788),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_767),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_771),
.B(n_758),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_792),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_813),
.B(n_618),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_831),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_773),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_784),
.B(n_772),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_766),
.Y(n_850)
);

CKINVDCx6p67_ASAP7_75t_R g851 ( 
.A(n_831),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_766),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_794),
.B(n_760),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_774),
.B(n_641),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_826),
.B(n_641),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_805),
.B(n_688),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_782),
.B(n_760),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_763),
.B(n_688),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_808),
.A2(n_760),
.B(n_196),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_803),
.A2(n_760),
.B(n_199),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_817),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_810),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_791),
.B(n_403),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_822),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_768),
.B(n_410),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_768),
.B(n_410),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_824),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_811),
.B(n_664),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_786),
.B(n_382),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_804),
.Y(n_870)
);

NAND2x1p5_ASAP7_75t_L g871 ( 
.A(n_781),
.B(n_667),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_790),
.B(n_591),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_779),
.B(n_591),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_780),
.B(n_698),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_829),
.B(n_667),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_777),
.B(n_698),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_830),
.B(n_683),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_778),
.B(n_698),
.Y(n_878)
);

INVxp33_ASAP7_75t_L g879 ( 
.A(n_783),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_795),
.A2(n_184),
.B(n_424),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_806),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_789),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_859),
.A2(n_797),
.B(n_815),
.Y(n_883)
);

AOI21x1_ASAP7_75t_L g884 ( 
.A1(n_849),
.A2(n_828),
.B(n_827),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_868),
.B(n_800),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_849),
.A2(n_819),
.B(n_809),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_850),
.B(n_812),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_860),
.A2(n_802),
.B(n_796),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_852),
.B(n_812),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_870),
.B(n_818),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_836),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_835),
.B(n_847),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_880),
.A2(n_765),
.B(n_769),
.C(n_785),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_841),
.A2(n_820),
.B(n_821),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_837),
.A2(n_823),
.B(n_775),
.C(n_799),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_838),
.B(n_832),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_841),
.A2(n_821),
.B(n_801),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_845),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_845),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_851),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_848),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_865),
.B(n_832),
.Y(n_902)
);

INVx5_ASAP7_75t_L g903 ( 
.A(n_835),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_863),
.A2(n_683),
.B(n_816),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_848),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_865),
.B(n_698),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_866),
.A2(n_601),
.B1(n_617),
.B2(n_551),
.Y(n_907)
);

BUFx8_ASAP7_75t_L g908 ( 
.A(n_843),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_881),
.B(n_365),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_881),
.B(n_365),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_836),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_866),
.A2(n_601),
.B(n_551),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_857),
.B(n_728),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_833),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_836),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_853),
.B(n_728),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_854),
.A2(n_400),
.B(n_459),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_851),
.A2(n_403),
.B1(n_400),
.B2(n_557),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_879),
.B(n_401),
.Y(n_919)
);

AND2x6_ASAP7_75t_L g920 ( 
.A(n_835),
.B(n_557),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_882),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_882),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_868),
.A2(n_404),
.B(n_557),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_879),
.B(n_0),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_876),
.A2(n_404),
.B(n_454),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_878),
.A2(n_473),
.B(n_471),
.Y(n_926)
);

INVxp67_ASAP7_75t_L g927 ( 
.A(n_844),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_842),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_869),
.A2(n_392),
.B(n_477),
.C(n_493),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_844),
.A2(n_490),
.B(n_485),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_892),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_883),
.A2(n_886),
.B1(n_888),
.B2(n_924),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_903),
.B(n_835),
.Y(n_933)
);

AOI33xp33_ASAP7_75t_L g934 ( 
.A1(n_893),
.A2(n_861),
.A3(n_846),
.B1(n_867),
.B2(n_864),
.B3(n_862),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_900),
.B(n_869),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_904),
.A2(n_871),
.B1(n_847),
.B2(n_874),
.Y(n_936)
);

NOR2x1_ASAP7_75t_L g937 ( 
.A(n_905),
.B(n_847),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_905),
.B(n_847),
.Y(n_938)
);

AO21x1_ASAP7_75t_L g939 ( 
.A1(n_884),
.A2(n_834),
.B(n_877),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_927),
.B(n_839),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_897),
.B(n_855),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_895),
.B(n_858),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_885),
.B(n_840),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_L g944 ( 
.A(n_926),
.B(n_872),
.C(n_873),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_894),
.A2(n_877),
.B(n_875),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_903),
.B(n_877),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_921),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_905),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_934),
.B(n_925),
.Y(n_949)
);

INVx5_ASAP7_75t_L g950 ( 
.A(n_948),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_948),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_932),
.B(n_887),
.Y(n_952)
);

NAND2x1p5_ASAP7_75t_L g953 ( 
.A(n_937),
.B(n_903),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_940),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_932),
.B(n_889),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_943),
.B(n_885),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_944),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_SL g958 ( 
.A1(n_933),
.A2(n_901),
.B(n_922),
.C(n_910),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_931),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_931),
.B(n_890),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_935),
.B(n_914),
.Y(n_961)
);

OAI21x1_ASAP7_75t_L g962 ( 
.A1(n_939),
.A2(n_911),
.B(n_891),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_947),
.Y(n_963)
);

BUFx8_ASAP7_75t_SL g964 ( 
.A(n_942),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_SL g965 ( 
.A(n_938),
.B(n_909),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_946),
.B(n_898),
.Y(n_966)
);

OAI22xp33_ASAP7_75t_L g967 ( 
.A1(n_941),
.A2(n_906),
.B1(n_907),
.B2(n_902),
.Y(n_967)
);

BUFx8_ASAP7_75t_L g968 ( 
.A(n_936),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_945),
.A2(n_916),
.B(n_913),
.Y(n_969)
);

BUFx12f_ASAP7_75t_L g970 ( 
.A(n_940),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_940),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_932),
.A2(n_929),
.B(n_919),
.C(n_912),
.Y(n_972)
);

NAND2xp33_ASAP7_75t_SL g973 ( 
.A(n_932),
.B(n_896),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_932),
.A2(n_923),
.B(n_918),
.C(n_917),
.Y(n_974)
);

INVxp67_ASAP7_75t_SL g975 ( 
.A(n_968),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_964),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_SL g977 ( 
.A1(n_957),
.A2(n_908),
.B1(n_899),
.B2(n_930),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_953),
.Y(n_978)
);

BUFx6f_ASAP7_75t_SL g979 ( 
.A(n_959),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_954),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_971),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_960),
.B(n_928),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_980),
.B(n_949),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_978),
.A2(n_962),
.B(n_951),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_983),
.B(n_975),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_984),
.A2(n_952),
.B1(n_955),
.B2(n_974),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_986),
.A2(n_985),
.B(n_981),
.Y(n_987)
);

AO21x2_ASAP7_75t_L g988 ( 
.A1(n_986),
.A2(n_958),
.B(n_979),
.Y(n_988)
);

OA21x2_ASAP7_75t_L g989 ( 
.A1(n_987),
.A2(n_976),
.B(n_969),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_988),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_989),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_990),
.Y(n_992)
);

INVxp67_ASAP7_75t_L g993 ( 
.A(n_991),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_992),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_994),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_993),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_994),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_997),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_996),
.A2(n_988),
.B1(n_979),
.B2(n_989),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_995),
.B(n_987),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_1000),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_998),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_1001),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_1002),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_1003),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_1004),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_1005),
.B(n_999),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_1006),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_1008),
.B(n_992),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_1007),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_1009),
.B(n_956),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_1010),
.B(n_950),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_1011),
.B(n_970),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1012),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_1011),
.B(n_950),
.Y(n_1015)
);

AND2x4_ASAP7_75t_SL g1016 ( 
.A(n_1013),
.B(n_963),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_1015),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1014),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_1016),
.Y(n_1019)
);

OR2x2_ASAP7_75t_L g1020 ( 
.A(n_1017),
.B(n_973),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1020),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1019),
.B(n_1018),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_1022),
.B(n_950),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_1021),
.B(n_966),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_1023),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1024),
.B(n_965),
.Y(n_1026)
);

AND2x2_ASAP7_75t_SL g1027 ( 
.A(n_1025),
.B(n_982),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_1026),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1027),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1028),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_1030),
.B(n_977),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_1029),
.Y(n_1032)
);

OAI222xp33_ASAP7_75t_L g1033 ( 
.A1(n_1030),
.A2(n_982),
.B1(n_972),
.B2(n_961),
.C1(n_198),
.C2(n_195),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1032),
.Y(n_1034)
);

AOI221xp5_ASAP7_75t_L g1035 ( 
.A1(n_1031),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.C(n_197),
.Y(n_1035)
);

OAI21xp33_ASAP7_75t_L g1036 ( 
.A1(n_1033),
.A2(n_178),
.B(n_966),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_1034),
.A2(n_967),
.B(n_390),
.Y(n_1037)
);

AO21x1_ASAP7_75t_L g1038 ( 
.A1(n_1035),
.A2(n_968),
.B(n_0),
.Y(n_1038)
);

OR2x2_ASAP7_75t_L g1039 ( 
.A(n_1038),
.B(n_1036),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1037),
.Y(n_1040)
);

NAND2xp33_ASAP7_75t_L g1041 ( 
.A(n_1039),
.B(n_390),
.Y(n_1041)
);

NOR2x1_ASAP7_75t_L g1042 ( 
.A(n_1040),
.B(n_1),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_1042),
.A2(n_4),
.B(n_2),
.C(n_3),
.Y(n_1043)
);

AOI211xp5_ASAP7_75t_L g1044 ( 
.A1(n_1041),
.A2(n_4),
.B(n_2),
.C(n_3),
.Y(n_1044)
);

NAND4xp25_ASAP7_75t_L g1045 ( 
.A(n_1044),
.B(n_7),
.C(n_5),
.D(n_6),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1043),
.A2(n_390),
.B(n_5),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_1046),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1045),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_1048),
.B(n_6),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1047),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_1048),
.B(n_8),
.Y(n_1051)
);

NAND4xp25_ASAP7_75t_L g1052 ( 
.A(n_1050),
.B(n_9),
.C(n_10),
.D(n_11),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_1049),
.B(n_10),
.Y(n_1053)
);

NAND4xp25_ASAP7_75t_L g1054 ( 
.A(n_1051),
.B(n_11),
.C(n_12),
.D(n_13),
.Y(n_1054)
);

NAND4xp75_ASAP7_75t_L g1055 ( 
.A(n_1053),
.B(n_12),
.C(n_13),
.D(n_14),
.Y(n_1055)
);

NOR2x1_ASAP7_75t_L g1056 ( 
.A(n_1054),
.B(n_15),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_1056),
.B(n_1052),
.Y(n_1057)
);

NAND4xp75_ASAP7_75t_L g1058 ( 
.A(n_1055),
.B(n_16),
.C(n_17),
.D(n_18),
.Y(n_1058)
);

NAND3xp33_ASAP7_75t_L g1059 ( 
.A(n_1057),
.B(n_908),
.C(n_16),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_SL g1060 ( 
.A(n_1058),
.B(n_17),
.C(n_19),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_1060),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1059),
.B(n_20),
.Y(n_1062)
);

NOR3xp33_ASAP7_75t_L g1063 ( 
.A(n_1062),
.B(n_21),
.C(n_22),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_1061),
.Y(n_1064)
);

NAND4xp25_ASAP7_75t_L g1065 ( 
.A(n_1064),
.B(n_22),
.C(n_23),
.D(n_24),
.Y(n_1065)
);

NAND4xp25_ASAP7_75t_L g1066 ( 
.A(n_1063),
.B(n_23),
.C(n_25),
.D(n_27),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1066),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1065),
.Y(n_1068)
);

NOR2x1_ASAP7_75t_L g1069 ( 
.A(n_1066),
.B(n_25),
.Y(n_1069)
);

NAND4xp75_ASAP7_75t_L g1070 ( 
.A(n_1068),
.B(n_495),
.C(n_490),
.D(n_485),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_SL g1071 ( 
.A1(n_1067),
.A2(n_446),
.B1(n_444),
.B2(n_443),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_L g1072 ( 
.A(n_1069),
.B(n_28),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_1072),
.Y(n_1073)
);

OAI221xp5_ASAP7_75t_L g1074 ( 
.A1(n_1071),
.A2(n_442),
.B1(n_439),
.B2(n_31),
.C(n_33),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_1073),
.Y(n_1075)
);

XOR2xp5_ASAP7_75t_L g1076 ( 
.A(n_1074),
.B(n_1070),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_1075),
.Y(n_1077)
);

AOI22x1_ASAP7_75t_L g1078 ( 
.A1(n_1076),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_1078)
);

AOI22x1_ASAP7_75t_L g1079 ( 
.A1(n_1077),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_1078),
.Y(n_1080)
);

NAND5xp2_ASAP7_75t_L g1081 ( 
.A(n_1080),
.B(n_39),
.C(n_40),
.D(n_41),
.E(n_42),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_1079),
.A2(n_390),
.B1(n_432),
.B2(n_370),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1082),
.B(n_1081),
.Y(n_1083)
);

OAI31xp33_ASAP7_75t_L g1084 ( 
.A1(n_1081),
.A2(n_495),
.A3(n_432),
.B(n_370),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_1083),
.A2(n_432),
.B1(n_370),
.B2(n_369),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_1084),
.A2(n_390),
.B1(n_369),
.B2(n_433),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_SL g1087 ( 
.A1(n_1083),
.A2(n_433),
.B1(n_431),
.B2(n_421),
.Y(n_1087)
);

AOI21xp33_ASAP7_75t_SL g1088 ( 
.A1(n_1086),
.A2(n_1085),
.B(n_1087),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_SL g1089 ( 
.A1(n_1086),
.A2(n_920),
.B1(n_44),
.B2(n_46),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_SL g1090 ( 
.A1(n_1086),
.A2(n_433),
.B1(n_431),
.B2(n_421),
.Y(n_1090)
);

AO21x2_ASAP7_75t_L g1091 ( 
.A1(n_1088),
.A2(n_434),
.B(n_43),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1090),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_1089),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1092),
.A2(n_47),
.B(n_49),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1093),
.A2(n_431),
.B1(n_421),
.B2(n_369),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_SL g1096 ( 
.A1(n_1091),
.A2(n_475),
.B1(n_51),
.B2(n_52),
.Y(n_1096)
);

XNOR2xp5_ASAP7_75t_L g1097 ( 
.A(n_1096),
.B(n_50),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1094),
.A2(n_1095),
.B(n_920),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1096),
.B(n_53),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1097),
.B(n_54),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1099),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1098),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_1097),
.B(n_56),
.Y(n_1103)
);

AOI221xp5_ASAP7_75t_L g1104 ( 
.A1(n_1097),
.A2(n_57),
.B1(n_61),
.B2(n_62),
.C(n_63),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1097),
.A2(n_475),
.B1(n_452),
.B2(n_438),
.Y(n_1105)
);

AOI21xp33_ASAP7_75t_L g1106 ( 
.A1(n_1097),
.A2(n_64),
.B(n_67),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1097),
.A2(n_920),
.B1(n_438),
.B2(n_452),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1097),
.B(n_68),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1097),
.B(n_71),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1097),
.A2(n_920),
.B(n_75),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1097),
.B(n_73),
.Y(n_1111)
);

AO21x1_ASAP7_75t_L g1112 ( 
.A1(n_1099),
.A2(n_76),
.B(n_77),
.Y(n_1112)
);

INVx4_ASAP7_75t_L g1113 ( 
.A(n_1102),
.Y(n_1113)
);

AOI22x1_ASAP7_75t_L g1114 ( 
.A1(n_1101),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1111),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_1108),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_1109),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1100),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1103),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1105),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1112),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1113),
.A2(n_1110),
.B(n_1106),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_R g1123 ( 
.A1(n_1117),
.A2(n_1118),
.B1(n_1119),
.B2(n_1116),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1115),
.A2(n_1107),
.B1(n_1104),
.B2(n_83),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1121),
.A2(n_856),
.B1(n_452),
.B2(n_438),
.Y(n_1125)
);

AOI221xp5_ASAP7_75t_L g1126 ( 
.A1(n_1120),
.A2(n_81),
.B1(n_82),
.B2(n_84),
.C(n_85),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_SL g1127 ( 
.A1(n_1114),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1122),
.A2(n_90),
.B(n_91),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1123),
.A2(n_92),
.B(n_93),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1124),
.B(n_94),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_SL g1131 ( 
.A1(n_1130),
.A2(n_1127),
.B1(n_1126),
.B2(n_1125),
.Y(n_1131)
);

AO21x2_ASAP7_75t_L g1132 ( 
.A1(n_1131),
.A2(n_1128),
.B(n_1129),
.Y(n_1132)
);

OA21x2_ASAP7_75t_L g1133 ( 
.A1(n_1132),
.A2(n_95),
.B(n_96),
.Y(n_1133)
);

OAI221xp5_ASAP7_75t_R g1134 ( 
.A1(n_1133),
.A2(n_97),
.B1(n_99),
.B2(n_103),
.C(n_104),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1134),
.A2(n_105),
.B(n_107),
.Y(n_1135)
);

AOI21xp33_ASAP7_75t_SL g1136 ( 
.A1(n_1135),
.A2(n_110),
.B(n_112),
.Y(n_1136)
);

AOI211xp5_ASAP7_75t_L g1137 ( 
.A1(n_1136),
.A2(n_915),
.B(n_117),
.C(n_118),
.Y(n_1137)
);

AOI211xp5_ASAP7_75t_L g1138 ( 
.A1(n_1137),
.A2(n_114),
.B(n_119),
.C(n_120),
.Y(n_1138)
);


endmodule