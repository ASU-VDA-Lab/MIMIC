module real_aes_2275_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g555 ( .A(n_0), .B(n_170), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_1), .B(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g131 ( .A(n_2), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_3), .B(n_478), .Y(n_510) );
NAND2xp33_ASAP7_75t_SL g504 ( .A(n_4), .B(n_152), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_5), .B(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g497 ( .A(n_6), .Y(n_497) );
INVx1_ASAP7_75t_L g229 ( .A(n_7), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g806 ( .A(n_8), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_9), .Y(n_221) );
AND2x2_ASAP7_75t_L g508 ( .A(n_10), .B(n_121), .Y(n_508) );
INVx2_ASAP7_75t_L g122 ( .A(n_11), .Y(n_122) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_12), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g804 ( .A(n_12), .B(n_805), .C(n_807), .Y(n_804) );
INVx1_ASAP7_75t_L g171 ( .A(n_13), .Y(n_171) );
AOI221x1_ASAP7_75t_L g500 ( .A1(n_14), .A2(n_154), .B1(n_477), .B2(n_501), .C(n_503), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_15), .B(n_478), .Y(n_486) );
INVx1_ASAP7_75t_L g467 ( .A(n_16), .Y(n_467) );
INVx1_ASAP7_75t_L g168 ( .A(n_17), .Y(n_168) );
INVx1_ASAP7_75t_SL g143 ( .A(n_18), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_19), .B(n_146), .Y(n_185) );
AOI33xp33_ASAP7_75t_L g238 ( .A1(n_20), .A2(n_51), .A3(n_128), .B1(n_139), .B2(n_239), .B3(n_240), .Y(n_238) );
AOI221xp5_ASAP7_75t_SL g476 ( .A1(n_21), .A2(n_40), .B1(n_477), .B2(n_478), .C(n_479), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_22), .A2(n_477), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_23), .B(n_170), .Y(n_513) );
INVx1_ASAP7_75t_L g768 ( .A(n_24), .Y(n_768) );
INVx1_ASAP7_75t_L g214 ( .A(n_25), .Y(n_214) );
OR2x2_ASAP7_75t_L g123 ( .A(n_26), .B(n_93), .Y(n_123) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_26), .A2(n_93), .B(n_122), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_27), .B(n_173), .Y(n_490) );
INVxp67_ASAP7_75t_L g499 ( .A(n_28), .Y(n_499) );
AND2x2_ASAP7_75t_L g544 ( .A(n_29), .B(n_120), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_30), .B(n_126), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_31), .A2(n_477), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_32), .B(n_173), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_33), .A2(n_43), .B1(n_758), .B2(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_33), .Y(n_758) );
AND2x2_ASAP7_75t_L g133 ( .A(n_34), .B(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g138 ( .A(n_34), .Y(n_138) );
AND2x2_ASAP7_75t_L g152 ( .A(n_34), .B(n_131), .Y(n_152) );
OR2x6_ASAP7_75t_L g465 ( .A(n_35), .B(n_466), .Y(n_465) );
INVxp67_ASAP7_75t_L g807 ( .A(n_35), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_36), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_37), .B(n_126), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_38), .A2(n_155), .B1(n_161), .B2(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_39), .B(n_187), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_41), .A2(n_82), .B1(n_136), .B2(n_477), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_42), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g759 ( .A(n_43), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_44), .B(n_170), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_45), .A2(n_786), .B1(n_787), .B2(n_790), .Y(n_785) );
INVx1_ASAP7_75t_L g790 ( .A(n_45), .Y(n_790) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_46), .B(n_189), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_47), .B(n_146), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_48), .Y(n_182) );
AND2x2_ASAP7_75t_L g558 ( .A(n_49), .B(n_120), .Y(n_558) );
OAI22xp5_ASAP7_75t_SL g787 ( .A1(n_49), .A2(n_78), .B1(n_788), .B2(n_789), .Y(n_787) );
INVxp67_ASAP7_75t_L g788 ( .A(n_49), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_50), .B(n_120), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_52), .B(n_146), .Y(n_260) );
INVx1_ASAP7_75t_L g129 ( .A(n_53), .Y(n_129) );
INVx1_ASAP7_75t_L g148 ( .A(n_53), .Y(n_148) );
AND2x2_ASAP7_75t_L g261 ( .A(n_54), .B(n_120), .Y(n_261) );
AOI221xp5_ASAP7_75t_L g227 ( .A1(n_55), .A2(n_74), .B1(n_126), .B2(n_136), .C(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_56), .B(n_126), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_57), .B(n_478), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_58), .B(n_155), .Y(n_223) );
AOI21xp5_ASAP7_75t_SL g194 ( .A1(n_59), .A2(n_136), .B(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g523 ( .A(n_60), .B(n_120), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_61), .B(n_173), .Y(n_556) );
INVx1_ASAP7_75t_L g164 ( .A(n_62), .Y(n_164) );
AND2x2_ASAP7_75t_SL g491 ( .A(n_63), .B(n_121), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_64), .B(n_170), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_65), .Y(n_809) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_66), .A2(n_477), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g259 ( .A(n_67), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_68), .B(n_173), .Y(n_514) );
AND2x2_ASAP7_75t_SL g529 ( .A(n_69), .B(n_189), .Y(n_529) );
OAI22xp5_ASAP7_75t_SL g796 ( .A1(n_70), .A2(n_92), .B1(n_797), .B2(n_798), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_70), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_71), .A2(n_136), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g134 ( .A(n_72), .Y(n_134) );
INVx1_ASAP7_75t_L g150 ( .A(n_72), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_73), .B(n_126), .Y(n_241) );
AND2x2_ASAP7_75t_L g153 ( .A(n_75), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g165 ( .A(n_76), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_77), .A2(n_136), .B(n_142), .Y(n_135) );
INVx1_ASAP7_75t_L g789 ( .A(n_78), .Y(n_789) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_79), .A2(n_136), .B(n_184), .C(n_188), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_80), .B(n_478), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_81), .A2(n_85), .B1(n_126), .B2(n_478), .Y(n_527) );
INVx1_ASAP7_75t_L g468 ( .A(n_83), .Y(n_468) );
AND2x2_ASAP7_75t_SL g192 ( .A(n_84), .B(n_154), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_86), .A2(n_136), .B1(n_236), .B2(n_237), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_87), .B(n_170), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_88), .B(n_170), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_89), .B(n_777), .Y(n_776) );
XNOR2x2_ASAP7_75t_SL g755 ( .A(n_90), .B(n_756), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_91), .A2(n_477), .B(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_SL g402 ( .A(n_92), .B(n_403), .Y(n_402) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_92), .A2(n_456), .B(n_457), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_92), .A2(n_403), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g798 ( .A(n_92), .Y(n_798) );
INVx1_ASAP7_75t_L g196 ( .A(n_94), .Y(n_196) );
XNOR2xp5_ASAP7_75t_L g756 ( .A(n_95), .B(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_96), .B(n_173), .Y(n_520) );
AND2x2_ASAP7_75t_L g242 ( .A(n_97), .B(n_154), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_98), .A2(n_212), .B(n_213), .C(n_215), .Y(n_211) );
INVxp67_ASAP7_75t_L g502 ( .A(n_99), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_100), .B(n_478), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_101), .B(n_173), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_102), .A2(n_477), .B(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g775 ( .A(n_103), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_104), .B(n_146), .Y(n_197) );
AOI21xp33_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_800), .B(n_808), .Y(n_105) );
OA22x2_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_772), .B1(n_775), .B2(n_780), .Y(n_106) );
OAI21xp5_ASAP7_75t_SL g107 ( .A1(n_108), .A2(n_755), .B(n_760), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OAI22xp5_ASAP7_75t_SL g109 ( .A1(n_110), .A2(n_460), .B1(n_469), .B2(n_751), .Y(n_109) );
INVx1_ASAP7_75t_L g762 ( .A(n_110), .Y(n_762) );
NAND3xp33_ASAP7_75t_L g110 ( .A(n_111), .B(n_455), .C(n_458), .Y(n_110) );
NAND4xp25_ASAP7_75t_L g111 ( .A(n_112), .B(n_342), .C(n_402), .D(n_430), .Y(n_111) );
INVx1_ASAP7_75t_L g459 ( .A(n_112), .Y(n_459) );
NAND3x1_ASAP7_75t_L g792 ( .A(n_112), .B(n_342), .C(n_793), .Y(n_792) );
AND3x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_281), .C(n_309), .Y(n_112) );
AOI221x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_204), .B1(n_243), .B2(n_247), .C(n_267), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_175), .B(n_199), .Y(n_115) );
AND2x4_ASAP7_75t_L g351 ( .A(n_116), .B(n_201), .Y(n_351) );
AND2x4_ASAP7_75t_SL g116 ( .A(n_117), .B(n_157), .Y(n_116) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_117), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_117), .B(n_333), .Y(n_450) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g200 ( .A(n_118), .B(n_159), .Y(n_200) );
INVx2_ASAP7_75t_L g274 ( .A(n_118), .Y(n_274) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_118), .Y(n_334) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_118), .Y(n_341) );
AND2x2_ASAP7_75t_L g346 ( .A(n_118), .B(n_158), .Y(n_346) );
INVx1_ASAP7_75t_L g376 ( .A(n_118), .Y(n_376) );
OR2x2_ASAP7_75t_L g429 ( .A(n_118), .B(n_191), .Y(n_429) );
AO21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_153), .Y(n_118) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_119), .A2(n_517), .B(n_523), .Y(n_516) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_119), .A2(n_538), .B(n_544), .Y(n_537) );
AO21x2_ASAP7_75t_L g601 ( .A1(n_119), .A2(n_538), .B(n_544), .Y(n_601) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_120), .A2(n_476), .B(n_482), .Y(n_475) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_SL g121 ( .A(n_122), .B(n_123), .Y(n_121) );
AND2x4_ASAP7_75t_L g161 ( .A(n_122), .B(n_123), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_135), .Y(n_124) );
INVx1_ASAP7_75t_L g224 ( .A(n_126), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_126), .A2(n_136), .B1(n_496), .B2(n_498), .Y(n_495) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_132), .Y(n_126) );
INVx1_ASAP7_75t_L g180 ( .A(n_127), .Y(n_180) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_130), .Y(n_127) );
OR2x6_ASAP7_75t_L g144 ( .A(n_128), .B(n_140), .Y(n_144) );
INVxp33_ASAP7_75t_L g239 ( .A(n_128), .Y(n_239) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g141 ( .A(n_129), .B(n_131), .Y(n_141) );
AND2x4_ASAP7_75t_L g173 ( .A(n_129), .B(n_149), .Y(n_173) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
BUFx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x6_ASAP7_75t_L g477 ( .A(n_133), .B(n_141), .Y(n_477) );
INVx2_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
AND2x6_ASAP7_75t_L g170 ( .A(n_134), .B(n_147), .Y(n_170) );
INVxp67_ASAP7_75t_L g222 ( .A(n_136), .Y(n_222) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
NOR2x1p5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
INVx1_ASAP7_75t_L g240 ( .A(n_139), .Y(n_240) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
O2A1O1Ixp33_ASAP7_75t_SL g142 ( .A1(n_143), .A2(n_144), .B(n_145), .C(n_151), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g163 ( .A1(n_144), .A2(n_164), .B1(n_165), .B2(n_166), .Y(n_163) );
INVx2_ASAP7_75t_L g187 ( .A(n_144), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_144), .A2(n_151), .B(n_196), .C(n_197), .Y(n_195) );
INVxp67_ASAP7_75t_L g212 ( .A(n_144), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_SL g228 ( .A1(n_144), .A2(n_151), .B(n_229), .C(n_230), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_144), .A2(n_151), .B(n_259), .C(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g166 ( .A(n_146), .Y(n_166) );
AND2x4_ASAP7_75t_L g478 ( .A(n_146), .B(n_152), .Y(n_478) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_151), .B(n_161), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_151), .A2(n_185), .B(n_186), .Y(n_184) );
INVx1_ASAP7_75t_L g236 ( .A(n_151), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_151), .A2(n_480), .B(n_481), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_151), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_151), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_151), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_151), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_151), .A2(n_555), .B(n_556), .Y(n_554) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_152), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_154), .A2(n_211), .B1(n_216), .B2(n_217), .Y(n_210) );
INVx3_ASAP7_75t_L g217 ( .A(n_154), .Y(n_217) );
INVx4_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_155), .B(n_220), .Y(n_219) );
AOI21x1_ASAP7_75t_L g551 ( .A1(n_155), .A2(n_552), .B(n_558), .Y(n_551) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx4f_ASAP7_75t_L g189 ( .A(n_156), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_157), .B(n_191), .Y(n_356) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x4_ASAP7_75t_L g246 ( .A(n_158), .B(n_177), .Y(n_246) );
AND2x2_ASAP7_75t_L g333 ( .A(n_158), .B(n_203), .Y(n_333) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g304 ( .A(n_159), .Y(n_304) );
NOR2x1_ASAP7_75t_SL g365 ( .A(n_159), .B(n_191), .Y(n_365) );
AND2x2_ASAP7_75t_L g386 ( .A(n_159), .B(n_177), .Y(n_386) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_162), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_161), .A2(n_194), .B(n_198), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_161), .B(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_161), .B(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_161), .B(n_502), .Y(n_501) );
NOR3xp33_ASAP7_75t_L g503 ( .A(n_161), .B(n_166), .C(n_504), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_161), .A2(n_510), .B(n_511), .Y(n_509) );
OAI21xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_167), .B(n_174), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_166), .B(n_214), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B1(n_171), .B2(n_172), .Y(n_167) );
INVxp67_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVxp67_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g382 ( .A(n_175), .B(n_272), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_175), .B(n_411), .Y(n_410) );
AND2x4_ASAP7_75t_SL g175 ( .A(n_176), .B(n_190), .Y(n_175) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g203 ( .A(n_177), .Y(n_203) );
INVx1_ASAP7_75t_L g271 ( .A(n_177), .Y(n_271) );
AND2x2_ASAP7_75t_L g329 ( .A(n_177), .B(n_191), .Y(n_329) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_183), .Y(n_177) );
NOR3xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .C(n_182), .Y(n_179) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_188), .A2(n_234), .B(n_242), .Y(n_233) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_188), .A2(n_234), .B(n_242), .Y(n_280) );
AOI21x1_ASAP7_75t_L g525 ( .A1(n_188), .A2(n_526), .B(n_529), .Y(n_525) );
INVx2_ASAP7_75t_SL g188 ( .A(n_189), .Y(n_188) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_189), .A2(n_227), .B(n_231), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_189), .A2(n_486), .B(n_487), .Y(n_485) );
NOR2x1_ASAP7_75t_L g244 ( .A(n_190), .B(n_245), .Y(n_244) );
AND2x4_ASAP7_75t_L g270 ( .A(n_190), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g308 ( .A(n_190), .B(n_200), .Y(n_308) );
INVx4_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g289 ( .A(n_191), .Y(n_289) );
AND2x4_ASAP7_75t_L g318 ( .A(n_191), .B(n_271), .Y(n_318) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_191), .Y(n_354) );
AND2x2_ASAP7_75t_L g453 ( .A(n_191), .B(n_304), .Y(n_453) );
OR2x6_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
OAI21xp33_ASAP7_75t_SL g451 ( .A1(n_199), .A2(n_452), .B(n_454), .Y(n_451) );
AND2x2_ASAP7_75t_SL g199 ( .A(n_200), .B(n_201), .Y(n_199) );
NOR2xp33_ASAP7_75t_SL g326 ( .A(n_200), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_SL g408 ( .A(n_201), .Y(n_408) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_206), .A2(n_276), .B1(n_317), .B2(n_333), .Y(n_372) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_225), .Y(n_206) );
INVx1_ASAP7_75t_L g427 ( .A(n_207), .Y(n_427) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g369 ( .A(n_208), .B(n_362), .Y(n_369) );
AND2x2_ASAP7_75t_L g407 ( .A(n_208), .B(n_225), .Y(n_407) );
INVx1_ASAP7_75t_L g421 ( .A(n_208), .Y(n_421) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g251 ( .A(n_209), .Y(n_251) );
AND2x4_ASAP7_75t_L g285 ( .A(n_209), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g294 ( .A(n_209), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_209), .B(n_254), .Y(n_324) );
OR2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_218), .Y(n_209) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_217), .A2(n_255), .B(n_261), .Y(n_254) );
AO21x2_ASAP7_75t_L g300 ( .A1(n_217), .A2(n_255), .B(n_261), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_222), .B1(n_223), .B2(n_224), .Y(n_218) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g265 ( .A(n_225), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g305 ( .A(n_225), .B(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g348 ( .A(n_225), .B(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_232), .Y(n_225) );
INVx1_ASAP7_75t_L g263 ( .A(n_226), .Y(n_263) );
INVx2_ASAP7_75t_L g286 ( .A(n_226), .Y(n_286) );
INVx1_ASAP7_75t_L g301 ( .A(n_226), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_226), .B(n_280), .Y(n_325) );
INVxp67_ASAP7_75t_L g381 ( .A(n_226), .Y(n_381) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g250 ( .A(n_233), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g284 ( .A(n_233), .Y(n_284) );
AND2x4_ASAP7_75t_L g400 ( .A(n_233), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_235), .B(n_241), .Y(n_234) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
BUFx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g328 ( .A(n_245), .Y(n_328) );
OAI21xp5_ASAP7_75t_L g438 ( .A1(n_245), .A2(n_439), .B(n_440), .Y(n_438) );
INVx4_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g288 ( .A(n_246), .B(n_289), .Y(n_288) );
NAND2xp33_ASAP7_75t_SL g247 ( .A(n_248), .B(n_264), .Y(n_247) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_252), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g454 ( .A(n_250), .B(n_299), .Y(n_454) );
AND2x2_ASAP7_75t_L g277 ( .A(n_251), .B(n_263), .Y(n_277) );
AND2x2_ASAP7_75t_L g322 ( .A(n_251), .B(n_300), .Y(n_322) );
NOR2xp67_ASAP7_75t_L g349 ( .A(n_251), .B(n_300), .Y(n_349) );
NAND2x1p5_ASAP7_75t_L g252 ( .A(n_253), .B(n_262), .Y(n_252) );
INVx3_ASAP7_75t_L g266 ( .A(n_253), .Y(n_266) );
AND2x4_ASAP7_75t_L g278 ( .A(n_253), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_253), .B(n_294), .Y(n_314) );
INVx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_254), .B(n_280), .Y(n_296) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_254), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_262), .B(n_313), .Y(n_312) );
INVx3_ASAP7_75t_L g358 ( .A(n_262), .Y(n_358) );
BUFx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_266), .B(n_277), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_266), .B(n_334), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_268), .B(n_275), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_269), .A2(n_419), .B(n_420), .Y(n_418) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
AND2x2_ASAP7_75t_L g302 ( .A(n_270), .B(n_303), .Y(n_302) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_270), .Y(n_310) );
AND2x2_ASAP7_75t_L g424 ( .A(n_270), .B(n_425), .Y(n_424) );
NOR3xp33_ASAP7_75t_L g311 ( .A(n_272), .B(n_312), .C(n_314), .Y(n_311) );
INVx1_ASAP7_75t_L g436 ( .A(n_272), .Y(n_436) );
INVx1_ASAP7_75t_L g446 ( .A(n_272), .Y(n_446) );
AND2x2_ASAP7_75t_L g452 ( .A(n_272), .B(n_453), .Y(n_452) );
INVx3_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_273), .Y(n_425) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_276), .B(n_354), .Y(n_432) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx2_ASAP7_75t_L g336 ( .A(n_277), .Y(n_336) );
INVx1_ASAP7_75t_L g335 ( .A(n_278), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_278), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g313 ( .A(n_279), .Y(n_313) );
AND2x2_ASAP7_75t_L g362 ( .A(n_279), .B(n_300), .Y(n_362) );
AND2x2_ASAP7_75t_L g380 ( .A(n_279), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AOI222xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_288), .B1(n_290), .B2(n_302), .C1(n_305), .C2(n_308), .Y(n_281) );
NAND2xp33_ASAP7_75t_SL g282 ( .A(n_283), .B(n_287), .Y(n_282) );
INVx2_ASAP7_75t_SL g370 ( .A(n_283), .Y(n_370) );
NAND2x1_ASAP7_75t_SL g283 ( .A(n_284), .B(n_285), .Y(n_283) );
OR2x2_ASAP7_75t_L g353 ( .A(n_284), .B(n_336), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_284), .B(n_298), .Y(n_439) );
INVx3_ASAP7_75t_L g389 ( .A(n_285), .Y(n_389) );
AND2x2_ASAP7_75t_L g399 ( .A(n_285), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_288), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g378 ( .A(n_289), .Y(n_378) );
NAND2xp33_ASAP7_75t_L g290 ( .A(n_291), .B(n_297), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OAI21xp33_ASAP7_75t_SL g433 ( .A1(n_292), .A2(n_434), .B(n_437), .Y(n_433) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_293), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g298 ( .A(n_294), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NOR2x1_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g401 ( .A(n_300), .Y(n_401) );
AND2x2_ASAP7_75t_L g317 ( .A(n_303), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NOR2x1_ASAP7_75t_L g377 ( .A(n_304), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AOI211xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B(n_315), .C(n_330), .Y(n_309) );
NAND2x1p5_ASAP7_75t_L g321 ( .A(n_313), .B(n_322), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_319), .B1(n_323), .B2(n_326), .Y(n_315) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g419 ( .A(n_318), .B(n_411), .Y(n_419) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_320), .A2(n_375), .B1(n_379), .B2(n_382), .Y(n_374) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g357 ( .A(n_321), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g379 ( .A(n_322), .B(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx2_ASAP7_75t_SL g391 ( .A(n_324), .Y(n_391) );
INVx2_ASAP7_75t_L g422 ( .A(n_325), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AND2x2_ASAP7_75t_L g338 ( .A(n_329), .B(n_339), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_329), .A2(n_364), .B1(n_388), .B2(n_392), .Y(n_387) );
AND2x2_ASAP7_75t_L g413 ( .A(n_329), .B(n_414), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_335), .B1(n_336), .B2(n_337), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_333), .B(n_354), .Y(n_371) );
INVx2_ASAP7_75t_L g397 ( .A(n_333), .Y(n_397) );
BUFx2_ASAP7_75t_L g411 ( .A(n_334), .Y(n_411) );
NOR2xp33_ASAP7_75t_SL g426 ( .A(n_335), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g364 ( .A(n_339), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVxp67_ASAP7_75t_L g456 ( .A(n_342), .Y(n_456) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_366), .Y(n_342) );
AOI21xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_354), .B(n_355), .Y(n_343) );
OAI21xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_347), .B(n_350), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
OAI21xp33_ASAP7_75t_L g350 ( .A1(n_346), .A2(n_351), .B(n_352), .Y(n_350) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI22xp33_ASAP7_75t_SL g423 ( .A1(n_348), .A2(n_424), .B1(n_426), .B2(n_428), .Y(n_423) );
AOI22xp33_ASAP7_75t_SL g368 ( .A1(n_351), .A2(n_369), .B1(n_370), .B2(n_371), .Y(n_368) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g384 ( .A(n_354), .B(n_385), .Y(n_384) );
OR2x6_ASAP7_75t_L g396 ( .A(n_354), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g398 ( .A(n_354), .B(n_386), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B1(n_359), .B2(n_363), .Y(n_355) );
NOR2xp67_ASAP7_75t_SL g360 ( .A(n_358), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g443 ( .A(n_358), .Y(n_443) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g415 ( .A(n_365), .Y(n_415) );
NOR2xp67_ASAP7_75t_L g366 ( .A(n_367), .B(n_373), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_372), .Y(n_367) );
NAND4xp25_ASAP7_75t_L g373 ( .A(n_374), .B(n_383), .C(n_387), .D(n_394), .Y(n_373) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
AND2x2_ASAP7_75t_L g385 ( .A(n_376), .B(n_386), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g416 ( .A(n_380), .B(n_391), .Y(n_416) );
NAND2xp33_ASAP7_75t_SL g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g406 ( .A(n_393), .Y(n_406) );
OAI21xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_398), .B(n_399), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g445 ( .A(n_400), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g793 ( .A(n_404), .B(n_794), .Y(n_793) );
AOI211x1_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_408), .B(n_409), .C(n_417), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_408), .B(n_436), .Y(n_437) );
AOI31xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .A3(n_415), .B(n_416), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_423), .Y(n_417) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_422), .B(n_448), .Y(n_447) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_425), .Y(n_441) );
INVx2_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g457 ( .A(n_430), .Y(n_457) );
AOI21xp33_ASAP7_75t_SL g430 ( .A1(n_431), .A2(n_438), .B(n_442), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g794 ( .A1(n_431), .A2(n_438), .B(n_442), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVxp33_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI211xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B(n_447), .C(n_451), .Y(n_442) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI21x1_ASAP7_75t_L g761 ( .A1(n_460), .A2(n_762), .B(n_763), .Y(n_761) );
CKINVDCx6p67_ASAP7_75t_R g460 ( .A(n_461), .Y(n_460) );
INVx3_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_463), .Y(n_462) );
AND2x6_ASAP7_75t_SL g463 ( .A(n_464), .B(n_465), .Y(n_463) );
OR2x6_ASAP7_75t_SL g753 ( .A(n_464), .B(n_754), .Y(n_753) );
OR2x2_ASAP7_75t_L g771 ( .A(n_464), .B(n_465), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_464), .B(n_754), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g754 ( .A(n_465), .Y(n_754) );
INVx1_ASAP7_75t_L g803 ( .A(n_466), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
NAND2x1_ASAP7_75t_SL g763 ( .A(n_469), .B(n_764), .Y(n_763) );
INVx4_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OR2x6_ASAP7_75t_L g470 ( .A(n_471), .B(n_664), .Y(n_470) );
NAND3xp33_ASAP7_75t_SL g471 ( .A(n_472), .B(n_574), .C(n_614), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_492), .B(n_505), .C(n_530), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_473), .B(n_579), .Y(n_613) );
NOR2x1p5_ASAP7_75t_L g473 ( .A(n_474), .B(n_483), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g549 ( .A(n_475), .Y(n_549) );
INVx2_ASAP7_75t_L g565 ( .A(n_475), .Y(n_565) );
OR2x2_ASAP7_75t_L g577 ( .A(n_475), .B(n_484), .Y(n_577) );
AND2x2_ASAP7_75t_L g591 ( .A(n_475), .B(n_550), .Y(n_591) );
INVx1_ASAP7_75t_L g619 ( .A(n_475), .Y(n_619) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_475), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_475), .B(n_484), .Y(n_725) );
OR2x2_ASAP7_75t_L g546 ( .A(n_483), .B(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_483), .Y(n_681) );
AND2x2_ASAP7_75t_L g686 ( .A(n_483), .B(n_548), .Y(n_686) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x4_ASAP7_75t_L g492 ( .A(n_484), .B(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g545 ( .A(n_484), .B(n_494), .Y(n_545) );
OR2x2_ASAP7_75t_L g564 ( .A(n_484), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g593 ( .A(n_484), .Y(n_593) );
AND2x4_ASAP7_75t_SL g632 ( .A(n_484), .B(n_494), .Y(n_632) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_484), .Y(n_636) );
OR2x2_ASAP7_75t_L g653 ( .A(n_484), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g663 ( .A(n_484), .B(n_570), .Y(n_663) );
INVx1_ASAP7_75t_L g692 ( .A(n_484), .Y(n_692) );
OR2x6_ASAP7_75t_L g484 ( .A(n_485), .B(n_491), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_492), .B(n_621), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_493), .B(n_550), .Y(n_567) );
AND2x2_ASAP7_75t_L g579 ( .A(n_493), .B(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g597 ( .A(n_493), .B(n_564), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_493), .B(n_618), .Y(n_617) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x4_ASAP7_75t_L g570 ( .A(n_494), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g592 ( .A(n_494), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g627 ( .A(n_494), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_494), .B(n_550), .Y(n_651) );
AND2x4_ASAP7_75t_L g494 ( .A(n_495), .B(n_500), .Y(n_494) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_515), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_506), .B(n_583), .Y(n_582) );
AND2x4_ASAP7_75t_L g600 ( .A(n_506), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_506), .B(n_516), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g620 ( .A(n_506), .B(n_621), .C(n_622), .Y(n_620) );
AND2x2_ASAP7_75t_L g668 ( .A(n_506), .B(n_573), .Y(n_668) );
INVx5_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g535 ( .A(n_507), .B(n_536), .Y(n_535) );
AND2x4_ASAP7_75t_SL g572 ( .A(n_507), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g588 ( .A(n_507), .Y(n_588) );
OR2x2_ASAP7_75t_L g611 ( .A(n_507), .B(n_601), .Y(n_611) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_507), .Y(n_628) );
AND2x2_ASAP7_75t_SL g646 ( .A(n_507), .B(n_534), .Y(n_646) );
AND2x4_ASAP7_75t_L g661 ( .A(n_507), .B(n_537), .Y(n_661) );
AND2x2_ASAP7_75t_L g675 ( .A(n_507), .B(n_516), .Y(n_675) );
OR2x2_ASAP7_75t_L g696 ( .A(n_507), .B(n_524), .Y(n_696) );
OR2x6_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
AND2x2_ASAP7_75t_L g750 ( .A(n_515), .B(n_628), .Y(n_750) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_524), .Y(n_515) );
AND2x4_ASAP7_75t_L g573 ( .A(n_516), .B(n_536), .Y(n_573) );
INVx2_ASAP7_75t_L g584 ( .A(n_516), .Y(n_584) );
AND2x2_ASAP7_75t_L g589 ( .A(n_516), .B(n_534), .Y(n_589) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_516), .Y(n_622) );
OR2x2_ASAP7_75t_L g645 ( .A(n_516), .B(n_537), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_516), .B(n_537), .Y(n_648) );
INVx1_ASAP7_75t_L g657 ( .A(n_516), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_522), .Y(n_517) );
AND2x2_ASAP7_75t_L g560 ( .A(n_524), .B(n_537), .Y(n_560) );
BUFx2_ASAP7_75t_L g609 ( .A(n_524), .Y(n_609) );
AND2x2_ASAP7_75t_L g704 ( .A(n_524), .B(n_584), .Y(n_704) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_525), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
OAI221xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_545), .B1(n_546), .B2(n_559), .C(n_561), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
NOR2x1_ASAP7_75t_L g606 ( .A(n_533), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_533), .B(n_600), .Y(n_640) );
OR2x2_ASAP7_75t_L g652 ( .A(n_533), .B(n_648), .Y(n_652) );
OR2x2_ASAP7_75t_L g655 ( .A(n_533), .B(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g744 ( .A(n_533), .B(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x4_ASAP7_75t_L g583 ( .A(n_534), .B(n_584), .Y(n_583) );
OA33x2_ASAP7_75t_L g616 ( .A1(n_534), .A2(n_577), .A3(n_617), .B1(n_620), .B2(n_623), .B3(n_626), .Y(n_616) );
OR2x2_ASAP7_75t_L g647 ( .A(n_534), .B(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g671 ( .A(n_534), .B(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g679 ( .A(n_534), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g699 ( .A(n_534), .B(n_573), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_534), .B(n_588), .Y(n_737) );
INVx2_ASAP7_75t_L g607 ( .A(n_535), .Y(n_607) );
AOI322xp5_ASAP7_75t_L g677 ( .A1(n_535), .A2(n_590), .A3(n_678), .B1(n_681), .B2(n_682), .C1(n_684), .C2(n_686), .Y(n_677) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_537), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_543), .Y(n_538) );
OR2x2_ASAP7_75t_L g659 ( .A(n_545), .B(n_638), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_545), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g732 ( .A(n_545), .Y(n_732) );
INVx1_ASAP7_75t_SL g598 ( .A(n_546), .Y(n_598) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g631 ( .A(n_548), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
INVx2_ASAP7_75t_L g571 ( .A(n_550), .Y(n_571) );
INVx1_ASAP7_75t_L g580 ( .A(n_550), .Y(n_580) );
INVx1_ASAP7_75t_L g621 ( .A(n_550), .Y(n_621) );
OR2x2_ASAP7_75t_L g638 ( .A(n_550), .B(n_565), .Y(n_638) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_550), .Y(n_713) );
INVx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_557), .Y(n_552) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_SL g682 ( .A(n_560), .B(n_683), .Y(n_682) );
OAI21xp5_ASAP7_75t_SL g561 ( .A1(n_562), .A2(n_568), .B(n_572), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g635 ( .A1(n_562), .A2(n_636), .B(n_637), .C(n_639), .Y(n_635) );
AND2x4_ASAP7_75t_L g562 ( .A(n_563), .B(n_566), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g700 ( .A(n_564), .B(n_701), .Y(n_700) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_565), .Y(n_569) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g724 ( .A(n_567), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AND2x2_ASAP7_75t_SL g693 ( .A(n_570), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g701 ( .A(n_570), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_570), .B(n_692), .Y(n_709) );
INVx3_ASAP7_75t_SL g634 ( .A(n_573), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_581), .B1(n_585), .B2(n_590), .C(n_594), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_580), .Y(n_625) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_583), .A2(n_610), .B(n_682), .Y(n_688) );
AND2x2_ASAP7_75t_L g714 ( .A(n_583), .B(n_661), .Y(n_714) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_584), .Y(n_602) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_588), .B(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g723 ( .A(n_588), .B(n_645), .Y(n_723) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx2_ASAP7_75t_L g672 ( .A(n_591), .Y(n_672) );
OAI21xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_599), .B(n_603), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
INVx2_ASAP7_75t_L g745 ( .A(n_600), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_601), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g674 ( .A(n_601), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_602), .B(n_624), .Y(n_623) );
OAI31xp33_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_606), .A3(n_608), .B(n_612), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_607), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
OR2x2_ASAP7_75t_L g685 ( .A(n_609), .B(n_611), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_609), .B(n_661), .Y(n_740) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NOR5xp2_ASAP7_75t_L g614 ( .A(n_615), .B(n_629), .C(n_641), .D(n_650), .E(n_658), .Y(n_614) );
INVxp67_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_619), .B(n_621), .Y(n_654) );
INVx1_ASAP7_75t_L g694 ( .A(n_619), .Y(n_694) );
INVxp67_ASAP7_75t_SL g731 ( .A(n_619), .Y(n_731) );
INVx1_ASAP7_75t_L g683 ( .A(n_622), .Y(n_683) );
INVxp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp33_ASAP7_75t_SL g626 ( .A(n_627), .B(n_628), .Y(n_626) );
OAI321xp33_ASAP7_75t_L g666 ( .A1(n_627), .A2(n_667), .A3(n_669), .B1(n_673), .B2(n_676), .C(n_677), .Y(n_666) );
INVx1_ASAP7_75t_L g720 ( .A(n_628), .Y(n_720) );
OAI21xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_633), .B(n_635), .Y(n_629) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_631), .A2(n_704), .B1(n_711), .B2(n_714), .Y(n_710) );
AND2x2_ASAP7_75t_L g739 ( .A(n_632), .B(n_713), .Y(n_739) );
INVx1_ASAP7_75t_L g649 ( .A(n_637), .Y(n_649) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_647), .B(n_649), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_648), .A2(n_659), .B1(n_660), .B2(n_662), .Y(n_658) );
INVx1_ASAP7_75t_L g721 ( .A(n_648), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B1(n_653), .B2(n_655), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_657), .B(n_661), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g735 ( .A1(n_659), .A2(n_736), .B1(n_738), .B2(n_740), .C(n_741), .Y(n_735) );
INVx1_ASAP7_75t_L g742 ( .A(n_659), .Y(n_742) );
OAI221xp5_ASAP7_75t_L g716 ( .A1(n_660), .A2(n_717), .B1(n_724), .B2(n_726), .C(n_727), .Y(n_716) );
OAI21xp5_ASAP7_75t_L g687 ( .A1(n_662), .A2(n_688), .B(n_689), .Y(n_687) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_715), .Y(n_664) );
NOR3xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_687), .C(n_705), .Y(n_665) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_668), .Y(n_734) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx3_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g733 ( .A(n_676), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_678), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g726 ( .A(n_686), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_695), .B(n_697), .Y(n_689) );
INVxp67_ASAP7_75t_L g747 ( .A(n_690), .Y(n_747) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_SL g702 ( .A(n_693), .Y(n_702) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_700), .B1(n_702), .B2(n_703), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI21xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B(n_710), .Y(n_705) );
INVx1_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g748 ( .A(n_711), .Y(n_748) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_735), .C(n_746), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_718), .B(n_722), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI21xp5_ASAP7_75t_SL g727 ( .A1(n_728), .A2(n_733), .B(n_734), .Y(n_727) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI21xp5_ASAP7_75t_L g741 ( .A1(n_739), .A2(n_742), .B(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI21xp33_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_748), .B(n_749), .Y(n_746) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_752), .Y(n_766) );
CKINVDCx11_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
AOI21xp33_ASAP7_75t_SL g760 ( .A1(n_755), .A2(n_761), .B(n_767), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_765), .Y(n_764) );
BUFx4f_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
INVx1_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_776), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_774), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_775), .Y(n_774) );
OAI21xp5_ASAP7_75t_L g780 ( .A1(n_776), .A2(n_781), .B(n_783), .Y(n_780) );
INVx1_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
BUFx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
BUFx2_ASAP7_75t_R g782 ( .A(n_779), .Y(n_782) );
INVx1_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_785), .B1(n_791), .B2(n_799), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g799 ( .A(n_791), .Y(n_799) );
XOR2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_795), .Y(n_791) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
INVx3_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_SL g810 ( .A(n_801), .Y(n_810) );
INVx2_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
AND2x2_ASAP7_75t_SL g802 ( .A(n_803), .B(n_804), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
endmodule