module fake_aes_847_n_1469 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_241, n_95, n_238, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1469, n_667);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_241;
input n_95;
input n_238;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1469;
output n_667;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_315;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1408;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_1455;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_1459;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_322;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1454;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_584;
wire n_1130;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1439;
wire n_374;
wire n_718;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_325;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g314 ( .A(n_129), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_106), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_246), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_121), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_7), .Y(n_318) );
CKINVDCx16_ASAP7_75t_R g319 ( .A(n_172), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_178), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_138), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_0), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_290), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_220), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_223), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_284), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_254), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_149), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_304), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_168), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_45), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_162), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_283), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_243), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_5), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_94), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_57), .Y(n_337) );
CKINVDCx16_ASAP7_75t_R g338 ( .A(n_111), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_80), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_221), .Y(n_340) );
INVxp33_ASAP7_75t_SL g341 ( .A(n_84), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_114), .Y(n_342) );
CKINVDCx16_ASAP7_75t_R g343 ( .A(n_171), .Y(n_343) );
CKINVDCx16_ASAP7_75t_R g344 ( .A(n_233), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_75), .Y(n_345) );
BUFx2_ASAP7_75t_SL g346 ( .A(n_26), .Y(n_346) );
INVxp67_ASAP7_75t_L g347 ( .A(n_197), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_292), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_130), .Y(n_349) );
INVxp33_ASAP7_75t_L g350 ( .A(n_161), .Y(n_350) );
INVx1_ASAP7_75t_SL g351 ( .A(n_95), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_101), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_18), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_270), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_182), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_288), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_303), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_14), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_309), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_188), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_107), .Y(n_361) );
INVxp33_ASAP7_75t_SL g362 ( .A(n_78), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_238), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_263), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_122), .Y(n_365) );
BUFx2_ASAP7_75t_SL g366 ( .A(n_192), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_208), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_286), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_159), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_40), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_287), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_126), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_224), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_251), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_84), .Y(n_375) );
CKINVDCx16_ASAP7_75t_R g376 ( .A(n_183), .Y(n_376) );
INVxp33_ASAP7_75t_L g377 ( .A(n_22), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_143), .Y(n_378) );
INVxp33_ASAP7_75t_L g379 ( .A(n_173), .Y(n_379) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_242), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_185), .Y(n_381) );
CKINVDCx20_ASAP7_75t_R g382 ( .A(n_256), .Y(n_382) );
INVxp33_ASAP7_75t_SL g383 ( .A(n_40), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_234), .Y(n_384) );
INVx2_ASAP7_75t_SL g385 ( .A(n_268), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_216), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_235), .Y(n_387) );
NOR2xp67_ASAP7_75t_L g388 ( .A(n_82), .B(n_313), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_24), .Y(n_389) );
INVxp33_ASAP7_75t_SL g390 ( .A(n_3), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_97), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_170), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_217), .Y(n_393) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_190), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_112), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_261), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_75), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_39), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_181), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_44), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_0), .Y(n_401) );
CKINVDCx16_ASAP7_75t_R g402 ( .A(n_43), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_123), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_310), .Y(n_404) );
INVxp33_ASAP7_75t_SL g405 ( .A(n_237), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_218), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_109), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_29), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_15), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_47), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_210), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_275), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_29), .B(n_110), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_6), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_239), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_305), .B(n_26), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_108), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_244), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_148), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_100), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_133), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_164), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_226), .Y(n_423) );
INVxp33_ASAP7_75t_L g424 ( .A(n_265), .Y(n_424) );
INVxp67_ASAP7_75t_SL g425 ( .A(n_291), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_6), .B(n_176), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_3), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_82), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_120), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_53), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_262), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_140), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_60), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_124), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_93), .Y(n_435) );
CKINVDCx16_ASAP7_75t_R g436 ( .A(n_45), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_204), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_266), .Y(n_438) );
CKINVDCx14_ASAP7_75t_R g439 ( .A(n_184), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_74), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_228), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_90), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_56), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_306), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_8), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_195), .Y(n_446) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_128), .Y(n_447) );
INVxp33_ASAP7_75t_L g448 ( .A(n_255), .Y(n_448) );
INVxp67_ASAP7_75t_SL g449 ( .A(n_206), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_47), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_139), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_58), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_89), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_10), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_245), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_213), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_293), .Y(n_457) );
INVxp67_ASAP7_75t_L g458 ( .A(n_35), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_36), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_21), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_127), .Y(n_461) );
CKINVDCx14_ASAP7_75t_R g462 ( .A(n_10), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_125), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_116), .Y(n_464) );
INVxp67_ASAP7_75t_SL g465 ( .A(n_25), .Y(n_465) );
INVxp67_ASAP7_75t_SL g466 ( .A(n_118), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_285), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_282), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_46), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_193), .Y(n_470) );
INVxp67_ASAP7_75t_SL g471 ( .A(n_264), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_56), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_215), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_232), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_160), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_231), .Y(n_476) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_374), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_400), .Y(n_478) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_374), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_377), .B(n_1), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_400), .Y(n_481) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_374), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_462), .Y(n_483) );
OAI22xp5_ASAP7_75t_SL g484 ( .A1(n_443), .A2(n_436), .B1(n_402), .B2(n_341), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_341), .A2(n_4), .B1(n_1), .B2(n_2), .Y(n_485) );
AND2x4_ASAP7_75t_L g486 ( .A(n_385), .B(n_2), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_385), .B(n_4), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_314), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_321), .Y(n_489) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_374), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_321), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_318), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_323), .B(n_5), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_332), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_323), .B(n_7), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_315), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_319), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_377), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_316), .Y(n_499) );
BUFx2_ASAP7_75t_L g500 ( .A(n_335), .Y(n_500) );
NAND2xp33_ASAP7_75t_L g501 ( .A(n_350), .B(n_91), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_320), .Y(n_502) );
BUFx8_ASAP7_75t_L g503 ( .A(n_426), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_352), .B(n_8), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_326), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_327), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_328), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_338), .Y(n_508) );
INVx3_ASAP7_75t_L g509 ( .A(n_332), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_443), .Y(n_510) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_374), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_342), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_330), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_333), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_477), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_488), .B(n_324), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_480), .A2(n_383), .B1(n_390), .B2(n_362), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_498), .B(n_350), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_500), .Y(n_519) );
NAND3xp33_ASAP7_75t_L g520 ( .A(n_488), .B(n_340), .C(n_336), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_500), .B(n_379), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_496), .B(n_379), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_509), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_503), .B(n_343), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_503), .B(n_344), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_486), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_496), .B(n_424), .Y(n_527) );
BUFx3_ASAP7_75t_L g528 ( .A(n_486), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_509), .Y(n_529) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_477), .Y(n_530) );
BUFx4f_ASAP7_75t_L g531 ( .A(n_493), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_480), .A2(n_322), .B1(n_337), .B2(n_331), .Y(n_532) );
INVx3_ASAP7_75t_L g533 ( .A(n_486), .Y(n_533) );
BUFx3_ASAP7_75t_L g534 ( .A(n_486), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_492), .B(n_424), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_497), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_499), .B(n_325), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_508), .B(n_335), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_509), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_499), .B(n_448), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_503), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_502), .B(n_505), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_477), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_503), .B(n_376), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_502), .B(n_505), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_506), .B(n_448), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_506), .B(n_358), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_507), .B(n_439), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_484), .A2(n_362), .B1(n_390), .B2(n_383), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_507), .B(n_437), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_487), .B(n_329), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g552 ( .A(n_513), .B(n_355), .C(n_348), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_477), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_477), .Y(n_554) );
INVx3_ASAP7_75t_L g555 ( .A(n_487), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_513), .B(n_334), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_483), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_514), .B(n_358), .Y(n_558) );
INVx6_ASAP7_75t_L g559 ( .A(n_493), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_510), .Y(n_560) );
INVx6_ASAP7_75t_L g561 ( .A(n_493), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_509), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_489), .Y(n_563) );
O2A1O1Ixp33_ASAP7_75t_L g564 ( .A1(n_547), .A2(n_514), .B(n_501), .C(n_458), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_558), .B(n_487), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_542), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_542), .Y(n_567) );
NAND2x1p5_ASAP7_75t_L g568 ( .A(n_541), .B(n_487), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_528), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_531), .B(n_493), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_563), .Y(n_571) );
BUFx3_ASAP7_75t_L g572 ( .A(n_541), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_535), .B(n_495), .Y(n_573) );
BUFx2_ASAP7_75t_L g574 ( .A(n_519), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_518), .B(n_397), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_535), .B(n_495), .Y(n_576) );
NOR3xp33_ASAP7_75t_SL g577 ( .A(n_536), .B(n_408), .C(n_397), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_521), .A2(n_504), .B1(n_495), .B2(n_382), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_522), .B(n_495), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_528), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_531), .A2(n_504), .B1(n_491), .B2(n_494), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_563), .Y(n_582) );
AND2x4_ASAP7_75t_L g583 ( .A(n_548), .B(n_504), .Y(n_583) );
AND2x4_ASAP7_75t_L g584 ( .A(n_548), .B(n_504), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_523), .Y(n_585) );
INVx4_ASAP7_75t_L g586 ( .A(n_531), .Y(n_586) );
NOR2x2_ASAP7_75t_L g587 ( .A(n_560), .B(n_382), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_527), .B(n_329), .Y(n_588) );
AND2x4_ASAP7_75t_L g589 ( .A(n_524), .B(n_485), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_560), .Y(n_590) );
AOI22xp33_ASAP7_75t_SL g591 ( .A1(n_559), .A2(n_346), .B1(n_421), .B2(n_415), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_531), .A2(n_491), .B(n_489), .Y(n_592) );
NAND3xp33_ASAP7_75t_SL g593 ( .A(n_532), .B(n_485), .C(n_409), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_523), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_518), .A2(n_421), .B1(n_431), .B2(n_415), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_529), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_551), .B(n_405), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_529), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_517), .A2(n_431), .B1(n_408), .B2(n_430), .Y(n_599) );
NOR3xp33_ASAP7_75t_SL g600 ( .A(n_525), .B(n_430), .C(n_409), .Y(n_600) );
INVxp67_ASAP7_75t_L g601 ( .A(n_547), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_550), .B(n_440), .Y(n_602) );
BUFx12f_ASAP7_75t_L g603 ( .A(n_538), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_539), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_540), .B(n_349), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_539), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_550), .B(n_405), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_546), .B(n_349), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_528), .Y(n_609) );
INVx5_ASAP7_75t_L g610 ( .A(n_559), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_534), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_534), .Y(n_612) );
BUFx3_ASAP7_75t_L g613 ( .A(n_534), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_562), .Y(n_614) );
INVx3_ASAP7_75t_L g615 ( .A(n_559), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_516), .B(n_354), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_516), .B(n_354), .Y(n_617) );
BUFx2_ASAP7_75t_L g618 ( .A(n_538), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_526), .B(n_357), .Y(n_619) );
INVxp67_ASAP7_75t_L g620 ( .A(n_537), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_559), .Y(n_621) );
NOR2x1p5_ASAP7_75t_L g622 ( .A(n_537), .B(n_440), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_544), .Y(n_623) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_559), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_517), .A2(n_445), .B1(n_472), .B2(n_465), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_556), .B(n_356), .Y(n_626) );
INVx2_ASAP7_75t_SL g627 ( .A(n_561), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_562), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_561), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_545), .B(n_356), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_561), .A2(n_445), .B1(n_472), .B2(n_426), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_526), .B(n_369), .Y(n_632) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_561), .Y(n_633) );
BUFx2_ASAP7_75t_L g634 ( .A(n_557), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_526), .B(n_359), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g636 ( .A1(n_526), .A2(n_361), .B(n_360), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_561), .Y(n_637) );
INVx3_ASAP7_75t_L g638 ( .A(n_533), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_533), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_549), .A2(n_339), .B1(n_353), .B2(n_345), .Y(n_640) );
OAI22xp5_ASAP7_75t_SL g641 ( .A1(n_549), .A2(n_370), .B1(n_389), .B2(n_375), .Y(n_641) );
BUFx3_ASAP7_75t_L g642 ( .A(n_555), .Y(n_642) );
INVx3_ASAP7_75t_L g643 ( .A(n_533), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_520), .B(n_478), .Y(n_644) );
INVx4_ASAP7_75t_L g645 ( .A(n_555), .Y(n_645) );
BUFx12f_ASAP7_75t_L g646 ( .A(n_530), .Y(n_646) );
AND2x4_ASAP7_75t_L g647 ( .A(n_555), .B(n_478), .Y(n_647) );
BUFx3_ASAP7_75t_L g648 ( .A(n_555), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_520), .B(n_369), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_552), .B(n_373), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_552), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_554), .B(n_481), .Y(n_652) );
AND2x4_ASAP7_75t_SL g653 ( .A(n_554), .B(n_398), .Y(n_653) );
INVx1_ASAP7_75t_SL g654 ( .A(n_515), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_515), .B(n_365), .Y(n_655) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_515), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_543), .Y(n_657) );
A2O1A1Ixp33_ASAP7_75t_L g658 ( .A1(n_543), .A2(n_481), .B(n_512), .C(n_494), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_553), .B(n_367), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_638), .Y(n_660) );
INVx3_ASAP7_75t_SL g661 ( .A(n_587), .Y(n_661) );
O2A1O1Ixp33_ASAP7_75t_L g662 ( .A1(n_566), .A2(n_410), .B(n_414), .C(n_401), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_638), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_620), .B(n_427), .Y(n_664) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_572), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_643), .Y(n_666) );
UNKNOWN g667 ( );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_589), .A2(n_428), .B1(n_442), .B2(n_433), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_620), .B(n_601), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_567), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_643), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_589), .A2(n_450), .B1(n_453), .B2(n_452), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_642), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_647), .Y(n_674) );
BUFx3_ASAP7_75t_L g675 ( .A(n_634), .Y(n_675) );
INVx1_ASAP7_75t_SL g676 ( .A(n_574), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_572), .B(n_412), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_642), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_570), .A2(n_416), .B(n_413), .Y(n_679) );
BUFx3_ASAP7_75t_L g680 ( .A(n_603), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_590), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g682 ( .A1(n_601), .A2(n_459), .B(n_460), .C(n_454), .Y(n_682) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_618), .Y(n_683) );
INVx4_ASAP7_75t_L g684 ( .A(n_586), .Y(n_684) );
BUFx3_ASAP7_75t_L g685 ( .A(n_623), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_570), .A2(n_425), .B(n_380), .Y(n_686) );
O2A1O1Ixp33_ASAP7_75t_L g687 ( .A1(n_573), .A2(n_469), .B(n_512), .C(n_368), .Y(n_687) );
BUFx3_ASAP7_75t_L g688 ( .A(n_624), .Y(n_688) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_646), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_607), .B(n_412), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_586), .B(n_417), .Y(n_691) );
AOI21xp33_ASAP7_75t_L g692 ( .A1(n_565), .A2(n_466), .B(n_449), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_607), .B(n_347), .Y(n_693) );
AO22x1_ASAP7_75t_L g694 ( .A1(n_587), .A2(n_447), .B1(n_451), .B2(n_417), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_647), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_583), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_583), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_584), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_581), .A2(n_471), .B1(n_388), .B2(n_371), .Y(n_699) );
OR2x6_ASAP7_75t_L g700 ( .A(n_584), .B(n_366), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_575), .B(n_447), .Y(n_701) );
INVx3_ASAP7_75t_L g702 ( .A(n_624), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_565), .B(n_451), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_648), .Y(n_704) );
INVxp67_ASAP7_75t_SL g705 ( .A(n_613), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_585), .Y(n_706) );
AOI21xp33_ASAP7_75t_L g707 ( .A1(n_564), .A2(n_381), .B(n_372), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_594), .Y(n_708) );
CKINVDCx5p33_ASAP7_75t_R g709 ( .A(n_591), .Y(n_709) );
BUFx5_ASAP7_75t_L g710 ( .A(n_613), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_619), .A2(n_387), .B(n_386), .Y(n_711) );
INVx3_ASAP7_75t_L g712 ( .A(n_624), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_602), .B(n_457), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_596), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_598), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_604), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_606), .Y(n_717) );
AND2x4_ASAP7_75t_L g718 ( .A(n_622), .B(n_391), .Y(n_718) );
BUFx12f_ASAP7_75t_L g719 ( .A(n_568), .Y(n_719) );
CKINVDCx5p33_ASAP7_75t_R g720 ( .A(n_591), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_614), .Y(n_721) );
BUFx2_ASAP7_75t_SL g722 ( .A(n_595), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_628), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_624), .Y(n_724) );
INVx4_ASAP7_75t_L g725 ( .A(n_610), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_593), .B(n_457), .Y(n_726) );
BUFx3_ASAP7_75t_L g727 ( .A(n_633), .Y(n_727) );
INVx4_ASAP7_75t_L g728 ( .A(n_610), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_619), .A2(n_395), .B(n_393), .Y(n_729) );
AOI221xp5_ASAP7_75t_L g730 ( .A1(n_593), .A2(n_463), .B1(n_473), .B2(n_403), .C(n_404), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_615), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_576), .B(n_463), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_615), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_635), .A2(n_406), .B(n_396), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_571), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_625), .B(n_473), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_633), .Y(n_737) );
INVx2_ASAP7_75t_SL g738 ( .A(n_616), .Y(n_738) );
CKINVDCx8_ASAP7_75t_R g739 ( .A(n_597), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_582), .Y(n_740) );
BUFx6f_ASAP7_75t_L g741 ( .A(n_633), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_579), .B(n_407), .Y(n_742) );
BUFx6f_ASAP7_75t_L g743 ( .A(n_633), .Y(n_743) );
INVx2_ASAP7_75t_SL g744 ( .A(n_617), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_629), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g746 ( .A1(n_651), .A2(n_418), .B(n_419), .C(n_411), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_645), .B(n_420), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_621), .Y(n_748) );
O2A1O1Ixp33_ASAP7_75t_SL g749 ( .A1(n_658), .A2(n_429), .B(n_432), .C(n_422), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_578), .A2(n_435), .B1(n_438), .B2(n_434), .Y(n_750) );
A2O1A1Ixp33_ASAP7_75t_L g751 ( .A1(n_636), .A2(n_444), .B(n_446), .C(n_441), .Y(n_751) );
BUFx6f_ASAP7_75t_L g752 ( .A(n_610), .Y(n_752) );
BUFx8_ASAP7_75t_L g753 ( .A(n_644), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_635), .A2(n_456), .B(n_455), .Y(n_754) );
INVx3_ASAP7_75t_L g755 ( .A(n_610), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_639), .A2(n_464), .B(n_461), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_645), .B(n_467), .Y(n_757) );
NOR2xp33_ASAP7_75t_SL g758 ( .A(n_568), .B(n_352), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_597), .B(n_317), .Y(n_759) );
BUFx3_ASAP7_75t_L g760 ( .A(n_652), .Y(n_760) );
BUFx6f_ASAP7_75t_L g761 ( .A(n_627), .Y(n_761) );
INVx3_ASAP7_75t_L g762 ( .A(n_569), .Y(n_762) );
A2O1A1Ixp33_ASAP7_75t_SL g763 ( .A1(n_652), .A2(n_554), .B(n_553), .C(n_363), .Y(n_763) );
CKINVDCx5p33_ASAP7_75t_R g764 ( .A(n_577), .Y(n_764) );
AOI222xp33_ASAP7_75t_L g765 ( .A1(n_641), .A2(n_468), .B1(n_470), .B2(n_351), .C1(n_423), .C2(n_364), .Y(n_765) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_653), .Y(n_766) );
AND2x4_ASAP7_75t_L g767 ( .A(n_600), .B(n_364), .Y(n_767) );
A2O1A1Ixp33_ASAP7_75t_L g768 ( .A1(n_592), .A2(n_363), .B(n_378), .C(n_342), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_637), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_632), .A2(n_384), .B(n_378), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_581), .A2(n_392), .B1(n_474), .B2(n_384), .Y(n_771) );
INVx3_ASAP7_75t_L g772 ( .A(n_580), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_609), .Y(n_773) );
INVx1_ASAP7_75t_SL g774 ( .A(n_653), .Y(n_774) );
BUFx6f_ASAP7_75t_L g775 ( .A(n_611), .Y(n_775) );
BUFx8_ASAP7_75t_SL g776 ( .A(n_649), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_612), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_631), .B(n_475), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_626), .B(n_9), .Y(n_779) );
BUFx3_ASAP7_75t_L g780 ( .A(n_640), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_658), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_656), .Y(n_782) );
NAND2xp5_ASAP7_75t_SL g783 ( .A(n_630), .B(n_475), .Y(n_783) );
INVx3_ASAP7_75t_L g784 ( .A(n_654), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_588), .B(n_9), .Y(n_785) );
BUFx2_ASAP7_75t_L g786 ( .A(n_600), .Y(n_786) );
BUFx3_ASAP7_75t_L g787 ( .A(n_650), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_656), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_577), .B(n_11), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_605), .A2(n_476), .B1(n_399), .B2(n_394), .Y(n_790) );
OAI22x1_ASAP7_75t_L g791 ( .A1(n_608), .A2(n_476), .B1(n_13), .B2(n_11), .Y(n_791) );
BUFx2_ASAP7_75t_L g792 ( .A(n_657), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_655), .A2(n_399), .B1(n_394), .B2(n_477), .Y(n_793) );
INVx3_ASAP7_75t_L g794 ( .A(n_659), .Y(n_794) );
INVxp67_ASAP7_75t_SL g795 ( .A(n_659), .Y(n_795) );
BUFx3_ASAP7_75t_L g796 ( .A(n_634), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_566), .Y(n_797) );
INVx2_ASAP7_75t_SL g798 ( .A(n_574), .Y(n_798) );
AND2x4_ASAP7_75t_L g799 ( .A(n_620), .B(n_12), .Y(n_799) );
INVx1_ASAP7_75t_SL g800 ( .A(n_574), .Y(n_800) );
INVx3_ASAP7_75t_L g801 ( .A(n_624), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_566), .Y(n_802) );
NAND2xp5_ASAP7_75t_SL g803 ( .A(n_572), .B(n_394), .Y(n_803) );
BUFx6f_ASAP7_75t_L g804 ( .A(n_572), .Y(n_804) );
OAI21x1_ASAP7_75t_L g805 ( .A1(n_770), .A2(n_553), .B(n_399), .Y(n_805) );
CKINVDCx11_ASAP7_75t_R g806 ( .A(n_680), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_675), .Y(n_807) );
BUFx6f_ASAP7_75t_L g808 ( .A(n_689), .Y(n_808) );
AND2x4_ASAP7_75t_L g809 ( .A(n_670), .B(n_13), .Y(n_809) );
AOI21x1_ASAP7_75t_L g810 ( .A1(n_770), .A2(n_399), .B(n_394), .Y(n_810) );
INVx4_ASAP7_75t_L g811 ( .A(n_689), .Y(n_811) );
INVxp67_ASAP7_75t_SL g812 ( .A(n_799), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_797), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_799), .A2(n_482), .B1(n_490), .B2(n_479), .Y(n_814) );
BUFx6f_ASAP7_75t_L g815 ( .A(n_689), .Y(n_815) );
AND2x4_ASAP7_75t_L g816 ( .A(n_802), .B(n_14), .Y(n_816) );
INVx3_ASAP7_75t_L g817 ( .A(n_684), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_774), .A2(n_482), .B1(n_490), .B2(n_479), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_669), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_782), .Y(n_820) );
AND2x4_ASAP7_75t_L g821 ( .A(n_738), .B(n_15), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_706), .B(n_16), .Y(n_822) );
AND2x2_ASAP7_75t_SL g823 ( .A(n_758), .B(n_16), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_788), .Y(n_824) );
OR2x6_ASAP7_75t_L g825 ( .A(n_719), .B(n_17), .Y(n_825) );
OAI21x1_ASAP7_75t_L g826 ( .A1(n_803), .A2(n_490), .B(n_482), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_735), .Y(n_827) );
BUFx3_ASAP7_75t_L g828 ( .A(n_796), .Y(n_828) );
NAND2x1p5_ASAP7_75t_L g829 ( .A(n_774), .B(n_490), .Y(n_829) );
OAI21xp5_ASAP7_75t_L g830 ( .A1(n_679), .A2(n_511), .B(n_490), .Y(n_830) );
AOI21xp5_ASAP7_75t_L g831 ( .A1(n_763), .A2(n_530), .B(n_511), .Y(n_831) );
AND2x4_ASAP7_75t_L g832 ( .A(n_744), .B(n_17), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_708), .Y(n_833) );
OR2x2_ASAP7_75t_L g834 ( .A(n_676), .B(n_18), .Y(n_834) );
AOI21xp33_ASAP7_75t_L g835 ( .A1(n_687), .A2(n_511), .B(n_19), .Y(n_835) );
BUFx2_ASAP7_75t_L g836 ( .A(n_676), .Y(n_836) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_800), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_740), .Y(n_838) );
NAND3xp33_ASAP7_75t_L g839 ( .A(n_687), .B(n_511), .C(n_530), .Y(n_839) );
INVx3_ASAP7_75t_L g840 ( .A(n_684), .Y(n_840) );
OAI21x1_ASAP7_75t_L g841 ( .A1(n_756), .A2(n_511), .B(n_92), .Y(n_841) );
AND2x4_ASAP7_75t_L g842 ( .A(n_696), .B(n_19), .Y(n_842) );
AO31x2_ASAP7_75t_L g843 ( .A1(n_768), .A2(n_530), .A3(n_21), .B(n_22), .Y(n_843) );
O2A1O1Ixp33_ASAP7_75t_L g844 ( .A1(n_662), .A2(n_20), .B(n_23), .C(n_24), .Y(n_844) );
BUFx2_ASAP7_75t_L g845 ( .A(n_800), .Y(n_845) );
INVx3_ASAP7_75t_L g846 ( .A(n_725), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_714), .Y(n_847) );
OAI21x1_ASAP7_75t_SL g848 ( .A1(n_747), .A2(n_20), .B(n_23), .Y(n_848) );
A2O1A1Ixp33_ASAP7_75t_L g849 ( .A1(n_785), .A2(n_530), .B(n_27), .C(n_28), .Y(n_849) );
OA21x2_ASAP7_75t_L g850 ( .A1(n_746), .A2(n_530), .B(n_96), .Y(n_850) );
OR2x6_ASAP7_75t_L g851 ( .A(n_798), .B(n_25), .Y(n_851) );
AO31x2_ASAP7_75t_L g852 ( .A1(n_771), .A2(n_27), .A3(n_28), .B(n_30), .Y(n_852) );
INVxp67_ASAP7_75t_L g853 ( .A(n_683), .Y(n_853) );
OAI221xp5_ASAP7_75t_L g854 ( .A1(n_668), .A2(n_30), .B1(n_31), .B2(n_32), .C(n_33), .Y(n_854) );
OAI21x1_ASAP7_75t_L g855 ( .A1(n_702), .A2(n_99), .B(n_98), .Y(n_855) );
OA21x2_ASAP7_75t_L g856 ( .A1(n_790), .A2(n_103), .B(n_102), .Y(n_856) );
BUFx3_ASAP7_75t_L g857 ( .A(n_681), .Y(n_857) );
OAI21x1_ASAP7_75t_L g858 ( .A1(n_712), .A2(n_105), .B(n_104), .Y(n_858) );
OAI21x1_ASAP7_75t_L g859 ( .A1(n_712), .A2(n_115), .B(n_113), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_715), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_716), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_717), .Y(n_862) );
OAI21x1_ASAP7_75t_L g863 ( .A1(n_801), .A2(n_119), .B(n_117), .Y(n_863) );
NOR2x1_ASAP7_75t_SL g864 ( .A(n_700), .B(n_31), .Y(n_864) );
AO31x2_ASAP7_75t_L g865 ( .A1(n_771), .A2(n_32), .A3(n_33), .B(n_34), .Y(n_865) );
OAI21xp5_ASAP7_75t_L g866 ( .A1(n_679), .A2(n_34), .B(n_35), .Y(n_866) );
AOI21xp5_ASAP7_75t_L g867 ( .A1(n_742), .A2(n_132), .B(n_131), .Y(n_867) );
OAI21x1_ASAP7_75t_L g868 ( .A1(n_747), .A2(n_757), .B(n_729), .Y(n_868) );
INVx2_ASAP7_75t_L g869 ( .A(n_721), .Y(n_869) );
OAI21x1_ASAP7_75t_L g870 ( .A1(n_757), .A2(n_135), .B(n_134), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_723), .B(n_36), .Y(n_871) );
OAI21x1_ASAP7_75t_L g872 ( .A1(n_711), .A2(n_137), .B(n_136), .Y(n_872) );
OAI21x1_ASAP7_75t_L g873 ( .A1(n_711), .A2(n_142), .B(n_141), .Y(n_873) );
OR2x2_ASAP7_75t_L g874 ( .A(n_780), .B(n_37), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_769), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_750), .A2(n_37), .B1(n_38), .B2(n_39), .Y(n_876) );
INVx6_ASAP7_75t_L g877 ( .A(n_753), .Y(n_877) );
OA21x2_ASAP7_75t_L g878 ( .A1(n_751), .A2(n_145), .B(n_144), .Y(n_878) );
OAI222xp33_ASAP7_75t_L g879 ( .A1(n_709), .A2(n_38), .B1(n_41), .B2(n_42), .C1(n_43), .C2(n_44), .Y(n_879) );
AOI21xp5_ASAP7_75t_L g880 ( .A1(n_783), .A2(n_147), .B(n_146), .Y(n_880) );
OAI21x1_ASAP7_75t_L g881 ( .A1(n_729), .A2(n_151), .B(n_150), .Y(n_881) );
HB1xp67_ASAP7_75t_L g882 ( .A(n_766), .Y(n_882) );
BUFx6f_ASAP7_75t_L g883 ( .A(n_665), .Y(n_883) );
NOR2x1_ASAP7_75t_SL g884 ( .A(n_700), .B(n_41), .Y(n_884) );
AO21x2_ASAP7_75t_L g885 ( .A1(n_749), .A2(n_153), .B(n_152), .Y(n_885) );
INVx2_ASAP7_75t_L g886 ( .A(n_748), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_745), .Y(n_887) );
O2A1O1Ixp33_ASAP7_75t_SL g888 ( .A1(n_692), .A2(n_200), .B(n_311), .C(n_308), .Y(n_888) );
BUFx6f_ASAP7_75t_L g889 ( .A(n_665), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_672), .B(n_42), .Y(n_890) );
AND2x4_ASAP7_75t_L g891 ( .A(n_697), .B(n_46), .Y(n_891) );
INVx4_ASAP7_75t_SL g892 ( .A(n_665), .Y(n_892) );
AND2x4_ASAP7_75t_L g893 ( .A(n_698), .B(n_48), .Y(n_893) );
OR2x6_ASAP7_75t_SL g894 ( .A(n_720), .B(n_694), .Y(n_894) );
BUFx3_ASAP7_75t_L g895 ( .A(n_753), .Y(n_895) );
OAI21x1_ASAP7_75t_L g896 ( .A1(n_734), .A2(n_201), .B(n_307), .Y(n_896) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_760), .Y(n_897) );
OR2x6_ASAP7_75t_L g898 ( .A(n_700), .B(n_48), .Y(n_898) );
INVx2_ASAP7_75t_SL g899 ( .A(n_685), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_792), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_664), .B(n_49), .Y(n_901) );
CKINVDCx5p33_ASAP7_75t_R g902 ( .A(n_661), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_674), .Y(n_903) );
OAI21x1_ASAP7_75t_L g904 ( .A1(n_734), .A2(n_199), .B(n_302), .Y(n_904) );
AND2x4_ASAP7_75t_L g905 ( .A(n_695), .B(n_49), .Y(n_905) );
A2O1A1Ixp33_ASAP7_75t_L g906 ( .A1(n_779), .A2(n_50), .B(n_51), .C(n_52), .Y(n_906) );
AOI21xp5_ASAP7_75t_L g907 ( .A1(n_754), .A2(n_202), .B(n_301), .Y(n_907) );
OA21x2_ASAP7_75t_L g908 ( .A1(n_754), .A2(n_198), .B(n_300), .Y(n_908) );
OAI21xp5_ASAP7_75t_L g909 ( .A1(n_692), .A2(n_50), .B(n_51), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_722), .A2(n_52), .B1(n_53), .B2(n_54), .Y(n_910) );
NOR2xp33_ASAP7_75t_L g911 ( .A(n_739), .B(n_54), .Y(n_911) );
AND2x4_ASAP7_75t_L g912 ( .A(n_787), .B(n_55), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_791), .Y(n_913) );
NOR2xp33_ASAP7_75t_L g914 ( .A(n_736), .B(n_55), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_667), .A2(n_57), .B1(n_58), .B2(n_59), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_701), .Y(n_916) );
BUFx6f_ASAP7_75t_L g917 ( .A(n_804), .Y(n_917) );
BUFx2_ASAP7_75t_L g918 ( .A(n_784), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_701), .Y(n_919) );
INVx3_ASAP7_75t_L g920 ( .A(n_725), .Y(n_920) );
NOR2xp33_ASAP7_75t_L g921 ( .A(n_693), .B(n_59), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_730), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_713), .Y(n_923) );
OAI21x1_ASAP7_75t_L g924 ( .A1(n_724), .A2(n_211), .B(n_299), .Y(n_924) );
INVxp67_ASAP7_75t_L g925 ( .A(n_705), .Y(n_925) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_690), .B(n_61), .Y(n_926) );
OAI222xp33_ASAP7_75t_L g927 ( .A1(n_699), .A2(n_62), .B1(n_63), .B2(n_64), .C1(n_65), .C2(n_66), .Y(n_927) );
OAI21x1_ASAP7_75t_L g928 ( .A1(n_737), .A2(n_212), .B(n_298), .Y(n_928) );
OAI21x1_ASAP7_75t_SL g929 ( .A1(n_686), .A2(n_63), .B(n_64), .Y(n_929) );
OAI21x1_ASAP7_75t_L g930 ( .A1(n_762), .A2(n_214), .B(n_297), .Y(n_930) );
OA21x2_ASAP7_75t_L g931 ( .A1(n_793), .A2(n_209), .B(n_296), .Y(n_931) );
OAI21x1_ASAP7_75t_L g932 ( .A1(n_762), .A2(n_207), .B(n_295), .Y(n_932) );
OR2x6_ASAP7_75t_L g933 ( .A(n_804), .B(n_682), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_682), .B(n_65), .Y(n_934) );
AND2x4_ASAP7_75t_L g935 ( .A(n_728), .B(n_66), .Y(n_935) );
INVxp67_ASAP7_75t_SL g936 ( .A(n_705), .Y(n_936) );
OAI21x1_ASAP7_75t_L g937 ( .A1(n_772), .A2(n_205), .B(n_294), .Y(n_937) );
AO31x2_ASAP7_75t_L g938 ( .A1(n_699), .A2(n_67), .A3(n_68), .B(n_69), .Y(n_938) );
OAI21x1_ASAP7_75t_SL g939 ( .A1(n_686), .A2(n_67), .B(n_68), .Y(n_939) );
OR2x2_ASAP7_75t_L g940 ( .A(n_726), .B(n_69), .Y(n_940) );
OAI21x1_ASAP7_75t_SL g941 ( .A1(n_662), .A2(n_70), .B(n_71), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_730), .B(n_70), .Y(n_942) );
HB1xp67_ASAP7_75t_L g943 ( .A(n_784), .Y(n_943) );
A2O1A1Ixp33_ASAP7_75t_L g944 ( .A1(n_707), .A2(n_71), .B(n_72), .C(n_73), .Y(n_944) );
O2A1O1Ixp33_ASAP7_75t_L g945 ( .A1(n_707), .A2(n_72), .B(n_73), .C(n_74), .Y(n_945) );
BUFx3_ASAP7_75t_L g946 ( .A(n_776), .Y(n_946) );
INVx6_ASAP7_75t_L g947 ( .A(n_752), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_778), .Y(n_948) );
NAND2x1p5_ASAP7_75t_L g949 ( .A(n_804), .B(n_76), .Y(n_949) );
AOI21xp5_ASAP7_75t_L g950 ( .A1(n_703), .A2(n_219), .B(n_289), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_773), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_777), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_765), .B(n_76), .Y(n_953) );
NAND2x1p5_ASAP7_75t_L g954 ( .A(n_728), .B(n_77), .Y(n_954) );
NAND2x1p5_ASAP7_75t_L g955 ( .A(n_752), .B(n_77), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_732), .B(n_78), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_731), .Y(n_957) );
OAI21xp5_ASAP7_75t_L g958 ( .A1(n_732), .A2(n_79), .B(n_80), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_953), .A2(n_786), .B1(n_718), .B2(n_759), .Y(n_959) );
AOI21xp5_ASAP7_75t_L g960 ( .A1(n_830), .A2(n_758), .B(n_795), .Y(n_960) );
INVx2_ASAP7_75t_L g961 ( .A(n_833), .Y(n_961) );
OAI211xp5_ASAP7_75t_SL g962 ( .A1(n_853), .A2(n_765), .B(n_923), .C(n_913), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_898), .A2(n_718), .B1(n_767), .B2(n_789), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_812), .A2(n_703), .B1(n_690), .B2(n_764), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_916), .B(n_660), .Y(n_965) );
INVx1_ASAP7_75t_SL g966 ( .A(n_836), .Y(n_966) );
INVx2_ASAP7_75t_L g967 ( .A(n_860), .Y(n_967) );
NOR2xp33_ASAP7_75t_L g968 ( .A(n_853), .B(n_691), .Y(n_968) );
OAI22xp33_ASAP7_75t_L g969 ( .A1(n_812), .A2(n_761), .B1(n_677), .B2(n_795), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_898), .A2(n_733), .B1(n_761), .B2(n_671), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_898), .A2(n_761), .B1(n_663), .B2(n_666), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_914), .A2(n_794), .B1(n_673), .B2(n_678), .Y(n_972) );
AOI22xp33_ASAP7_75t_SL g973 ( .A1(n_823), .A2(n_710), .B1(n_755), .B2(n_775), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_936), .A2(n_775), .B1(n_743), .B2(n_741), .Y(n_974) );
INVx2_ASAP7_75t_L g975 ( .A(n_869), .Y(n_975) );
AO31x2_ASAP7_75t_L g976 ( .A1(n_818), .A2(n_704), .A3(n_710), .B(n_741), .Y(n_976) );
A2O1A1Ixp33_ASAP7_75t_L g977 ( .A1(n_926), .A2(n_921), .B(n_958), .C(n_866), .Y(n_977) );
HB1xp67_ASAP7_75t_L g978 ( .A(n_845), .Y(n_978) );
AOI21xp5_ASAP7_75t_L g979 ( .A1(n_830), .A2(n_794), .B(n_743), .Y(n_979) );
AOI21xp5_ASAP7_75t_L g980 ( .A1(n_831), .A2(n_741), .B(n_743), .Y(n_980) );
OR2x2_ASAP7_75t_L g981 ( .A(n_837), .B(n_897), .Y(n_981) );
CKINVDCx11_ASAP7_75t_R g982 ( .A(n_806), .Y(n_982) );
AOI22xp5_ASAP7_75t_SL g983 ( .A1(n_807), .A2(n_755), .B1(n_752), .B2(n_727), .Y(n_983) );
INVx2_ASAP7_75t_L g984 ( .A(n_813), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_819), .A2(n_775), .B1(n_710), .B2(n_688), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_936), .A2(n_710), .B1(n_81), .B2(n_83), .Y(n_986) );
NAND4xp25_ASAP7_75t_L g987 ( .A(n_844), .B(n_79), .C(n_81), .D(n_83), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_821), .A2(n_710), .B1(n_86), .B2(n_87), .Y(n_988) );
AOI22xp33_ASAP7_75t_SL g989 ( .A1(n_864), .A2(n_85), .B1(n_86), .B2(n_87), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_919), .B(n_85), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_837), .B(n_88), .Y(n_991) );
AOI22xp5_ASAP7_75t_L g992 ( .A1(n_912), .A2(n_88), .B1(n_89), .B2(n_90), .Y(n_992) );
AND2x4_ASAP7_75t_L g993 ( .A(n_811), .B(n_154), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_827), .Y(n_994) );
OR2x2_ASAP7_75t_L g995 ( .A(n_900), .B(n_155), .Y(n_995) );
AOI221xp5_ASAP7_75t_L g996 ( .A1(n_934), .A2(n_156), .B1(n_157), .B2(n_158), .C(n_163), .Y(n_996) );
INVx3_ASAP7_75t_L g997 ( .A(n_808), .Y(n_997) );
AOI222xp33_ASAP7_75t_L g998 ( .A1(n_876), .A2(n_165), .B1(n_166), .B2(n_167), .C1(n_169), .C2(n_174), .Y(n_998) );
AOI221xp5_ASAP7_75t_L g999 ( .A1(n_934), .A2(n_175), .B1(n_177), .B2(n_179), .C(n_180), .Y(n_999) );
OAI22xp33_ASAP7_75t_L g1000 ( .A1(n_825), .A2(n_186), .B1(n_187), .B2(n_189), .Y(n_1000) );
AOI322xp5_ASAP7_75t_L g1001 ( .A1(n_911), .A2(n_191), .A3(n_194), .B1(n_196), .B2(n_203), .C1(n_222), .C2(n_225), .Y(n_1001) );
NOR2xp33_ASAP7_75t_L g1002 ( .A(n_882), .B(n_227), .Y(n_1002) );
INVx2_ASAP7_75t_L g1003 ( .A(n_820), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_948), .B(n_229), .Y(n_1004) );
AOI22xp5_ASAP7_75t_L g1005 ( .A1(n_912), .A2(n_230), .B1(n_236), .B2(n_240), .Y(n_1005) );
BUFx6f_ASAP7_75t_L g1006 ( .A(n_808), .Y(n_1006) );
AOI22xp33_ASAP7_75t_SL g1007 ( .A1(n_884), .A2(n_241), .B1(n_247), .B2(n_248), .Y(n_1007) );
AOI21xp33_ASAP7_75t_L g1008 ( .A1(n_839), .A2(n_933), .B(n_940), .Y(n_1008) );
BUFx8_ASAP7_75t_SL g1009 ( .A(n_825), .Y(n_1009) );
AND2x4_ASAP7_75t_L g1010 ( .A(n_811), .B(n_249), .Y(n_1010) );
A2O1A1Ixp33_ASAP7_75t_L g1011 ( .A1(n_958), .A2(n_250), .B(n_252), .C(n_253), .Y(n_1011) );
OAI21xp5_ASAP7_75t_L g1012 ( .A1(n_868), .A2(n_839), .B(n_956), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_838), .Y(n_1013) );
OAI211xp5_ASAP7_75t_L g1014 ( .A1(n_844), .A2(n_257), .B(n_258), .C(n_259), .Y(n_1014) );
OR2x2_ASAP7_75t_L g1015 ( .A(n_874), .B(n_260), .Y(n_1015) );
A2O1A1Ixp33_ASAP7_75t_L g1016 ( .A1(n_866), .A2(n_267), .B(n_269), .C(n_271), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_821), .A2(n_272), .B1(n_273), .B2(n_274), .Y(n_1017) );
AOI22xp33_ASAP7_75t_SL g1018 ( .A1(n_851), .A2(n_276), .B1(n_277), .B2(n_278), .Y(n_1018) );
AOI21xp5_ASAP7_75t_L g1019 ( .A1(n_831), .A2(n_279), .B(n_280), .Y(n_1019) );
BUFx2_ASAP7_75t_L g1020 ( .A(n_828), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_832), .A2(n_281), .B1(n_312), .B2(n_933), .Y(n_1021) );
BUFx3_ASAP7_75t_L g1022 ( .A(n_808), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_832), .A2(n_933), .B1(n_851), .B2(n_942), .Y(n_1023) );
INVx2_ASAP7_75t_L g1024 ( .A(n_824), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_847), .B(n_861), .Y(n_1025) );
INVxp33_ASAP7_75t_L g1026 ( .A(n_815), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_862), .Y(n_1027) );
INVx3_ASAP7_75t_L g1028 ( .A(n_815), .Y(n_1028) );
OAI21x1_ASAP7_75t_L g1029 ( .A1(n_805), .A2(n_810), .B(n_826), .Y(n_1029) );
BUFx3_ASAP7_75t_L g1030 ( .A(n_815), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_822), .Y(n_1031) );
CKINVDCx14_ASAP7_75t_R g1032 ( .A(n_825), .Y(n_1032) );
AOI21xp33_ASAP7_75t_L g1033 ( .A1(n_945), .A2(n_835), .B(n_901), .Y(n_1033) );
HB1xp67_ASAP7_75t_L g1034 ( .A(n_851), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_822), .Y(n_1035) );
INVx2_ASAP7_75t_SL g1036 ( .A(n_877), .Y(n_1036) );
OA21x2_ASAP7_75t_L g1037 ( .A1(n_870), .A2(n_841), .B(n_924), .Y(n_1037) );
A2O1A1Ixp33_ASAP7_75t_L g1038 ( .A1(n_835), .A2(n_956), .B(n_945), .C(n_901), .Y(n_1038) );
OA21x2_ASAP7_75t_L g1039 ( .A1(n_928), .A2(n_950), .B(n_930), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_809), .B(n_816), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_942), .A2(n_891), .B1(n_893), .B2(n_842), .Y(n_1041) );
AND2x4_ASAP7_75t_L g1042 ( .A(n_892), .B(n_817), .Y(n_1042) );
INVx2_ASAP7_75t_L g1043 ( .A(n_951), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_809), .B(n_816), .Y(n_1044) );
CKINVDCx6p67_ASAP7_75t_R g1045 ( .A(n_895), .Y(n_1045) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_925), .A2(n_891), .B1(n_842), .B2(n_893), .Y(n_1046) );
HB1xp67_ASAP7_75t_L g1047 ( .A(n_857), .Y(n_1047) );
OR2x2_ASAP7_75t_L g1048 ( .A(n_834), .B(n_882), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_887), .B(n_952), .Y(n_1049) );
OAI22xp33_ASAP7_75t_L g1050 ( .A1(n_894), .A2(n_854), .B1(n_877), .B2(n_890), .Y(n_1050) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_925), .A2(n_905), .B1(n_954), .B2(n_955), .Y(n_1051) );
BUFx12f_ASAP7_75t_L g1052 ( .A(n_902), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1053 ( .A1(n_905), .A2(n_954), .B1(n_955), .B2(n_854), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_903), .B(n_871), .Y(n_1054) );
AOI221xp5_ASAP7_75t_L g1055 ( .A1(n_876), .A2(n_890), .B1(n_909), .B2(n_927), .C(n_941), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_918), .B(n_943), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_935), .A2(n_943), .B1(n_922), .B2(n_871), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_935), .A2(n_909), .B1(n_910), .B2(n_875), .Y(n_1058) );
AOI221xp5_ASAP7_75t_L g1059 ( .A1(n_927), .A2(n_879), .B1(n_939), .B2(n_929), .C(n_848), .Y(n_1059) );
CKINVDCx16_ASAP7_75t_R g1060 ( .A(n_946), .Y(n_1060) );
OAI22xp33_ASAP7_75t_L g1061 ( .A1(n_949), .A2(n_817), .B1(n_840), .B2(n_899), .Y(n_1061) );
OA21x2_ASAP7_75t_L g1062 ( .A1(n_950), .A2(n_932), .B(n_937), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_957), .Y(n_1063) );
AOI211xp5_ASAP7_75t_L g1064 ( .A1(n_879), .A2(n_906), .B(n_944), .C(n_849), .Y(n_1064) );
INVx2_ASAP7_75t_L g1065 ( .A(n_886), .Y(n_1065) );
O2A1O1Ixp33_ASAP7_75t_L g1066 ( .A1(n_814), .A2(n_888), .B(n_915), .C(n_818), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_840), .A2(n_920), .B1(n_846), .B2(n_814), .Y(n_1067) );
BUFx2_ASAP7_75t_L g1068 ( .A(n_947), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_938), .B(n_865), .Y(n_1069) );
A2O1A1Ixp33_ASAP7_75t_L g1070 ( .A1(n_867), .A2(n_907), .B(n_880), .C(n_920), .Y(n_1070) );
AOI22xp33_ASAP7_75t_SL g1071 ( .A1(n_949), .A2(n_846), .B1(n_878), .B2(n_829), .Y(n_1071) );
AOI21xp33_ASAP7_75t_L g1072 ( .A1(n_878), .A2(n_850), .B(n_885), .Y(n_1072) );
CKINVDCx11_ASAP7_75t_R g1073 ( .A(n_892), .Y(n_1073) );
AOI221xp5_ASAP7_75t_L g1074 ( .A1(n_867), .A2(n_907), .B1(n_880), .B2(n_917), .C(n_883), .Y(n_1074) );
OR2x2_ASAP7_75t_L g1075 ( .A(n_938), .B(n_852), .Y(n_1075) );
BUFx12f_ASAP7_75t_L g1076 ( .A(n_947), .Y(n_1076) );
OR2x2_ASAP7_75t_L g1077 ( .A(n_938), .B(n_852), .Y(n_1077) );
OR2x2_ASAP7_75t_L g1078 ( .A(n_852), .B(n_865), .Y(n_1078) );
A2O1A1Ixp33_ASAP7_75t_L g1079 ( .A1(n_872), .A2(n_881), .B(n_904), .C(n_896), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g1080 ( .A1(n_829), .A2(n_883), .B1(n_889), .B2(n_917), .Y(n_1080) );
INVx2_ASAP7_75t_SL g1081 ( .A(n_883), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_889), .A2(n_917), .B1(n_850), .B2(n_856), .Y(n_1082) );
AND2x4_ASAP7_75t_L g1083 ( .A(n_892), .B(n_889), .Y(n_1083) );
OAI221xp5_ASAP7_75t_L g1084 ( .A1(n_908), .A2(n_931), .B1(n_865), .B2(n_843), .C(n_885), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_843), .B(n_908), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_843), .B(n_873), .Y(n_1086) );
HB1xp67_ASAP7_75t_L g1087 ( .A(n_855), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1088 ( .A1(n_931), .A2(n_858), .B1(n_859), .B2(n_863), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_813), .Y(n_1089) );
AO31x2_ASAP7_75t_L g1090 ( .A1(n_818), .A2(n_781), .A3(n_768), .B(n_950), .Y(n_1090) );
AND2x4_ASAP7_75t_L g1091 ( .A(n_811), .B(n_670), .Y(n_1091) );
AOI22xp33_ASAP7_75t_SL g1092 ( .A1(n_823), .A2(n_709), .B1(n_720), .B2(n_812), .Y(n_1092) );
INVx11_ASAP7_75t_L g1093 ( .A(n_806), .Y(n_1093) );
AND2x4_ASAP7_75t_L g1094 ( .A(n_811), .B(n_670), .Y(n_1094) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_812), .A2(n_823), .B1(n_898), .B2(n_936), .Y(n_1095) );
INVx3_ASAP7_75t_L g1096 ( .A(n_808), .Y(n_1096) );
AND2x4_ASAP7_75t_L g1097 ( .A(n_811), .B(n_670), .Y(n_1097) );
OAI22xp33_ASAP7_75t_L g1098 ( .A1(n_812), .A2(n_595), .B1(n_661), .B2(n_709), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_961), .B(n_967), .Y(n_1099) );
INVx2_ASAP7_75t_L g1100 ( .A(n_1085), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_975), .B(n_1043), .Y(n_1101) );
OA21x2_ASAP7_75t_L g1102 ( .A1(n_1072), .A2(n_1012), .B(n_1084), .Y(n_1102) );
BUFx3_ASAP7_75t_L g1103 ( .A(n_1006), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1078), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1065), .B(n_1003), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1069), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1024), .B(n_1031), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1035), .B(n_984), .Y(n_1108) );
INVxp67_ASAP7_75t_L g1109 ( .A(n_1046), .Y(n_1109) );
BUFx2_ASAP7_75t_L g1110 ( .A(n_976), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_1050), .A2(n_1095), .B1(n_959), .B2(n_1092), .Y(n_1111) );
OR2x2_ASAP7_75t_L g1112 ( .A(n_1046), .B(n_981), .Y(n_1112) );
CKINVDCx5p33_ASAP7_75t_R g1113 ( .A(n_1009), .Y(n_1113) );
OR2x2_ASAP7_75t_L g1114 ( .A(n_966), .B(n_1095), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1040), .B(n_1044), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1075), .Y(n_1116) );
INVx3_ASAP7_75t_L g1117 ( .A(n_1006), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_994), .B(n_1013), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1027), .B(n_1089), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1063), .B(n_1025), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1025), .B(n_1041), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1077), .Y(n_1122) );
INVxp67_ASAP7_75t_SL g1123 ( .A(n_1051), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1049), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1049), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_977), .B(n_1038), .Y(n_1126) );
OR2x2_ASAP7_75t_L g1127 ( .A(n_966), .B(n_1048), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1054), .B(n_1055), .Y(n_1128) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1054), .Y(n_1129) );
BUFx3_ASAP7_75t_L g1130 ( .A(n_1006), .Y(n_1130) );
OAI21xp33_ASAP7_75t_L g1131 ( .A1(n_987), .A2(n_986), .B(n_1059), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1023), .B(n_1033), .Y(n_1132) );
INVxp67_ASAP7_75t_L g1133 ( .A(n_1034), .Y(n_1133) );
BUFx3_ASAP7_75t_L g1134 ( .A(n_1073), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_962), .A2(n_964), .B1(n_1032), .B2(n_987), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_1033), .B(n_964), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1056), .B(n_991), .Y(n_1137) );
AND2x4_ASAP7_75t_L g1138 ( .A(n_1083), .B(n_1081), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_965), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_965), .B(n_1091), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1091), .B(n_1094), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_986), .Y(n_1142) );
AND2x4_ASAP7_75t_L g1143 ( .A(n_1083), .B(n_1042), .Y(n_1143) );
INVx2_ASAP7_75t_L g1144 ( .A(n_1086), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1004), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1094), .B(n_1097), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1004), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1097), .B(n_990), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1051), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_990), .B(n_983), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1087), .Y(n_1151) );
INVx3_ASAP7_75t_L g1152 ( .A(n_1042), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1012), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_976), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_978), .B(n_997), .Y(n_1155) );
INVx2_ASAP7_75t_L g1156 ( .A(n_976), .Y(n_1156) );
INVx3_ASAP7_75t_L g1157 ( .A(n_1022), .Y(n_1157) );
INVx3_ASAP7_75t_L g1158 ( .A(n_1030), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_997), .B(n_1028), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1028), .B(n_1096), .Y(n_1160) );
INVx2_ASAP7_75t_L g1161 ( .A(n_1037), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1090), .Y(n_1162) );
AOI22xp5_ASAP7_75t_SL g1163 ( .A1(n_1053), .A2(n_1060), .B1(n_993), .B2(n_1010), .Y(n_1163) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1090), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1096), .B(n_1064), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1090), .Y(n_1166) );
BUFx3_ASAP7_75t_L g1167 ( .A(n_1076), .Y(n_1167) );
INVx3_ASAP7_75t_L g1168 ( .A(n_993), .Y(n_1168) );
AOI221xp5_ASAP7_75t_L g1169 ( .A1(n_1098), .A2(n_1053), .B1(n_963), .B2(n_968), .C(n_1057), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_974), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_974), .Y(n_1171) );
HB1xp67_ASAP7_75t_L g1172 ( .A(n_1020), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1084), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1026), .B(n_1058), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_998), .B(n_1010), .Y(n_1175) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_1008), .B(n_1070), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_998), .B(n_1015), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_992), .B(n_988), .Y(n_1178) );
HB1xp67_ASAP7_75t_L g1179 ( .A(n_1080), .Y(n_1179) );
OAI31xp33_ASAP7_75t_L g1180 ( .A1(n_1000), .A2(n_1014), .A3(n_1061), .B(n_1002), .Y(n_1180) );
INVx2_ASAP7_75t_L g1181 ( .A(n_1039), .Y(n_1181) );
NOR2xp33_ASAP7_75t_L g1182 ( .A(n_1047), .B(n_1036), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_995), .B(n_989), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1088), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g1185 ( .A(n_1008), .B(n_972), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_971), .B(n_970), .Y(n_1186) );
INVx2_ASAP7_75t_SL g1187 ( .A(n_1080), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1067), .B(n_973), .Y(n_1188) );
OR2x2_ASAP7_75t_L g1189 ( .A(n_1068), .B(n_960), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1088), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1001), .B(n_1018), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1062), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1062), .Y(n_1193) );
BUFx3_ASAP7_75t_L g1194 ( .A(n_1045), .Y(n_1194) );
BUFx2_ASAP7_75t_L g1195 ( .A(n_1074), .Y(n_1195) );
OR2x6_ASAP7_75t_L g1196 ( .A(n_979), .B(n_1066), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1021), .B(n_1005), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1016), .B(n_1011), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1071), .B(n_969), .Y(n_1199) );
INVx2_ASAP7_75t_L g1200 ( .A(n_1039), .Y(n_1200) );
HB1xp67_ASAP7_75t_L g1201 ( .A(n_980), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1007), .B(n_1017), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_996), .B(n_999), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1079), .Y(n_1204) );
NAND4xp25_ASAP7_75t_L g1205 ( .A(n_1135), .B(n_1082), .C(n_985), .D(n_1019), .Y(n_1205) );
AO31x2_ASAP7_75t_L g1206 ( .A1(n_1204), .A2(n_1029), .A3(n_1052), .B(n_1093), .Y(n_1206) );
HB1xp67_ASAP7_75t_L g1207 ( .A(n_1140), .Y(n_1207) );
BUFx2_ASAP7_75t_L g1208 ( .A(n_1141), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1106), .B(n_982), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1120), .B(n_1118), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1119), .Y(n_1211) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1161), .Y(n_1212) );
AND2x4_ASAP7_75t_L g1213 ( .A(n_1106), .B(n_1163), .Y(n_1213) );
OR2x2_ASAP7_75t_L g1214 ( .A(n_1127), .B(n_1137), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1100), .B(n_1144), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1100), .B(n_1144), .Y(n_1216) );
INVx2_ASAP7_75t_SL g1217 ( .A(n_1103), .Y(n_1217) );
AND2x4_ASAP7_75t_L g1218 ( .A(n_1163), .B(n_1100), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1119), .Y(n_1219) );
BUFx3_ASAP7_75t_L g1220 ( .A(n_1167), .Y(n_1220) );
AND2x4_ASAP7_75t_L g1221 ( .A(n_1144), .B(n_1104), .Y(n_1221) );
OAI221xp5_ASAP7_75t_L g1222 ( .A1(n_1111), .A2(n_1169), .B1(n_1131), .B2(n_1133), .C(n_1128), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1120), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1108), .Y(n_1224) );
NOR2xp33_ASAP7_75t_L g1225 ( .A(n_1128), .B(n_1121), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1108), .Y(n_1226) );
INVxp67_ASAP7_75t_SL g1227 ( .A(n_1168), .Y(n_1227) );
AOI22xp33_ASAP7_75t_L g1228 ( .A1(n_1175), .A2(n_1177), .B1(n_1191), .B2(n_1169), .Y(n_1228) );
BUFx3_ASAP7_75t_L g1229 ( .A(n_1167), .Y(n_1229) );
OAI221xp5_ASAP7_75t_L g1230 ( .A1(n_1131), .A2(n_1133), .B1(n_1180), .B2(n_1132), .C(n_1136), .Y(n_1230) );
INVxp67_ASAP7_75t_SL g1231 ( .A(n_1168), .Y(n_1231) );
BUFx3_ASAP7_75t_L g1232 ( .A(n_1141), .Y(n_1232) );
OAI221xp5_ASAP7_75t_L g1233 ( .A1(n_1180), .A2(n_1132), .B1(n_1136), .B2(n_1126), .C(n_1172), .Y(n_1233) );
AND2x4_ASAP7_75t_L g1234 ( .A(n_1104), .B(n_1116), .Y(n_1234) );
NOR2xp33_ASAP7_75t_L g1235 ( .A(n_1121), .B(n_1129), .Y(n_1235) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1124), .B(n_1125), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1116), .B(n_1122), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1122), .B(n_1140), .Y(n_1238) );
INVx1_ASAP7_75t_SL g1239 ( .A(n_1194), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1099), .Y(n_1240) );
INVx5_ASAP7_75t_SL g1241 ( .A(n_1143), .Y(n_1241) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1127), .B(n_1137), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1173), .B(n_1101), .Y(n_1243) );
OR2x2_ASAP7_75t_SL g1244 ( .A(n_1114), .B(n_1112), .Y(n_1244) );
OAI21xp5_ASAP7_75t_L g1245 ( .A1(n_1191), .A2(n_1203), .B(n_1175), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1124), .B(n_1125), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1115), .B(n_1146), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1129), .B(n_1107), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1173), .B(n_1149), .Y(n_1249) );
INVx3_ASAP7_75t_L g1250 ( .A(n_1168), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1107), .B(n_1139), .Y(n_1251) );
NAND2xp5_ASAP7_75t_SL g1252 ( .A(n_1168), .B(n_1150), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1149), .B(n_1105), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1105), .Y(n_1254) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1139), .Y(n_1255) );
AOI21xp33_ASAP7_75t_SL g1256 ( .A1(n_1113), .A2(n_1182), .B(n_1177), .Y(n_1256) );
NAND2xp5_ASAP7_75t_SL g1257 ( .A(n_1150), .B(n_1142), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1109), .B(n_1142), .Y(n_1258) );
INVx2_ASAP7_75t_L g1259 ( .A(n_1161), .Y(n_1259) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1155), .Y(n_1260) );
AOI22xp5_ASAP7_75t_L g1261 ( .A1(n_1183), .A2(n_1178), .B1(n_1148), .B2(n_1197), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1109), .B(n_1126), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1115), .Y(n_1263) );
AND2x4_ASAP7_75t_L g1264 ( .A(n_1123), .B(n_1165), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1162), .B(n_1164), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1162), .B(n_1164), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1165), .Y(n_1267) );
AND2x4_ASAP7_75t_L g1268 ( .A(n_1123), .B(n_1187), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1166), .B(n_1146), .Y(n_1269) );
NOR2xp33_ASAP7_75t_L g1270 ( .A(n_1183), .B(n_1148), .Y(n_1270) );
NAND2xp33_ASAP7_75t_SL g1271 ( .A(n_1114), .B(n_1112), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1166), .B(n_1153), .Y(n_1272) );
OAI321xp33_ASAP7_75t_L g1273 ( .A1(n_1176), .A2(n_1195), .A3(n_1185), .B1(n_1188), .B2(n_1199), .C(n_1202), .Y(n_1273) );
NAND3xp33_ASAP7_75t_L g1274 ( .A(n_1195), .B(n_1204), .C(n_1185), .Y(n_1274) );
AOI221xp5_ASAP7_75t_L g1275 ( .A1(n_1178), .A2(n_1176), .B1(n_1174), .B2(n_1153), .C(n_1184), .Y(n_1275) );
NOR2x1_ASAP7_75t_R g1276 ( .A(n_1194), .B(n_1134), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1184), .B(n_1190), .Y(n_1277) );
INVx3_ASAP7_75t_L g1278 ( .A(n_1103), .Y(n_1278) );
OAI31xp33_ASAP7_75t_SL g1279 ( .A1(n_1202), .A2(n_1188), .A3(n_1197), .B(n_1143), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1190), .B(n_1171), .Y(n_1280) );
INVx4_ASAP7_75t_L g1281 ( .A(n_1152), .Y(n_1281) );
AND2x4_ASAP7_75t_SL g1282 ( .A(n_1143), .B(n_1152), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1170), .B(n_1171), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1215), .B(n_1154), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1215), .B(n_1154), .Y(n_1285) );
BUFx2_ASAP7_75t_L g1286 ( .A(n_1220), .Y(n_1286) );
NAND2xp5_ASAP7_75t_L g1287 ( .A(n_1225), .B(n_1174), .Y(n_1287) );
OR2x2_ASAP7_75t_L g1288 ( .A(n_1214), .B(n_1242), .Y(n_1288) );
INVx2_ASAP7_75t_L g1289 ( .A(n_1212), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1225), .B(n_1145), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1211), .Y(n_1291) );
INVxp67_ASAP7_75t_L g1292 ( .A(n_1220), .Y(n_1292) );
AND2x4_ASAP7_75t_L g1293 ( .A(n_1221), .B(n_1187), .Y(n_1293) );
INVxp67_ASAP7_75t_L g1294 ( .A(n_1229), .Y(n_1294) );
NAND2x1_ASAP7_75t_L g1295 ( .A(n_1218), .B(n_1152), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1216), .B(n_1170), .Y(n_1296) );
AND2x4_ASAP7_75t_SL g1297 ( .A(n_1213), .B(n_1143), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_1223), .B(n_1145), .Y(n_1298) );
OR2x2_ASAP7_75t_L g1299 ( .A(n_1207), .B(n_1189), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1219), .Y(n_1300) );
CKINVDCx16_ASAP7_75t_R g1301 ( .A(n_1229), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1224), .B(n_1147), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1237), .Y(n_1303) );
NOR2xp67_ASAP7_75t_SL g1304 ( .A(n_1276), .B(n_1134), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1216), .B(n_1151), .Y(n_1305) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1237), .Y(n_1306) );
OR2x2_ASAP7_75t_L g1307 ( .A(n_1244), .B(n_1189), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1226), .B(n_1147), .Y(n_1308) );
AOI211x1_ASAP7_75t_SL g1309 ( .A1(n_1245), .A2(n_1199), .B(n_1156), .C(n_1200), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1269), .B(n_1151), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1269), .B(n_1156), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1258), .B(n_1156), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1258), .B(n_1110), .Y(n_1313) );
NAND4xp25_ASAP7_75t_L g1314 ( .A(n_1279), .B(n_1186), .C(n_1203), .D(n_1110), .Y(n_1314) );
AND2x4_ASAP7_75t_L g1315 ( .A(n_1221), .B(n_1187), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1234), .Y(n_1316) );
INVx2_ASAP7_75t_L g1317 ( .A(n_1212), .Y(n_1317) );
NOR2xp33_ASAP7_75t_L g1318 ( .A(n_1256), .B(n_1186), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1221), .B(n_1102), .Y(n_1319) );
NOR2xp33_ASAP7_75t_L g1320 ( .A(n_1222), .B(n_1152), .Y(n_1320) );
OR2x2_ASAP7_75t_L g1321 ( .A(n_1210), .B(n_1179), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1234), .Y(n_1322) );
OAI22xp5_ASAP7_75t_L g1323 ( .A1(n_1228), .A2(n_1158), .B1(n_1157), .B2(n_1179), .Y(n_1323) );
INVx2_ASAP7_75t_SL g1324 ( .A(n_1278), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1235), .B(n_1138), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1235), .B(n_1138), .Y(n_1326) );
INVxp67_ASAP7_75t_SL g1327 ( .A(n_1218), .Y(n_1327) );
INVx2_ASAP7_75t_L g1328 ( .A(n_1259), .Y(n_1328) );
OR2x2_ASAP7_75t_L g1329 ( .A(n_1267), .B(n_1193), .Y(n_1329) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1255), .Y(n_1330) );
NOR2xp33_ASAP7_75t_L g1331 ( .A(n_1261), .B(n_1158), .Y(n_1331) );
NAND3xp33_ASAP7_75t_L g1332 ( .A(n_1230), .B(n_1201), .C(n_1193), .Y(n_1332) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1238), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1249), .B(n_1102), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1238), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1336 ( .A(n_1249), .B(n_1102), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1253), .B(n_1102), .Y(n_1337) );
INVx2_ASAP7_75t_L g1338 ( .A(n_1259), .Y(n_1338) );
INVx1_ASAP7_75t_SL g1339 ( .A(n_1239), .Y(n_1339) );
AND4x1_ASAP7_75t_L g1340 ( .A(n_1209), .B(n_1198), .C(n_1159), .D(n_1160), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1253), .B(n_1192), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1240), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1283), .B(n_1192), .Y(n_1343) );
AOI31xp33_ASAP7_75t_L g1344 ( .A1(n_1213), .A2(n_1198), .A3(n_1159), .B(n_1160), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1283), .B(n_1181), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1287), .B(n_1262), .Y(n_1346) );
NAND2xp5_ASAP7_75t_SL g1347 ( .A(n_1301), .B(n_1213), .Y(n_1347) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1337), .B(n_1264), .Y(n_1348) );
AOI22xp5_ASAP7_75t_SL g1349 ( .A1(n_1318), .A2(n_1209), .B1(n_1218), .B2(n_1270), .Y(n_1349) );
BUFx2_ASAP7_75t_L g1350 ( .A(n_1286), .Y(n_1350) );
OR2x2_ASAP7_75t_L g1351 ( .A(n_1321), .B(n_1264), .Y(n_1351) );
INVx2_ASAP7_75t_L g1352 ( .A(n_1289), .Y(n_1352) );
NAND4xp25_ASAP7_75t_L g1353 ( .A(n_1318), .B(n_1233), .C(n_1275), .D(n_1270), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1333), .B(n_1262), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1330), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1335), .B(n_1243), .Y(n_1356) );
OR2x2_ASAP7_75t_L g1357 ( .A(n_1321), .B(n_1264), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1337), .B(n_1280), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1343), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1334), .B(n_1280), .Y(n_1360) );
OAI22xp5_ASAP7_75t_L g1361 ( .A1(n_1344), .A2(n_1257), .B1(n_1252), .B2(n_1232), .Y(n_1361) );
NAND2xp5_ASAP7_75t_L g1362 ( .A(n_1303), .B(n_1243), .Y(n_1362) );
INVx3_ASAP7_75t_SL g1363 ( .A(n_1339), .Y(n_1363) );
INVx2_ASAP7_75t_L g1364 ( .A(n_1289), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1343), .Y(n_1365) );
CKINVDCx16_ASAP7_75t_R g1366 ( .A(n_1288), .Y(n_1366) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1341), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1334), .B(n_1268), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1336), .B(n_1268), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1370 ( .A(n_1336), .B(n_1268), .Y(n_1370) );
OR2x2_ASAP7_75t_L g1371 ( .A(n_1299), .B(n_1277), .Y(n_1371) );
INVx2_ASAP7_75t_L g1372 ( .A(n_1317), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1319), .B(n_1277), .Y(n_1373) );
XNOR2x2_ASAP7_75t_L g1374 ( .A(n_1314), .B(n_1257), .Y(n_1374) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1306), .B(n_1254), .Y(n_1375) );
AOI21xp5_ASAP7_75t_L g1376 ( .A1(n_1332), .A2(n_1271), .B(n_1252), .Y(n_1376) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1341), .Y(n_1377) );
OR2x2_ASAP7_75t_L g1378 ( .A(n_1288), .B(n_1260), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1329), .Y(n_1379) );
INVxp67_ASAP7_75t_L g1380 ( .A(n_1304), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_1311), .B(n_1272), .Y(n_1381) );
NAND2xp5_ASAP7_75t_L g1382 ( .A(n_1290), .B(n_1263), .Y(n_1382) );
AND2x4_ASAP7_75t_L g1383 ( .A(n_1327), .B(n_1206), .Y(n_1383) );
OR2x2_ASAP7_75t_L g1384 ( .A(n_1307), .B(n_1271), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1311), .B(n_1266), .Y(n_1385) );
HB1xp67_ASAP7_75t_L g1386 ( .A(n_1292), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1284), .B(n_1266), .Y(n_1387) );
OR2x2_ASAP7_75t_L g1388 ( .A(n_1329), .B(n_1265), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1389 ( .A(n_1366), .B(n_1358), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1390 ( .A(n_1379), .B(n_1310), .Y(n_1390) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1355), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1392 ( .A(n_1379), .B(n_1296), .Y(n_1392) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1355), .Y(n_1393) );
INVx2_ASAP7_75t_L g1394 ( .A(n_1350), .Y(n_1394) );
OR2x2_ASAP7_75t_L g1395 ( .A(n_1388), .B(n_1310), .Y(n_1395) );
NAND2xp5_ASAP7_75t_L g1396 ( .A(n_1367), .B(n_1291), .Y(n_1396) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1367), .Y(n_1397) );
NAND2xp5_ASAP7_75t_L g1398 ( .A(n_1377), .B(n_1300), .Y(n_1398) );
NAND3xp33_ASAP7_75t_SL g1399 ( .A(n_1380), .B(n_1340), .C(n_1309), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1358), .B(n_1313), .Y(n_1400) );
AOI222xp33_ASAP7_75t_L g1401 ( .A1(n_1361), .A2(n_1273), .B1(n_1320), .B2(n_1331), .C1(n_1325), .C2(n_1326), .Y(n_1401) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1377), .Y(n_1402) );
AOI221xp5_ASAP7_75t_L g1403 ( .A1(n_1353), .A2(n_1320), .B1(n_1342), .B2(n_1331), .C(n_1323), .Y(n_1403) );
NOR2xp33_ASAP7_75t_L g1404 ( .A(n_1363), .B(n_1294), .Y(n_1404) );
AOI22xp5_ASAP7_75t_L g1405 ( .A1(n_1347), .A2(n_1297), .B1(n_1316), .B2(n_1322), .Y(n_1405) );
AOI32xp33_ASAP7_75t_L g1406 ( .A1(n_1350), .A2(n_1297), .A3(n_1208), .B1(n_1247), .B2(n_1232), .Y(n_1406) );
NAND2xp5_ASAP7_75t_L g1407 ( .A(n_1359), .B(n_1305), .Y(n_1407) );
OAI21xp5_ASAP7_75t_L g1408 ( .A1(n_1376), .A2(n_1274), .B(n_1295), .Y(n_1408) );
AOI32xp33_ASAP7_75t_L g1409 ( .A1(n_1374), .A2(n_1282), .A3(n_1293), .B1(n_1315), .B2(n_1305), .Y(n_1409) );
OR2x2_ASAP7_75t_L g1410 ( .A(n_1388), .B(n_1285), .Y(n_1410) );
BUFx2_ASAP7_75t_L g1411 ( .A(n_1386), .Y(n_1411) );
OAI22xp5_ASAP7_75t_L g1412 ( .A1(n_1349), .A2(n_1251), .B1(n_1248), .B2(n_1241), .Y(n_1412) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1359), .Y(n_1413) );
OAI22xp5_ASAP7_75t_L g1414 ( .A1(n_1384), .A2(n_1351), .B1(n_1357), .B2(n_1378), .Y(n_1414) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1365), .Y(n_1415) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1391), .Y(n_1416) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1393), .Y(n_1417) );
A2O1A1Ixp33_ASAP7_75t_L g1418 ( .A1(n_1409), .A2(n_1378), .B(n_1383), .C(n_1387), .Y(n_1418) );
HB1xp67_ASAP7_75t_L g1419 ( .A(n_1411), .Y(n_1419) );
AOI22xp5_ASAP7_75t_L g1420 ( .A1(n_1401), .A2(n_1346), .B1(n_1348), .B2(n_1365), .Y(n_1420) );
OR2x2_ASAP7_75t_L g1421 ( .A(n_1410), .B(n_1371), .Y(n_1421) );
INVx1_ASAP7_75t_SL g1422 ( .A(n_1389), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1423 ( .A(n_1400), .B(n_1360), .Y(n_1423) );
INVx2_ASAP7_75t_L g1424 ( .A(n_1397), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1402), .Y(n_1425) );
NOR2xp33_ASAP7_75t_L g1426 ( .A(n_1404), .B(n_1382), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_1394), .B(n_1360), .Y(n_1427) );
NAND2xp5_ASAP7_75t_L g1428 ( .A(n_1403), .B(n_1373), .Y(n_1428) );
OAI21xp5_ASAP7_75t_L g1429 ( .A1(n_1408), .A2(n_1324), .B(n_1387), .Y(n_1429) );
NAND3xp33_ASAP7_75t_L g1430 ( .A(n_1408), .B(n_1324), .C(n_1357), .Y(n_1430) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1413), .Y(n_1431) );
AOI21xp33_ASAP7_75t_L g1432 ( .A1(n_1412), .A2(n_1308), .B(n_1302), .Y(n_1432) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1415), .B(n_1373), .Y(n_1433) );
OAI211xp5_ASAP7_75t_L g1434 ( .A1(n_1420), .A2(n_1406), .B(n_1399), .C(n_1405), .Y(n_1434) );
OAI21xp5_ASAP7_75t_L g1435 ( .A1(n_1430), .A2(n_1414), .B(n_1395), .Y(n_1435) );
OAI21xp33_ASAP7_75t_L g1436 ( .A1(n_1418), .A2(n_1392), .B(n_1390), .Y(n_1436) );
OAI21xp5_ASAP7_75t_L g1437 ( .A1(n_1429), .A2(n_1398), .B(n_1396), .Y(n_1437) );
AOI221xp5_ASAP7_75t_L g1438 ( .A1(n_1428), .A2(n_1392), .B1(n_1407), .B2(n_1354), .C(n_1348), .Y(n_1438) );
OAI221xp5_ASAP7_75t_SL g1439 ( .A1(n_1422), .A2(n_1371), .B1(n_1362), .B2(n_1356), .C(n_1368), .Y(n_1439) );
NAND3xp33_ASAP7_75t_L g1440 ( .A(n_1419), .B(n_1205), .C(n_1375), .Y(n_1440) );
O2A1O1Ixp5_ASAP7_75t_L g1441 ( .A1(n_1432), .A2(n_1298), .B(n_1281), .C(n_1236), .Y(n_1441) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1425), .Y(n_1442) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1425), .Y(n_1443) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1431), .Y(n_1444) );
AOI22xp33_ASAP7_75t_L g1445 ( .A1(n_1426), .A2(n_1369), .B1(n_1368), .B2(n_1370), .Y(n_1445) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1442), .Y(n_1446) );
NAND3xp33_ASAP7_75t_L g1447 ( .A(n_1434), .B(n_1417), .C(n_1416), .Y(n_1447) );
AOI221xp5_ASAP7_75t_L g1448 ( .A1(n_1436), .A2(n_1433), .B1(n_1424), .B2(n_1427), .C(n_1423), .Y(n_1448) );
AOI211xp5_ASAP7_75t_L g1449 ( .A1(n_1435), .A2(n_1421), .B(n_1423), .C(n_1427), .Y(n_1449) );
OAI21xp33_ASAP7_75t_SL g1450 ( .A1(n_1445), .A2(n_1385), .B(n_1381), .Y(n_1450) );
OAI21xp33_ASAP7_75t_L g1451 ( .A1(n_1439), .A2(n_1424), .B(n_1369), .Y(n_1451) );
O2A1O1Ixp33_ASAP7_75t_L g1452 ( .A1(n_1441), .A2(n_1246), .B(n_1217), .C(n_1231), .Y(n_1452) );
INVx2_ASAP7_75t_SL g1453 ( .A(n_1443), .Y(n_1453) );
NOR3xp33_ASAP7_75t_SL g1454 ( .A(n_1447), .B(n_1440), .C(n_1438), .Y(n_1454) );
OAI22x1_ASAP7_75t_L g1455 ( .A1(n_1453), .A2(n_1444), .B1(n_1441), .B2(n_1281), .Y(n_1455) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1446), .Y(n_1456) );
AND2x4_ASAP7_75t_L g1457 ( .A(n_1450), .B(n_1437), .Y(n_1457) );
NOR2xp33_ASAP7_75t_R g1458 ( .A(n_1452), .B(n_1157), .Y(n_1458) );
NAND5xp2_ASAP7_75t_L g1459 ( .A(n_1454), .B(n_1449), .C(n_1448), .D(n_1451), .E(n_1227), .Y(n_1459) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1456), .Y(n_1460) );
NAND3xp33_ASAP7_75t_SL g1461 ( .A(n_1458), .B(n_1372), .C(n_1364), .Y(n_1461) );
AOI22x1_ASAP7_75t_L g1462 ( .A1(n_1460), .A2(n_1455), .B1(n_1457), .B2(n_1158), .Y(n_1462) );
INVx2_ASAP7_75t_L g1463 ( .A(n_1459), .Y(n_1463) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1461), .Y(n_1464) );
NAND3xp33_ASAP7_75t_L g1465 ( .A(n_1463), .B(n_1130), .C(n_1117), .Y(n_1465) );
OR3x1_ASAP7_75t_L g1466 ( .A(n_1465), .B(n_1464), .C(n_1462), .Y(n_1466) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1466), .Y(n_1467) );
AOI322xp5_ASAP7_75t_L g1468 ( .A1(n_1467), .A2(n_1250), .A3(n_1312), .B1(n_1284), .B2(n_1345), .C1(n_1352), .C2(n_1372), .Y(n_1468) );
OAI22xp33_ASAP7_75t_L g1469 ( .A1(n_1468), .A2(n_1196), .B1(n_1338), .B2(n_1328), .Y(n_1469) );
endmodule