module real_aes_5430_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_974, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_975, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_974;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_975;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_919;
wire n_857;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_931;
wire n_904;
wire n_780;
wire n_570;
wire n_675;
wire n_840;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_281;
wire n_496;
wire n_962;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_310;
wire n_960;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_947;
wire n_561;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_713;
wire n_288;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_354;
wire n_265;
wire n_972;
wire n_968;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_266;
wire n_312;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_949;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_259;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_0), .A2(n_25), .B1(n_452), .B2(n_453), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_1), .A2(n_52), .B1(n_727), .B2(n_730), .Y(n_764) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_2), .Y(n_260) );
AND2x4_ASAP7_75t_L g696 ( .A(n_2), .B(n_242), .Y(n_696) );
AND2x4_ASAP7_75t_L g701 ( .A(n_2), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g447 ( .A(n_3), .Y(n_447) );
INVx1_ASAP7_75t_SL g511 ( .A(n_4), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_5), .A2(n_84), .B1(n_584), .B2(n_585), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_6), .A2(n_86), .B1(n_660), .B2(n_662), .Y(n_659) );
AOI221x1_ASAP7_75t_L g916 ( .A1(n_7), .A2(n_8), .B1(n_917), .B2(n_918), .C(n_919), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_9), .A2(n_114), .B1(n_354), .B2(n_355), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_10), .A2(n_62), .B1(n_347), .B2(n_373), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g963 ( .A1(n_11), .A2(n_159), .B1(n_303), .B2(n_428), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_12), .A2(n_101), .B1(n_405), .B2(n_501), .Y(n_500) );
AOI21xp33_ASAP7_75t_SL g454 ( .A1(n_13), .A2(n_455), .B(n_456), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_14), .A2(n_232), .B1(n_343), .B2(n_344), .Y(n_957) );
INVx1_ASAP7_75t_L g528 ( .A(n_15), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_16), .A2(n_35), .B1(n_382), .B2(n_385), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g931 ( .A(n_17), .Y(n_931) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_18), .A2(n_92), .B1(n_705), .B2(n_720), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_19), .A2(n_218), .B1(n_334), .B2(n_335), .Y(n_956) );
INVx1_ASAP7_75t_L g417 ( .A(n_20), .Y(n_417) );
AO22x1_ASAP7_75t_L g966 ( .A1(n_21), .A2(n_145), .B1(n_432), .B2(n_433), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_22), .A2(n_139), .B1(n_388), .B2(n_392), .Y(n_387) );
INVx1_ASAP7_75t_L g753 ( .A(n_23), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_24), .A2(n_98), .B1(n_355), .B2(n_435), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_26), .A2(n_57), .B1(n_452), .B2(n_464), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_27), .A2(n_153), .B1(n_402), .B2(n_612), .Y(n_611) );
CKINVDCx5p33_ASAP7_75t_R g933 ( .A(n_28), .Y(n_933) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_29), .A2(n_179), .B1(n_488), .B2(n_554), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_30), .A2(n_200), .B1(n_378), .B2(n_492), .Y(n_559) );
INVx1_ASAP7_75t_L g408 ( .A(n_31), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_32), .A2(n_87), .B1(n_693), .B2(n_697), .Y(n_692) );
AOI22xp33_ASAP7_75t_SL g923 ( .A1(n_33), .A2(n_69), .B1(n_364), .B2(n_367), .Y(n_923) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_34), .A2(n_71), .B1(n_335), .B2(n_343), .Y(n_425) );
INVx1_ASAP7_75t_SL g803 ( .A(n_36), .Y(n_803) );
INVx1_ASAP7_75t_L g644 ( .A(n_37), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_38), .A2(n_156), .B1(n_492), .B2(n_632), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g958 ( .A1(n_39), .A2(n_321), .B(n_959), .Y(n_958) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_40), .B(n_194), .Y(n_258) );
INVx1_ASAP7_75t_L g295 ( .A(n_40), .Y(n_295) );
INVxp67_ASAP7_75t_L g341 ( .A(n_40), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_41), .A2(n_102), .B1(n_700), .B2(n_715), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g319 ( .A1(n_42), .A2(n_78), .B1(n_320), .B2(n_321), .C(n_323), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_43), .B(n_459), .Y(n_458) );
AO22x1_ASAP7_75t_L g964 ( .A1(n_44), .A2(n_138), .B1(n_354), .B2(n_355), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_45), .B(n_616), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_46), .A2(n_120), .B1(n_303), .B2(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_47), .B(n_280), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_48), .A2(n_238), .B1(n_546), .B2(n_547), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_49), .A2(n_241), .B1(n_554), .B2(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_50), .A2(n_226), .B1(n_376), .B2(n_378), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_51), .A2(n_127), .B1(n_590), .B2(n_591), .Y(n_589) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_52), .A2(n_270), .B(n_356), .Y(n_269) );
NAND4xp25_ASAP7_75t_L g356 ( .A(n_52), .B(n_271), .C(n_318), .D(n_345), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_53), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_54), .A2(n_248), .B1(n_712), .B2(n_713), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g539 ( .A1(n_55), .A2(n_81), .B1(n_540), .B2(n_541), .C(n_543), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_56), .A2(n_175), .B1(n_273), .B2(n_298), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_58), .A2(n_222), .B1(n_549), .B2(n_550), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_59), .A2(n_171), .B1(n_298), .B2(n_364), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_60), .A2(n_192), .B1(n_463), .B2(n_464), .Y(n_462) );
NAND2xp33_ASAP7_75t_L g420 ( .A(n_61), .B(n_421), .Y(n_420) );
OAI22x1_ASAP7_75t_L g653 ( .A1(n_63), .A2(n_654), .B1(n_679), .B2(n_680), .Y(n_653) );
INVx1_ASAP7_75t_L g680 ( .A(n_63), .Y(n_680) );
INVxp67_ASAP7_75t_R g755 ( .A(n_64), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_65), .A2(n_231), .B1(n_577), .B2(n_658), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_66), .A2(n_149), .B1(n_582), .B2(n_585), .Y(n_678) );
INVx2_ASAP7_75t_L g255 ( .A(n_67), .Y(n_255) );
INVx1_ASAP7_75t_L g642 ( .A(n_68), .Y(n_642) );
AOI21xp33_ASAP7_75t_L g617 ( .A1(n_70), .A2(n_618), .B(n_619), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_72), .A2(n_214), .B1(n_370), .B2(n_371), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_73), .A2(n_167), .B1(n_469), .B2(n_471), .Y(n_468) );
INVx1_ASAP7_75t_L g695 ( .A(n_74), .Y(n_695) );
AND2x4_ASAP7_75t_L g698 ( .A(n_74), .B(n_255), .Y(n_698) );
INVx1_ASAP7_75t_SL g721 ( .A(n_74), .Y(n_721) );
INVx1_ASAP7_75t_L g532 ( .A(n_75), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_76), .B(n_320), .Y(n_955) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_77), .A2(n_79), .B1(n_475), .B2(n_490), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_80), .B(n_569), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_82), .A2(n_186), .B1(n_705), .B2(n_720), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_83), .A2(n_151), .B1(n_347), .B2(n_351), .Y(n_346) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_85), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_88), .A2(n_176), .B1(n_343), .B2(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g439 ( .A(n_89), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_90), .A2(n_184), .B1(n_334), .B2(n_423), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_91), .A2(n_103), .B1(n_672), .B2(n_673), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_93), .A2(n_169), .B1(n_334), .B2(n_335), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_94), .A2(n_100), .B1(n_396), .B2(n_399), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_95), .A2(n_235), .B1(n_303), .B2(n_308), .Y(n_302) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_96), .A2(n_188), .B1(n_402), .B2(n_404), .C(n_407), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_97), .A2(n_210), .B1(n_351), .B2(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_99), .B(n_335), .Y(n_534) );
INVx1_ASAP7_75t_SL g915 ( .A(n_102), .Y(n_915) );
NOR3xp33_ASAP7_75t_L g940 ( .A(n_102), .B(n_941), .C(n_942), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g948 ( .A1(n_102), .A2(n_949), .B1(n_967), .B2(n_969), .Y(n_948) );
CKINVDCx16_ASAP7_75t_R g751 ( .A(n_104), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_105), .A2(n_157), .B1(n_700), .B2(n_703), .Y(n_699) );
AO22x1_ASAP7_75t_L g570 ( .A1(n_106), .A2(n_185), .B1(n_571), .B2(n_572), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_107), .A2(n_206), .B1(n_351), .B2(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g281 ( .A(n_108), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_108), .B(n_193), .Y(n_338) );
INVx1_ASAP7_75t_L g324 ( .A(n_109), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_110), .A2(n_211), .B1(n_385), .B2(n_557), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_111), .A2(n_950), .B1(n_951), .B2(n_952), .Y(n_949) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_111), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_112), .A2(n_219), .B1(n_574), .B2(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g620 ( .A(n_113), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_115), .A2(n_152), .B1(n_347), .B2(n_473), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g934 ( .A(n_116), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_117), .A2(n_233), .B1(n_371), .B2(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g722 ( .A(n_118), .Y(n_722) );
INVx1_ASAP7_75t_L g960 ( .A(n_119), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_121), .A2(n_158), .B1(n_693), .B2(n_713), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_122), .B(n_495), .Y(n_649) );
XOR2x2_ASAP7_75t_L g563 ( .A(n_123), .B(n_564), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_124), .A2(n_174), .B1(n_435), .B2(n_436), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_125), .A2(n_170), .B1(n_475), .B2(n_490), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_126), .A2(n_133), .B1(n_428), .B2(n_436), .Y(n_924) );
INVx1_ASAP7_75t_L g457 ( .A(n_128), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_129), .A2(n_201), .B1(n_464), .B2(n_614), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_130), .A2(n_172), .B1(n_298), .B2(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_131), .A2(n_164), .B1(n_697), .B2(n_712), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_132), .A2(n_220), .B1(n_363), .B2(n_365), .Y(n_362) );
AO22x1_ASAP7_75t_L g965 ( .A1(n_134), .A2(n_239), .B1(n_435), .B2(n_436), .Y(n_965) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_135), .A2(n_191), .B1(n_354), .B2(n_355), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_136), .A2(n_215), .B1(n_557), .B2(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g530 ( .A(n_137), .Y(n_530) );
INVx1_ASAP7_75t_L g503 ( .A(n_140), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_141), .A2(n_567), .B(n_570), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_142), .A2(n_162), .B1(n_475), .B2(n_587), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_143), .A2(n_205), .B1(n_354), .B2(n_355), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_144), .A2(n_154), .B1(n_467), .B2(n_471), .Y(n_486) );
AOI22x1_ASAP7_75t_L g358 ( .A1(n_146), .A2(n_359), .B1(n_360), .B2(n_409), .Y(n_358) );
INVx1_ASAP7_75t_L g409 ( .A(n_146), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_147), .A2(n_160), .B1(n_303), .B2(n_428), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_148), .A2(n_223), .B1(n_727), .B2(n_730), .Y(n_739) );
INVx1_ASAP7_75t_L g724 ( .A(n_150), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_155), .A2(n_163), .B1(n_490), .B2(n_630), .Y(n_629) );
AOI22xp33_ASAP7_75t_SL g576 ( .A1(n_161), .A2(n_183), .B1(n_577), .B2(n_578), .Y(n_576) );
INVx1_ASAP7_75t_L g526 ( .A(n_165), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_166), .A2(n_228), .B1(n_354), .B2(n_355), .Y(n_519) );
OA22x2_ASAP7_75t_L g286 ( .A1(n_168), .A2(n_194), .B1(n_280), .B2(n_284), .Y(n_286) );
INVx1_ASAP7_75t_L g315 ( .A(n_168), .Y(n_315) );
AOI21xp5_ASAP7_75t_SL g524 ( .A1(n_173), .A2(n_321), .B(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_177), .A2(n_195), .B1(n_463), .B2(n_495), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_178), .A2(n_196), .B1(n_432), .B2(n_433), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_180), .A2(n_234), .B1(n_469), .B2(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_181), .A2(n_221), .B1(n_581), .B2(n_582), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g929 ( .A(n_182), .Y(n_929) );
AND2x2_ASAP7_75t_L g919 ( .A(n_187), .B(n_920), .Y(n_919) );
CKINVDCx6p67_ASAP7_75t_R g750 ( .A(n_189), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_190), .A2(n_208), .B1(n_432), .B2(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g297 ( .A(n_193), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_193), .B(n_313), .Y(n_331) );
OAI21xp33_ASAP7_75t_L g316 ( .A1(n_194), .A2(n_212), .B(n_317), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_197), .A2(n_227), .B1(n_303), .B2(n_428), .Y(n_516) );
INVx1_ASAP7_75t_L g522 ( .A(n_198), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_199), .Y(n_536) );
INVx1_ASAP7_75t_L g647 ( .A(n_202), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_203), .A2(n_247), .B1(n_700), .B2(n_715), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_204), .A2(n_224), .B1(n_354), .B2(n_557), .Y(n_914) );
INVx1_ASAP7_75t_L g638 ( .A(n_207), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_209), .A2(n_245), .B1(n_435), .B2(n_436), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_212), .B(n_236), .Y(n_259) );
INVx1_ASAP7_75t_L g283 ( .A(n_212), .Y(n_283) );
INVx1_ASAP7_75t_SL g650 ( .A(n_213), .Y(n_650) );
INVx1_ASAP7_75t_L g804 ( .A(n_216), .Y(n_804) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_217), .A2(n_243), .B1(n_392), .B2(n_664), .C(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g602 ( .A(n_223), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_225), .A2(n_237), .B1(n_378), .B2(n_492), .Y(n_491) );
AOI21xp33_ASAP7_75t_SL g437 ( .A1(n_229), .A2(n_321), .B(n_438), .Y(n_437) );
AOI21xp33_ASAP7_75t_L g636 ( .A1(n_230), .A2(n_540), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_236), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_240), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g702 ( .A(n_242), .Y(n_702) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_242), .Y(n_971) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_244), .Y(n_544) );
INVx1_ASAP7_75t_L g666 ( .A(n_246), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_261), .B(n_683), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
BUFx4_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
NAND3xp33_ASAP7_75t_L g252 ( .A(n_253), .B(n_256), .C(n_260), .Y(n_252) );
AND2x2_ASAP7_75t_L g945 ( .A(n_253), .B(n_946), .Y(n_945) );
AND2x2_ASAP7_75t_L g968 ( .A(n_253), .B(n_947), .Y(n_968) );
AOI21xp5_ASAP7_75t_L g972 ( .A1(n_253), .A2(n_260), .B(n_721), .Y(n_972) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AO21x1_ASAP7_75t_L g970 ( .A1(n_254), .A2(n_971), .B(n_972), .Y(n_970) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g694 ( .A(n_255), .B(n_695), .Y(n_694) );
AND3x4_ASAP7_75t_L g720 ( .A(n_255), .B(n_701), .C(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g946 ( .A(n_256), .B(n_947), .Y(n_946) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AO21x2_ASAP7_75t_L g327 ( .A1(n_257), .A2(n_328), .B(n_330), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g947 ( .A(n_260), .Y(n_947) );
XNOR2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_505), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_264), .B1(n_442), .B2(n_504), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
XOR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_414), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_357), .B1(n_410), .B2(n_412), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g413 ( .A(n_267), .Y(n_413) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND3x1_ASAP7_75t_L g270 ( .A(n_271), .B(n_318), .C(n_345), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_302), .Y(n_271) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g364 ( .A(n_274), .Y(n_364) );
INVx1_ASAP7_75t_L g672 ( .A(n_274), .Y(n_672) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
BUFx12f_ASAP7_75t_L g475 ( .A(n_275), .Y(n_475) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_275), .Y(n_630) );
AND2x4_ASAP7_75t_L g275 ( .A(n_276), .B(n_287), .Y(n_275) );
AND2x2_ASAP7_75t_L g299 ( .A(n_276), .B(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g348 ( .A(n_276), .B(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g352 ( .A(n_276), .B(n_305), .Y(n_352) );
AND2x4_ASAP7_75t_L g432 ( .A(n_276), .B(n_287), .Y(n_432) );
AND2x4_ASAP7_75t_L g433 ( .A(n_276), .B(n_300), .Y(n_433) );
AND2x4_ASAP7_75t_L g435 ( .A(n_276), .B(n_349), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_276), .B(n_384), .Y(n_436) );
AND2x4_ASAP7_75t_L g276 ( .A(n_277), .B(n_285), .Y(n_276) );
AND2x2_ASAP7_75t_L g322 ( .A(n_277), .B(n_286), .Y(n_322) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g304 ( .A(n_278), .B(n_286), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_282), .Y(n_278) );
NAND2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx2_ASAP7_75t_L g284 ( .A(n_280), .Y(n_284) );
INVx3_ASAP7_75t_L g290 ( .A(n_280), .Y(n_290) );
NAND2xp33_ASAP7_75t_L g296 ( .A(n_280), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g317 ( .A(n_280), .Y(n_317) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_280), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_281), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
OAI21xp5_ASAP7_75t_L g340 ( .A1(n_283), .A2(n_317), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g339 ( .A(n_286), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g334 ( .A(n_287), .B(n_304), .Y(n_334) );
AND2x4_ASAP7_75t_L g343 ( .A(n_287), .B(n_322), .Y(n_343) );
AND2x2_ASAP7_75t_L g391 ( .A(n_287), .B(n_304), .Y(n_391) );
AND2x4_ASAP7_75t_L g403 ( .A(n_287), .B(n_322), .Y(n_403) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_292), .Y(n_287) );
INVx2_ASAP7_75t_L g301 ( .A(n_288), .Y(n_301) );
OR2x2_ASAP7_75t_L g306 ( .A(n_288), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g336 ( .A(n_288), .B(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_L g349 ( .A(n_288), .B(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_290), .B(n_295), .Y(n_294) );
INVxp67_ASAP7_75t_L g313 ( .A(n_290), .Y(n_313) );
NAND3xp33_ASAP7_75t_L g330 ( .A(n_291), .B(n_312), .C(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g300 ( .A(n_292), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g307 ( .A(n_293), .Y(n_307) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
BUFx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g368 ( .A(n_299), .Y(n_368) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_299), .Y(n_490) );
BUFx5_ASAP7_75t_L g588 ( .A(n_299), .Y(n_588) );
AND2x2_ASAP7_75t_L g320 ( .A(n_300), .B(n_304), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_300), .B(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g344 ( .A(n_300), .B(n_311), .Y(n_344) );
AND2x4_ASAP7_75t_L g398 ( .A(n_300), .B(n_322), .Y(n_398) );
AND2x4_ASAP7_75t_L g400 ( .A(n_300), .B(n_311), .Y(n_400) );
AND2x2_ASAP7_75t_L g406 ( .A(n_300), .B(n_304), .Y(n_406) );
AND2x4_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
AND2x4_ASAP7_75t_L g354 ( .A(n_304), .B(n_349), .Y(n_354) );
AND2x2_ASAP7_75t_L g377 ( .A(n_304), .B(n_349), .Y(n_377) );
AND2x4_ASAP7_75t_L g383 ( .A(n_304), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g470 ( .A(n_304), .B(n_349), .Y(n_470) );
AND2x4_ASAP7_75t_L g310 ( .A(n_305), .B(n_311), .Y(n_310) );
AND2x4_ASAP7_75t_L g428 ( .A(n_305), .B(n_311), .Y(n_428) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g384 ( .A(n_306), .Y(n_384) );
INVx1_ASAP7_75t_L g350 ( .A(n_307), .Y(n_350) );
INVx3_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx5_ASAP7_75t_L g467 ( .A(n_309), .Y(n_467) );
INVx2_ASAP7_75t_L g558 ( .A(n_309), .Y(n_558) );
INVx2_ASAP7_75t_L g606 ( .A(n_309), .Y(n_606) );
INVx6_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx12f_ASAP7_75t_L g385 ( .A(n_310), .Y(n_385) );
AND2x4_ASAP7_75t_L g355 ( .A(n_311), .B(n_349), .Y(n_355) );
AND2x4_ASAP7_75t_L g380 ( .A(n_311), .B(n_349), .Y(n_380) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_316), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_332), .Y(n_318) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_320), .Y(n_421) );
INVx2_ASAP7_75t_L g523 ( .A(n_320), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_325), .B(n_408), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_325), .B(n_620), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_325), .B(n_666), .Y(n_665) );
INVx4_ASAP7_75t_L g920 ( .A(n_325), .Y(n_920) );
INVx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx4_ASAP7_75t_L g502 ( .A(n_326), .Y(n_502) );
INVx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_327), .Y(n_441) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_329), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_342), .Y(n_332) );
INVx1_ASAP7_75t_L g533 ( .A(n_334), .Y(n_533) );
INVx2_ASAP7_75t_L g935 ( .A(n_334), .Y(n_935) );
INVx4_ASAP7_75t_L g930 ( .A(n_335), .Y(n_930) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_339), .Y(n_335) );
AND2x4_ASAP7_75t_L g394 ( .A(n_336), .B(n_339), .Y(n_394) );
INVx2_ASAP7_75t_L g529 ( .A(n_343), .Y(n_529) );
INVx2_ASAP7_75t_L g424 ( .A(n_344), .Y(n_424) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_353), .Y(n_345) );
BUFx12f_ASAP7_75t_L g370 ( .A(n_347), .Y(n_370) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_347), .Y(n_670) );
BUFx12f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_348), .Y(n_488) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_348), .Y(n_628) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_352), .Y(n_373) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_352), .Y(n_554) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g411 ( .A(n_358), .Y(n_411) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND4xp75_ASAP7_75t_L g360 ( .A(n_361), .B(n_374), .C(n_386), .D(n_401), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_369), .Y(n_361) );
BUFx4f_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_381), .Y(n_374) );
BUFx8_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_377), .Y(n_492) );
INVx4_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g473 ( .A(n_379), .Y(n_473) );
INVx2_ASAP7_75t_L g592 ( .A(n_379), .Y(n_592) );
INVx4_ASAP7_75t_L g632 ( .A(n_379), .Y(n_632) );
INVx1_ASAP7_75t_L g677 ( .A(n_379), .Y(n_677) );
INVx8_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx3_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx12f_ASAP7_75t_L g471 ( .A(n_383), .Y(n_471) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_383), .Y(n_557) );
BUFx3_ASAP7_75t_L g582 ( .A(n_385), .Y(n_582) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_395), .Y(n_386) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g614 ( .A(n_390), .Y(n_614) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_391), .Y(n_463) );
BUFx3_ASAP7_75t_L g546 ( .A(n_391), .Y(n_546) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx4_ASAP7_75t_L g495 ( .A(n_393), .Y(n_495) );
INVx2_ASAP7_75t_L g547 ( .A(n_393), .Y(n_547) );
INVx2_ASAP7_75t_L g571 ( .A(n_393), .Y(n_571) );
INVx5_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx2_ASAP7_75t_L g453 ( .A(n_394), .Y(n_453) );
BUFx4f_ASAP7_75t_L g612 ( .A(n_394), .Y(n_612) );
INVx2_ASAP7_75t_L g643 ( .A(n_396), .Y(n_643) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_398), .Y(n_455) );
INVx2_ASAP7_75t_L g499 ( .A(n_398), .Y(n_499) );
BUFx3_ASAP7_75t_L g549 ( .A(n_398), .Y(n_549) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_398), .Y(n_618) );
BUFx8_ASAP7_75t_SL g917 ( .A(n_398), .Y(n_917) );
BUFx3_ASAP7_75t_L g575 ( .A(n_399), .Y(n_575) );
INVx4_ASAP7_75t_L g645 ( .A(n_399), .Y(n_645) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_400), .Y(n_464) );
INVx3_ASAP7_75t_L g551 ( .A(n_400), .Y(n_551) );
BUFx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx3_ASAP7_75t_L g452 ( .A(n_403), .Y(n_452) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_403), .Y(n_540) );
BUFx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g461 ( .A(n_406), .Y(n_461) );
INVx3_ASAP7_75t_L g542 ( .A(n_406), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_409), .A2(n_726), .B1(n_728), .B2(n_729), .Y(n_725) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVx3_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
XNOR2x1_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
NOR2x1_ASAP7_75t_L g418 ( .A(n_419), .B(n_426), .Y(n_418) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .C(n_425), .Y(n_419) );
INVxp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI22xp33_ASAP7_75t_L g527 ( .A1(n_424), .A2(n_528), .B1(n_529), .B2(n_530), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_424), .A2(n_929), .B1(n_930), .B2(n_931), .Y(n_928) );
NAND4xp25_ASAP7_75t_SL g426 ( .A(n_427), .B(n_429), .C(n_430), .D(n_437), .Y(n_426) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_434), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_440), .B(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_440), .B(n_544), .Y(n_543) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_441), .B(n_526), .Y(n_525) );
INVx2_ASAP7_75t_SL g572 ( .A(n_441), .Y(n_572) );
INVx1_ASAP7_75t_L g640 ( .A(n_441), .Y(n_640) );
INVx1_ASAP7_75t_L g504 ( .A(n_442), .Y(n_504) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
XNOR2x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_482), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI21x1_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_448), .B(n_476), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_446), .B(n_462), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_447), .Y(n_446) );
NOR2xp67_ASAP7_75t_L g448 ( .A(n_449), .B(n_465), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_458), .C(n_462), .Y(n_449) );
INVx1_ASAP7_75t_L g480 ( .A(n_450), .Y(n_480) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .Y(n_450) );
BUFx2_ASAP7_75t_L g577 ( .A(n_452), .Y(n_577) );
BUFx3_ASAP7_75t_L g574 ( .A(n_455), .Y(n_574) );
INVxp67_ASAP7_75t_L g478 ( .A(n_458), .Y(n_478) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_459), .Y(n_664) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g569 ( .A(n_460), .Y(n_569) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx3_ASAP7_75t_L g648 ( .A(n_463), .Y(n_648) );
BUFx3_ASAP7_75t_L g658 ( .A(n_463), .Y(n_658) );
INVx1_ASAP7_75t_L g481 ( .A(n_465), .Y(n_481) );
NAND4xp25_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .C(n_472), .D(n_474), .Y(n_465) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx3_ASAP7_75t_L g585 ( .A(n_471), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_481), .Y(n_476) );
NOR3xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .C(n_480), .Y(n_477) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
XOR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_503), .Y(n_483) );
NOR2x1_ASAP7_75t_L g484 ( .A(n_485), .B(n_493), .Y(n_484) );
NAND4xp25_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .C(n_489), .D(n_491), .Y(n_485) );
BUFx2_ASAP7_75t_SL g590 ( .A(n_488), .Y(n_590) );
BUFx2_ASAP7_75t_SL g673 ( .A(n_490), .Y(n_673) );
BUFx3_ASAP7_75t_L g584 ( .A(n_492), .Y(n_584) );
NAND4xp25_ASAP7_75t_L g493 ( .A(n_494), .B(n_496), .C(n_497), .D(n_500), .Y(n_493) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx4_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g959 ( .A(n_502), .B(n_960), .Y(n_959) );
XNOR2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_595), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_562), .B1(n_593), .B2(n_594), .Y(n_506) );
INVx1_ASAP7_75t_L g593 ( .A(n_507), .Y(n_593) );
BUFx2_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
OA22x2_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_535), .B1(n_560), .B2(n_561), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
XNOR2x1_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
XNOR2xp5_ASAP7_75t_L g561 ( .A(n_511), .B(n_512), .Y(n_561) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_520), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_517), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
NOR3xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_527), .C(n_531), .Y(n_520) );
OAI21xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_524), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_529), .A2(n_933), .B1(n_934), .B2(n_935), .Y(n_932) );
OAI21xp5_ASAP7_75t_SL g531 ( .A1(n_532), .A2(n_533), .B(n_534), .Y(n_531) );
INVxp67_ASAP7_75t_SL g560 ( .A(n_535), .Y(n_560) );
XNOR2x1_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_552), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_545), .C(n_548), .Y(n_538) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g616 ( .A(n_542), .Y(n_616) );
INVx2_ASAP7_75t_L g918 ( .A(n_542), .Y(n_918) );
BUFx2_ASAP7_75t_L g578 ( .A(n_546), .Y(n_578) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g662 ( .A(n_551), .Y(n_662) );
NAND4xp25_ASAP7_75t_SL g552 ( .A(n_553), .B(n_555), .C(n_556), .D(n_559), .Y(n_552) );
BUFx3_ASAP7_75t_L g581 ( .A(n_554), .Y(n_581) );
BUFx2_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g594 ( .A(n_563), .Y(n_594) );
NOR2x1_ASAP7_75t_L g564 ( .A(n_565), .B(n_579), .Y(n_564) );
NAND3xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_573), .C(n_576), .Y(n_565) );
INVx2_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND4xp25_ASAP7_75t_SL g579 ( .A(n_580), .B(n_583), .C(n_586), .D(n_589), .Y(n_579) );
BUFx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
BUFx2_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_652), .B1(n_681), .B2(n_682), .Y(n_595) );
INVx1_ASAP7_75t_L g681 ( .A(n_596), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B1(n_621), .B2(n_651), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVxp67_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
XNOR2x1_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
NOR2x1_ASAP7_75t_L g603 ( .A(n_604), .B(n_610), .Y(n_603) );
NAND4xp25_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .C(n_608), .D(n_609), .Y(n_604) );
NAND4xp25_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .C(n_615), .D(n_617), .Y(n_610) );
INVx2_ASAP7_75t_L g661 ( .A(n_618), .Y(n_661) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g651 ( .A(n_623), .Y(n_651) );
XOR2x1_ASAP7_75t_L g623 ( .A(n_624), .B(n_650), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_633), .Y(n_624) );
AND4x1_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .C(n_629), .D(n_631), .Y(n_625) );
NOR3xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_641), .C(n_646), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_635), .B(n_636), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B1(n_644), .B2(n_645), .Y(n_641) );
OAI21xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B(n_649), .Y(n_646) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
BUFx3_ASAP7_75t_L g682 ( .A(n_653), .Y(n_682) );
OR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_667), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_655), .B(n_667), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_663), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2x1p5_ASAP7_75t_L g667 ( .A(n_668), .B(n_674), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_678), .Y(n_674) );
BUFx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_901), .B1(n_904), .B2(n_943), .C(n_948), .Y(n_683) );
NOR3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_806), .C(n_866), .Y(n_684) );
AOI31xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_774), .A3(n_792), .B(n_800), .Y(n_685) );
AOI211xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_706), .B(n_757), .C(n_765), .Y(n_686) );
INVx3_ASAP7_75t_L g881 ( .A(n_687), .Y(n_881) );
INVx3_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_688), .B(n_818), .Y(n_817) );
AOI221xp5_ASAP7_75t_L g826 ( .A1(n_688), .A2(n_827), .B1(n_830), .B2(n_832), .C(n_834), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_688), .B(n_759), .Y(n_843) );
INVx3_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_689), .B(n_746), .Y(n_812) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NOR3xp33_ASAP7_75t_L g813 ( .A(n_690), .B(n_737), .C(n_814), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_690), .B(n_709), .Y(n_847) );
INVx3_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_691), .B(n_709), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_691), .B(n_784), .Y(n_831) );
OR2x2_ASAP7_75t_L g864 ( .A(n_691), .B(n_709), .Y(n_864) );
AND2x2_ASAP7_75t_L g868 ( .A(n_691), .B(n_828), .Y(n_868) );
AND2x2_ASAP7_75t_L g874 ( .A(n_691), .B(n_710), .Y(n_874) );
INVx1_ASAP7_75t_L g886 ( .A(n_691), .Y(n_886) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_691), .B(n_836), .Y(n_900) );
AND2x4_ASAP7_75t_L g691 ( .A(n_692), .B(n_699), .Y(n_691) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
AND2x4_ASAP7_75t_L g700 ( .A(n_694), .B(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g712 ( .A(n_694), .B(n_696), .Y(n_712) );
AND2x2_ASAP7_75t_L g730 ( .A(n_694), .B(n_696), .Y(n_730) );
AND2x4_ASAP7_75t_L g697 ( .A(n_696), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g713 ( .A(n_696), .B(n_698), .Y(n_713) );
AND2x2_ASAP7_75t_L g727 ( .A(n_696), .B(n_698), .Y(n_727) );
INVx2_ASAP7_75t_L g756 ( .A(n_697), .Y(n_756) );
AND2x4_ASAP7_75t_L g705 ( .A(n_698), .B(n_701), .Y(n_705) );
AND2x4_ASAP7_75t_L g715 ( .A(n_698), .B(n_701), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_698), .B(n_701), .Y(n_723) );
INVx3_ASAP7_75t_L g749 ( .A(n_700), .Y(n_749) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
OAI22xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_731), .B1(n_742), .B2(n_744), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_716), .Y(n_707) );
OAI211xp5_ASAP7_75t_SL g834 ( .A1(n_708), .A2(n_835), .B(n_839), .C(n_852), .Y(n_834) );
INVx3_ASAP7_75t_L g850 ( .A(n_708), .Y(n_850) );
INVx3_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g818 ( .A(n_709), .B(n_747), .Y(n_818) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g745 ( .A(n_710), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g784 ( .A(n_710), .B(n_747), .Y(n_784) );
OR2x2_ASAP7_75t_L g791 ( .A(n_710), .B(n_747), .Y(n_791) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_714), .Y(n_710) );
INVx3_ASAP7_75t_L g754 ( .A(n_712), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_716), .B(n_745), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_716), .B(n_746), .Y(n_759) );
AND2x2_ASAP7_75t_L g781 ( .A(n_716), .B(n_782), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_716), .B(n_791), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_716), .B(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_716), .B(n_784), .Y(n_814) );
AND2x2_ASAP7_75t_L g823 ( .A(n_716), .B(n_773), .Y(n_823) );
A2O1A1Ixp33_ASAP7_75t_L g852 ( .A1(n_716), .A2(n_736), .B(n_828), .C(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g860 ( .A(n_716), .Y(n_860) );
CKINVDCx6p67_ASAP7_75t_R g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_717), .B(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g810 ( .A(n_717), .B(n_770), .Y(n_810) );
INVx1_ASAP7_75t_L g837 ( .A(n_717), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_717), .B(n_841), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_717), .B(n_746), .Y(n_849) );
AND2x2_ASAP7_75t_L g857 ( .A(n_717), .B(n_780), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_717), .A2(n_760), .B1(n_859), .B2(n_861), .Y(n_858) );
OR2x6_ASAP7_75t_SL g717 ( .A(n_718), .B(n_725), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_723), .A2(n_749), .B1(n_750), .B2(n_751), .Y(n_748) );
OAI221xp5_ASAP7_75t_L g802 ( .A1(n_723), .A2(n_749), .B1(n_803), .B2(n_804), .C(n_805), .Y(n_802) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_740), .Y(n_731) );
AND2x2_ASAP7_75t_L g761 ( .A(n_732), .B(n_762), .Y(n_761) );
AND2x2_ASAP7_75t_L g822 ( .A(n_732), .B(n_823), .Y(n_822) );
AND2x2_ASAP7_75t_SL g853 ( .A(n_732), .B(n_773), .Y(n_853) );
AND2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_736), .Y(n_732) );
INVx1_ASAP7_75t_L g741 ( .A(n_733), .Y(n_741) );
AND2x2_ASAP7_75t_L g770 ( .A(n_733), .B(n_737), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
AND2x2_ASAP7_75t_L g780 ( .A(n_736), .B(n_741), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_736), .B(n_782), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_736), .B(n_781), .Y(n_829) );
CKINVDCx5p33_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g740 ( .A(n_737), .B(n_741), .Y(n_740) );
OR2x2_ASAP7_75t_L g833 ( .A(n_737), .B(n_762), .Y(n_833) );
AND2x4_ASAP7_75t_SL g737 ( .A(n_738), .B(n_739), .Y(n_737) );
AND2x2_ASAP7_75t_L g787 ( .A(n_740), .B(n_773), .Y(n_787) );
INVx1_ASAP7_75t_L g841 ( .A(n_740), .Y(n_841) );
AND2x2_ASAP7_75t_L g862 ( .A(n_740), .B(n_762), .Y(n_862) );
INVx1_ASAP7_75t_L g743 ( .A(n_741), .Y(n_743) );
AND2x2_ASAP7_75t_L g838 ( .A(n_741), .B(n_782), .Y(n_838) );
AND2x2_ASAP7_75t_L g844 ( .A(n_741), .B(n_773), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_741), .B(n_782), .Y(n_898) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OAI211xp5_ASAP7_75t_L g884 ( .A1(n_745), .A2(n_865), .B(n_885), .C(n_887), .Y(n_884) );
INVx3_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g768 ( .A(n_747), .Y(n_768) );
OR2x2_ASAP7_75t_L g747 ( .A(n_748), .B(n_752), .Y(n_747) );
INVx1_ASAP7_75t_L g903 ( .A(n_749), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B1(n_755), .B2(n_756), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_760), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_761), .A2(n_793), .B1(n_795), .B2(n_799), .Y(n_792) );
CKINVDCx6p67_ASAP7_75t_R g773 ( .A(n_762), .Y(n_773) );
INVx1_ASAP7_75t_L g783 ( .A(n_762), .Y(n_783) );
AND2x2_ASAP7_75t_L g871 ( .A(n_762), .B(n_810), .Y(n_871) );
AND2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVxp67_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_769), .Y(n_766) );
AND2x2_ASAP7_75t_L g799 ( .A(n_767), .B(n_793), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_767), .A2(n_786), .B1(n_828), .B2(n_829), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_767), .B(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
BUFx2_ASAP7_75t_L g821 ( .A(n_768), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g885 ( .A(n_768), .B(n_886), .Y(n_885) );
O2A1O1Ixp33_ASAP7_75t_L g891 ( .A1(n_769), .A2(n_784), .B(n_878), .C(n_892), .Y(n_891) );
AND2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
INVx1_ASAP7_75t_L g778 ( .A(n_770), .Y(n_778) );
NAND3xp33_ASAP7_75t_L g848 ( .A(n_770), .B(n_849), .C(n_850), .Y(n_848) );
AND2x2_ASAP7_75t_L g878 ( .A(n_770), .B(n_781), .Y(n_878) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_773), .B(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_773), .B(n_780), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_773), .B(n_857), .Y(n_856) );
AOI21xp33_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_784), .B(n_785), .Y(n_774) );
INVxp67_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_777), .B(n_779), .Y(n_776) );
INVx1_ASAP7_75t_L g788 ( .A(n_777), .Y(n_788) );
AOI21xp33_ASAP7_75t_SL g896 ( .A1(n_778), .A2(n_897), .B(n_899), .Y(n_896) );
AND2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_780), .B(n_823), .Y(n_825) );
AOI211xp5_ASAP7_75t_L g815 ( .A1(n_782), .A2(n_816), .B(n_819), .C(n_824), .Y(n_815) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AOI221xp5_ASAP7_75t_L g839 ( .A1(n_784), .A2(n_840), .B1(n_842), .B2(n_844), .C(n_845), .Y(n_839) );
AOI21xp33_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_788), .B(n_789), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_786), .B(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g828 ( .A(n_791), .Y(n_828) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
A2O1A1Ixp33_ASAP7_75t_L g882 ( .A1(n_796), .A2(n_861), .B(n_883), .C(n_884), .Y(n_882) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
BUFx3_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g851 ( .A(n_802), .Y(n_851) );
AOI32xp33_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_815), .A3(n_826), .B1(n_854), .B2(n_865), .Y(n_806) );
O2A1O1Ixp33_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_810), .B(n_811), .C(n_813), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_809), .B(n_831), .Y(n_892) );
OAI21xp5_ASAP7_75t_L g889 ( .A1(n_810), .A2(n_868), .B(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
AOI221xp5_ASAP7_75t_SL g893 ( .A1(n_816), .A2(n_838), .B1(n_894), .B2(n_895), .C(n_896), .Y(n_893) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g883 ( .A(n_818), .Y(n_883) );
AND2x2_ASAP7_75t_L g819 ( .A(n_820), .B(n_822), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_820), .B(n_825), .Y(n_824) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
A2O1A1Ixp33_ASAP7_75t_SL g854 ( .A1(n_821), .A2(n_855), .B(n_858), .C(n_863), .Y(n_854) );
INVx1_ASAP7_75t_L g879 ( .A(n_825), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_828), .B(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
AOI31xp33_ASAP7_75t_L g869 ( .A1(n_833), .A2(n_870), .A3(n_872), .B(n_873), .Y(n_869) );
AOI21xp5_ASAP7_75t_L g890 ( .A1(n_833), .A2(n_870), .B(n_873), .Y(n_890) );
INVx1_ASAP7_75t_L g894 ( .A(n_835), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_838), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_836), .B(n_862), .Y(n_888) );
INVx3_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g846 ( .A(n_838), .Y(n_846) );
INVxp67_ASAP7_75t_SL g842 ( .A(n_843), .Y(n_842) );
A2O1A1Ixp33_ASAP7_75t_L g867 ( .A1(n_844), .A2(n_859), .B(n_868), .C(n_869), .Y(n_867) );
OAI211xp5_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_847), .B(n_848), .C(n_851), .Y(n_845) );
INVx1_ASAP7_75t_L g895 ( .A(n_847), .Y(n_895) );
CKINVDCx16_ASAP7_75t_R g865 ( .A(n_851), .Y(n_865) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
CKINVDCx14_ASAP7_75t_R g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
NAND5xp2_ASAP7_75t_L g866 ( .A(n_867), .B(n_875), .C(n_889), .D(n_891), .E(n_893), .Y(n_866) );
INVx1_ASAP7_75t_L g872 ( .A(n_868), .Y(n_872) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
O2A1O1Ixp33_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_879), .B(n_880), .C(n_882), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
CKINVDCx5p33_ASAP7_75t_R g901 ( .A(n_902), .Y(n_901) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVxp67_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx2_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
BUFx3_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
NAND2x1_ASAP7_75t_L g911 ( .A(n_912), .B(n_936), .Y(n_911) );
NOR3xp33_ASAP7_75t_L g912 ( .A(n_913), .B(n_921), .C(n_925), .Y(n_912) );
OAI22xp33_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_915), .B1(n_916), .B2(n_974), .Y(n_913) );
INVx1_ASAP7_75t_L g941 ( .A(n_914), .Y(n_941) );
NOR2xp67_ASAP7_75t_L g921 ( .A(n_915), .B(n_922), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_915), .A2(n_926), .B1(n_927), .B2(n_975), .Y(n_925) );
INVx1_ASAP7_75t_L g938 ( .A(n_916), .Y(n_938) );
NAND3xp33_ASAP7_75t_L g936 ( .A(n_922), .B(n_937), .C(n_940), .Y(n_936) );
AND2x2_ASAP7_75t_L g922 ( .A(n_923), .B(n_924), .Y(n_922) );
INVx1_ASAP7_75t_L g942 ( .A(n_926), .Y(n_942) );
INVx1_ASAP7_75t_L g939 ( .A(n_927), .Y(n_939) );
NOR2x1_ASAP7_75t_L g927 ( .A(n_928), .B(n_932), .Y(n_927) );
NOR2xp33_ASAP7_75t_L g937 ( .A(n_938), .B(n_939), .Y(n_937) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
HB1xp67_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
INVxp33_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_954), .B(n_961), .Y(n_953) );
AND4x1_ASAP7_75t_L g954 ( .A(n_955), .B(n_956), .C(n_957), .D(n_958), .Y(n_954) );
NOR4xp25_ASAP7_75t_L g961 ( .A(n_962), .B(n_964), .C(n_965), .D(n_966), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
HB1xp67_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
endmodule