module fake_jpeg_15633_n_270 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.C(n_1),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_43),
.Y(n_65)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_42),
.Y(n_54)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_1),
.C(n_2),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_49),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_30),
.B1(n_31),
.B2(n_19),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_57),
.B1(n_16),
.B2(n_36),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_43),
.B1(n_38),
.B2(n_36),
.Y(n_68)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_43),
.B1(n_30),
.B2(n_40),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_61),
.B1(n_62),
.B2(n_43),
.Y(n_67)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_66),
.Y(n_84)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_41),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_18),
.B1(n_23),
.B2(n_21),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_33),
.B(n_17),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_19),
.B1(n_16),
.B2(n_21),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_19),
.B1(n_16),
.B2(n_25),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_38),
.B1(n_36),
.B2(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_32),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_68),
.B1(n_38),
.B2(n_39),
.Y(n_95)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_76),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_35),
.B(n_34),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_78),
.B(n_81),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_35),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_50),
.C(n_35),
.Y(n_94)
);

INVx2_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_58),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_38),
.B1(n_23),
.B2(n_18),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_35),
.B(n_43),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_85),
.B(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_25),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_62),
.Y(n_108)
);

AOI32xp33_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_38),
.A3(n_41),
.B1(n_22),
.B2(n_26),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_24),
.Y(n_87)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_88),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_91),
.B(n_92),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_88),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_75),
.C(n_77),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_101),
.B1(n_48),
.B2(n_63),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_70),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_97),
.Y(n_123)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_103),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_45),
.B1(n_52),
.B2(n_49),
.Y(n_100)
);

AO21x1_ASAP7_75t_L g137 ( 
.A1(n_100),
.A2(n_105),
.B(n_39),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_45),
.B1(n_39),
.B2(n_60),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_70),
.Y(n_103)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_80),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_83),
.B1(n_82),
.B2(n_84),
.Y(n_118)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_50),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_73),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_98),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_114),
.A2(n_121),
.B(n_130),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_85),
.Y(n_116)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_116),
.A2(n_132),
.B(n_137),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_118),
.A2(n_122),
.B1(n_124),
.B2(n_101),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_111),
.B1(n_102),
.B2(n_99),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_127),
.C(n_94),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_90),
.B(n_93),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_82),
.B1(n_77),
.B2(n_89),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_77),
.B1(n_48),
.B2(n_63),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_102),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_125),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_87),
.C(n_73),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_98),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_44),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_136),
.Y(n_145)
);

INVxp67_ASAP7_75t_SL g138 ( 
.A(n_104),
.Y(n_138)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_136),
.B(n_107),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_147),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_90),
.B(n_93),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_158),
.B(n_22),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_160),
.C(n_162),
.Y(n_169)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_113),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_149),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_103),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_59),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_72),
.B1(n_74),
.B2(n_64),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_107),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_17),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_105),
.B(n_95),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_159),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_106),
.C(n_91),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_119),
.A2(n_106),
.B1(n_99),
.B2(n_97),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_161),
.A2(n_123),
.B1(n_128),
.B2(n_97),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_92),
.C(n_58),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_137),
.B1(n_124),
.B2(n_132),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_166),
.A2(n_167),
.B1(n_154),
.B2(n_157),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_137),
.B1(n_130),
.B2(n_114),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_134),
.B(n_126),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_170),
.A2(n_171),
.B(n_174),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_158),
.A2(n_134),
.B(n_125),
.Y(n_171)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_115),
.B(n_74),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_177),
.A2(n_80),
.B(n_28),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_58),
.C(n_48),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_185),
.C(n_151),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_140),
.B1(n_150),
.B2(n_153),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_44),
.Y(n_181)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_187),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_26),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_41),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_72),
.Y(n_186)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_27),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_175),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_198),
.Y(n_208)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_196),
.C(n_203),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_192),
.A2(n_194),
.B1(n_197),
.B2(n_200),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_176),
.A2(n_153),
.B1(n_164),
.B2(n_159),
.Y(n_194)
);

INVxp33_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_SL g212 ( 
.A(n_195),
.B(n_168),
.C(n_178),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_156),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_152),
.B1(n_157),
.B2(n_160),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_174),
.A2(n_150),
.B1(n_161),
.B2(n_155),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_141),
.C(n_59),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_204),
.A2(n_28),
.B(n_32),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_27),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_182),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_26),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_191),
.A2(n_177),
.B1(n_170),
.B2(n_166),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_201),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_179),
.C(n_185),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_216),
.C(n_220),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_212),
.A2(n_218),
.B1(n_217),
.B2(n_195),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_171),
.B(n_187),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_199),
.B(n_192),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_218),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_196),
.C(n_197),
.Y(n_216)
);

NOR3xp33_ASAP7_75t_SL g218 ( 
.A(n_205),
.B(n_167),
.C(n_173),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_183),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_221),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_184),
.C(n_29),
.Y(n_220)
);

NOR2xp67_ASAP7_75t_R g222 ( 
.A(n_205),
.B(n_27),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_206),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_223),
.A2(n_204),
.B(n_20),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_233),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_227),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_228),
.A2(n_1),
.B(n_3),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_20),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_201),
.C(n_189),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_235),
.C(n_220),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_231),
.B(n_209),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_214),
.A2(n_198),
.B1(n_2),
.B2(n_3),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_232),
.A2(n_208),
.B1(n_3),
.B2(n_4),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_210),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_26),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_5),
.Y(n_253)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_221),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_242),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_241),
.B(n_242),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_243),
.B(n_244),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_245),
.A2(n_235),
.B1(n_225),
.B2(n_6),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_224),
.B(n_225),
.C(n_233),
.Y(n_246)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_250),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_4),
.Y(n_250)
);

OAI21x1_ASAP7_75t_L g255 ( 
.A1(n_252),
.A2(n_241),
.B(n_245),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_5),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_256),
.Y(n_261)
);

OAI21x1_ASAP7_75t_L g260 ( 
.A1(n_255),
.A2(n_248),
.B(n_7),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_5),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_6),
.Y(n_257)
);

O2A1O1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_248),
.B(n_8),
.C(n_10),
.Y(n_262)
);

AO21x1_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_262),
.B(n_258),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_259),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_263),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_265),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_258),
.C(n_11),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_10),
.C(n_11),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_267),
.B(n_268),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_12),
.C(n_267),
.Y(n_270)
);


endmodule