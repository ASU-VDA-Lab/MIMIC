module real_jpeg_15994_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_10;
wire n_9;
wire n_12;
wire n_11;
wire n_14;
wire n_18;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx6p67_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_R g11 ( 
.A(n_1),
.B(n_12),
.Y(n_11)
);

AOI21xp33_ASAP7_75t_L g15 ( 
.A1(n_1),
.A2(n_16),
.B(n_20),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_2),
.B(n_5),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_3),
.B(n_6),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g9 ( 
.A(n_4),
.B(n_10),
.Y(n_9)
);

OR2x4_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

AOI221xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_8)
);

INVx2_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_13),
.B(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_19),
.Y(n_17)
);


endmodule