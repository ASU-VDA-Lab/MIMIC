module fake_netlist_1_5636_n_660 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_166, n_162, n_75, n_163, n_105, n_159, n_72, n_136, n_43, n_76, n_89, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_15, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_660);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_166;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_15;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_660;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_387;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_178;
wire n_616;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_524;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_602;
wire n_198;
wire n_424;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_175;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g172 ( .A(n_75), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_145), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_124), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_96), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_102), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_58), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_111), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_52), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_65), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_64), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_117), .Y(n_182) );
INVx1_ASAP7_75t_SL g183 ( .A(n_19), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_37), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_78), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_23), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_140), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_139), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_10), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_16), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_43), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_18), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_5), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_25), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_55), .Y(n_195) );
NOR2xp67_ASAP7_75t_L g196 ( .A(n_155), .B(n_42), .Y(n_196) );
BUFx5_ASAP7_75t_L g197 ( .A(n_151), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_87), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_32), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_17), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_132), .Y(n_201) );
INVx1_ASAP7_75t_SL g202 ( .A(n_122), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_127), .Y(n_203) );
BUFx5_ASAP7_75t_L g204 ( .A(n_48), .Y(n_204) );
CKINVDCx14_ASAP7_75t_R g205 ( .A(n_70), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g206 ( .A(n_56), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_118), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_60), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_92), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_156), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_125), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_138), .Y(n_212) );
BUFx3_ASAP7_75t_L g213 ( .A(n_159), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_51), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_153), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_57), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_150), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_149), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_129), .Y(n_219) );
CKINVDCx16_ASAP7_75t_R g220 ( .A(n_123), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_40), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_164), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_120), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_135), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_126), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_147), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_90), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_163), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_131), .Y(n_229) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_20), .Y(n_230) );
CKINVDCx16_ASAP7_75t_R g231 ( .A(n_171), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_13), .Y(n_232) );
INVxp67_ASAP7_75t_L g233 ( .A(n_116), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_146), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_137), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_26), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_38), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_165), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_1), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_68), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_130), .Y(n_241) );
INVxp67_ASAP7_75t_L g242 ( .A(n_72), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_133), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_128), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_115), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_157), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_80), .Y(n_247) );
BUFx10_ASAP7_75t_L g248 ( .A(n_47), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_21), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_134), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_99), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_152), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_73), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_112), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_3), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_154), .Y(n_256) );
OR2x2_ASAP7_75t_L g257 ( .A(n_148), .B(n_161), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_142), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_158), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_15), .Y(n_260) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_106), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_114), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_35), .Y(n_263) );
BUFx5_ASAP7_75t_L g264 ( .A(n_143), .Y(n_264) );
CKINVDCx16_ASAP7_75t_R g265 ( .A(n_162), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_121), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_39), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_101), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_14), .Y(n_269) );
INVx1_ASAP7_75t_SL g270 ( .A(n_50), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_71), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_30), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_41), .Y(n_273) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_141), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_119), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_160), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_136), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_144), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_193), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_255), .Y(n_280) );
BUFx12f_ASAP7_75t_L g281 ( .A(n_248), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_197), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_227), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_230), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_197), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_190), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_258), .B(n_0), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_229), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_206), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_197), .Y(n_290) );
INVx4_ASAP7_75t_L g291 ( .A(n_176), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_248), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_172), .Y(n_293) );
BUFx8_ASAP7_75t_L g294 ( .A(n_239), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_220), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_173), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_227), .Y(n_297) );
NAND2xp33_ASAP7_75t_L g298 ( .A(n_197), .B(n_9), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_231), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_174), .Y(n_300) );
NAND3xp33_ASAP7_75t_L g301 ( .A(n_284), .B(n_239), .C(n_205), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_282), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_291), .B(n_265), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_285), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_291), .B(n_178), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_290), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_292), .B(n_179), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_289), .A2(n_261), .B1(n_274), .B2(n_250), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_283), .Y(n_309) );
AND3x2_ASAP7_75t_L g310 ( .A(n_279), .B(n_242), .C(n_233), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_283), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_292), .B(n_180), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_293), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_300), .B(n_181), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_283), .Y(n_315) );
INVxp67_ASAP7_75t_L g316 ( .A(n_308), .Y(n_316) );
BUFx6f_ASAP7_75t_SL g317 ( .A(n_313), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_313), .B(n_280), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_302), .Y(n_319) );
INVxp67_ASAP7_75t_L g320 ( .A(n_303), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_301), .B(n_287), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_305), .B(n_296), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_304), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_306), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_307), .B(n_281), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_314), .B(n_188), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_315), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_312), .A2(n_299), .B1(n_295), .B2(n_298), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_320), .B(n_310), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_322), .A2(n_177), .B(n_175), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_321), .A2(n_184), .B(n_182), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_318), .A2(n_186), .B(n_185), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_324), .B(n_288), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_319), .A2(n_194), .B(n_187), .Y(n_334) );
OAI21xp5_ASAP7_75t_L g335 ( .A1(n_323), .A2(n_199), .B(n_198), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_328), .B(n_286), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_316), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_325), .A2(n_217), .B(n_208), .Y(n_338) );
INVx2_ASAP7_75t_SL g339 ( .A(n_326), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_327), .A2(n_219), .B(n_218), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_328), .A2(n_232), .B(n_226), .Y(n_341) );
AND2x6_ASAP7_75t_L g342 ( .A(n_317), .B(n_234), .Y(n_342) );
NAND2xp33_ASAP7_75t_SL g343 ( .A(n_339), .B(n_317), .Y(n_343) );
AND2x6_ASAP7_75t_L g344 ( .A(n_342), .B(n_235), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g345 ( .A1(n_341), .A2(n_238), .B(n_236), .Y(n_345) );
OA21x2_ASAP7_75t_L g346 ( .A1(n_335), .A2(n_244), .B(n_240), .Y(n_346) );
AOI211x1_ASAP7_75t_L g347 ( .A1(n_332), .A2(n_245), .B(n_260), .C(n_259), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_337), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_333), .B(n_191), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_330), .A2(n_257), .B(n_256), .Y(n_350) );
OAI222xp33_ASAP7_75t_L g351 ( .A1(n_336), .A2(n_277), .B1(n_271), .B2(n_273), .C1(n_246), .C2(n_267), .Y(n_351) );
OAI21xp5_ASAP7_75t_L g352 ( .A1(n_331), .A2(n_278), .B(n_196), .Y(n_352) );
INVx1_ASAP7_75t_SL g353 ( .A(n_342), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_338), .A2(n_195), .B(n_189), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_334), .A2(n_225), .B(n_222), .Y(n_355) );
BUFx10_ASAP7_75t_L g356 ( .A(n_342), .Y(n_356) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_329), .B(n_192), .Y(n_357) );
AO21x1_ASAP7_75t_L g358 ( .A1(n_340), .A2(n_262), .B(n_253), .Y(n_358) );
INVx5_ASAP7_75t_L g359 ( .A(n_342), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_330), .A2(n_202), .B(n_183), .Y(n_360) );
BUFx2_ASAP7_75t_R g361 ( .A(n_329), .Y(n_361) );
OAI22xp33_ASAP7_75t_L g362 ( .A1(n_359), .A2(n_239), .B1(n_200), .B2(n_201), .Y(n_362) );
BUFx2_ASAP7_75t_R g363 ( .A(n_357), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_348), .B(n_294), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_347), .Y(n_365) );
OAI21x1_ASAP7_75t_L g366 ( .A1(n_358), .A2(n_311), .B(n_309), .Y(n_366) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_352), .A2(n_204), .B(n_197), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_344), .A2(n_294), .B1(n_204), .B2(n_264), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_356), .Y(n_369) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_346), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_355), .A2(n_264), .B(n_204), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_359), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_354), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_353), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_359), .B(n_209), .Y(n_375) );
NAND2x1p5_ASAP7_75t_L g376 ( .A(n_344), .B(n_270), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_351), .B(n_203), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_344), .B(n_4), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_343), .Y(n_379) );
BUFx2_ASAP7_75t_L g380 ( .A(n_345), .Y(n_380) );
OA21x2_ASAP7_75t_L g381 ( .A1(n_350), .A2(n_210), .B(n_207), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_361), .Y(n_382) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
OAI21x1_ASAP7_75t_L g384 ( .A1(n_360), .A2(n_264), .B(n_204), .Y(n_384) );
CKINVDCx6p67_ASAP7_75t_R g385 ( .A(n_359), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_359), .A2(n_213), .B1(n_224), .B2(n_275), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_344), .A2(n_247), .B1(n_212), .B2(n_272), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_348), .B(n_5), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_356), .Y(n_389) );
INVx3_ASAP7_75t_SL g390 ( .A(n_359), .Y(n_390) );
NOR2xp67_ASAP7_75t_L g391 ( .A(n_359), .B(n_6), .Y(n_391) );
OA21x2_ASAP7_75t_L g392 ( .A1(n_352), .A2(n_243), .B(n_214), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_348), .Y(n_393) );
OAI21xp5_ASAP7_75t_L g394 ( .A1(n_345), .A2(n_251), .B(n_215), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g395 ( .A1(n_350), .A2(n_276), .B(n_227), .Y(n_395) );
OAI21x1_ASAP7_75t_L g396 ( .A1(n_358), .A2(n_264), .B(n_276), .Y(n_396) );
OAI21xp5_ASAP7_75t_L g397 ( .A1(n_345), .A2(n_252), .B(n_216), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_347), .Y(n_398) );
A2O1A1Ixp33_ASAP7_75t_L g399 ( .A1(n_345), .A2(n_276), .B(n_249), .C(n_269), .Y(n_399) );
OAI22xp5_ASAP7_75t_SL g400 ( .A1(n_348), .A2(n_254), .B1(n_221), .B2(n_223), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_365), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_398), .Y(n_402) );
INVxp67_ASAP7_75t_L g403 ( .A(n_380), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_388), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_393), .Y(n_405) );
OAI21xp5_ASAP7_75t_L g406 ( .A1(n_398), .A2(n_263), .B(n_228), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_373), .B(n_6), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_370), .A2(n_297), .B(n_268), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_384), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_391), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
INVx3_ASAP7_75t_L g412 ( .A(n_385), .Y(n_412) );
BUFx2_ASAP7_75t_L g413 ( .A(n_379), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_364), .B(n_7), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_378), .B(n_7), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_383), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_383), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_383), .Y(n_418) );
BUFx3_ASAP7_75t_L g419 ( .A(n_390), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_374), .Y(n_420) );
INVx2_ASAP7_75t_SL g421 ( .A(n_369), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_375), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_382), .B(n_8), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_396), .Y(n_424) );
AO21x1_ASAP7_75t_SL g425 ( .A1(n_368), .A2(n_8), .B(n_11), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_366), .Y(n_426) );
AOI211xp5_ASAP7_75t_L g427 ( .A1(n_377), .A2(n_266), .B(n_241), .C(n_237), .Y(n_427) );
INVx4_ASAP7_75t_L g428 ( .A(n_389), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_375), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_367), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_371), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_372), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_381), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_381), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_392), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_392), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_394), .Y(n_437) );
NOR2x1_ASAP7_75t_SL g438 ( .A(n_386), .B(n_297), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_400), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_397), .A2(n_211), .B1(n_297), .B2(n_24), .Y(n_440) );
OAI21x1_ASAP7_75t_L g441 ( .A1(n_395), .A2(n_12), .B(n_22), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_387), .B(n_27), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_363), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_399), .A2(n_170), .B1(n_29), .B2(n_31), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_362), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_388), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_398), .B(n_28), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_398), .B(n_33), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_388), .Y(n_449) );
NAND3xp33_ASAP7_75t_SL g450 ( .A(n_376), .B(n_34), .C(n_36), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_388), .Y(n_451) );
OAI222xp33_ASAP7_75t_L g452 ( .A1(n_380), .A2(n_44), .B1(n_45), .B2(n_46), .C1(n_49), .C2(n_53), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_372), .B(n_54), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_385), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_365), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_365), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_365), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_365), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_365), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_365), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_365), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_365), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_404), .B(n_59), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_405), .B(n_61), .Y(n_464) );
INVx2_ASAP7_75t_SL g465 ( .A(n_419), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_403), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_403), .B(n_62), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_420), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_402), .Y(n_469) );
INVxp67_ASAP7_75t_SL g470 ( .A(n_407), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_414), .B(n_63), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_446), .B(n_66), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_432), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_449), .B(n_67), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_401), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_455), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_451), .B(n_69), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_419), .B(n_74), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_411), .B(n_76), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_456), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_457), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_458), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_413), .B(n_77), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_459), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_416), .B(n_79), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_460), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_417), .B(n_81), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_461), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_418), .B(n_82), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_439), .B(n_83), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_415), .B(n_84), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_423), .B(n_85), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_435), .Y(n_493) );
BUFx3_ASAP7_75t_L g494 ( .A(n_412), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_422), .B(n_86), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_429), .B(n_169), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_443), .B(n_88), .Y(n_497) );
INVxp67_ASAP7_75t_L g498 ( .A(n_433), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_462), .B(n_168), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_447), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_447), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_448), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_448), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_409), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_437), .A2(n_89), .B1(n_91), .B2(n_93), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_407), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_412), .B(n_94), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_454), .B(n_95), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_445), .B(n_167), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_436), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_426), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_424), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_454), .B(n_97), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_430), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_437), .B(n_166), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_434), .Y(n_516) );
BUFx3_ASAP7_75t_L g517 ( .A(n_428), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_445), .B(n_98), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_410), .B(n_442), .Y(n_519) );
INVxp67_ASAP7_75t_SL g520 ( .A(n_453), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_431), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_450), .A2(n_100), .B1(n_103), .B2(n_104), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_453), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_469), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_466), .B(n_421), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_465), .B(n_425), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_468), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_466), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_476), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_465), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_519), .B(n_408), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_473), .B(n_408), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_481), .B(n_428), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_506), .B(n_427), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_484), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_488), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_469), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_518), .B(n_438), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_520), .B(n_441), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_517), .B(n_406), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_517), .B(n_406), .Y(n_541) );
AND2x4_ASAP7_75t_SL g542 ( .A(n_478), .B(n_440), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_475), .B(n_440), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_500), .B(n_427), .Y(n_544) );
BUFx2_ASAP7_75t_L g545 ( .A(n_494), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_475), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_480), .Y(n_547) );
NOR2xp67_ASAP7_75t_L g548 ( .A(n_494), .B(n_450), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_480), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_482), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_486), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_486), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_501), .B(n_444), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_516), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_520), .B(n_105), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_470), .B(n_444), .Y(n_556) );
INVx4_ASAP7_75t_L g557 ( .A(n_467), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_516), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_498), .Y(n_559) );
INVxp67_ASAP7_75t_SL g560 ( .A(n_493), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_470), .B(n_107), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_493), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_502), .B(n_108), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_498), .Y(n_564) );
AND2x6_ASAP7_75t_L g565 ( .A(n_523), .B(n_503), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_483), .B(n_109), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_510), .B(n_110), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_528), .B(n_510), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_527), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_529), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_530), .B(n_490), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_525), .B(n_497), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_560), .B(n_521), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_536), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_537), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_535), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_562), .B(n_521), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_554), .B(n_504), .Y(n_578) );
INVx3_ASAP7_75t_L g579 ( .A(n_545), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_559), .Y(n_580) );
AND2x4_ASAP7_75t_L g581 ( .A(n_558), .B(n_504), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_533), .B(n_531), .Y(n_582) );
AND2x2_ASAP7_75t_SL g583 ( .A(n_542), .B(n_557), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_559), .B(n_514), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_564), .Y(n_585) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_564), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_540), .B(n_492), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_541), .B(n_464), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_546), .B(n_471), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_524), .B(n_514), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_524), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_547), .B(n_511), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_549), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_550), .B(n_511), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_551), .B(n_512), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_552), .B(n_509), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_586), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_569), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_575), .B(n_556), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_582), .B(n_526), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_570), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_580), .B(n_532), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_585), .B(n_553), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_573), .B(n_567), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_574), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_577), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_579), .B(n_538), .Y(n_607) );
INVx2_ASAP7_75t_SL g608 ( .A(n_579), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_568), .B(n_557), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_583), .B(n_548), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_576), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_591), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_572), .B(n_534), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_593), .Y(n_614) );
INVx2_ASAP7_75t_SL g615 ( .A(n_608), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_610), .A2(n_587), .B1(n_588), .B2(n_571), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_599), .B(n_578), .Y(n_617) );
INVx1_ASAP7_75t_SL g618 ( .A(n_609), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_607), .B(n_555), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_597), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_597), .B(n_596), .Y(n_621) );
NOR2xp33_ASAP7_75t_SL g622 ( .A(n_600), .B(n_589), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_604), .A2(n_555), .B1(n_561), .B2(n_544), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_613), .A2(n_505), .B1(n_563), .B2(n_594), .Y(n_624) );
NOR2x1_ASAP7_75t_L g625 ( .A(n_611), .B(n_515), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_624), .A2(n_602), .B1(n_606), .B2(n_603), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_616), .A2(n_565), .B1(n_605), .B2(n_601), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_620), .B(n_614), .Y(n_628) );
INVxp67_ASAP7_75t_L g629 ( .A(n_615), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_617), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_621), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_618), .A2(n_598), .B1(n_612), .B2(n_584), .C(n_581), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_626), .A2(n_625), .B(n_622), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_628), .Y(n_634) );
AOI21xp33_ASAP7_75t_L g635 ( .A1(n_629), .A2(n_623), .B(n_507), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_627), .A2(n_619), .B1(n_584), .B2(n_539), .Y(n_636) );
OAI221xp5_ASAP7_75t_SL g637 ( .A1(n_632), .A2(n_491), .B1(n_513), .B2(n_508), .C(n_566), .Y(n_637) );
NOR2x1_ASAP7_75t_L g638 ( .A(n_633), .B(n_452), .Y(n_638) );
NOR3x1_ASAP7_75t_L g639 ( .A(n_636), .B(n_631), .C(n_630), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_637), .B(n_452), .C(n_505), .Y(n_640) );
NOR2x1_ASAP7_75t_L g641 ( .A(n_638), .B(n_634), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_640), .A2(n_635), .B(n_463), .Y(n_642) );
NOR3xp33_ASAP7_75t_L g643 ( .A(n_639), .B(n_479), .C(n_474), .Y(n_643) );
NOR2x1_ASAP7_75t_L g644 ( .A(n_641), .B(n_472), .Y(n_644) );
NOR2xp67_ASAP7_75t_L g645 ( .A(n_642), .B(n_113), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_645), .A2(n_643), .B1(n_522), .B2(n_539), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_644), .B(n_581), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_647), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_646), .B(n_477), .Y(n_649) );
INVx3_ASAP7_75t_SL g650 ( .A(n_648), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_649), .Y(n_651) );
INVxp33_ASAP7_75t_L g652 ( .A(n_651), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_650), .B(n_565), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_652), .B(n_522), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_653), .Y(n_655) );
AOI22xp33_ASAP7_75t_SL g656 ( .A1(n_655), .A2(n_495), .B1(n_565), .B2(n_489), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_654), .A2(n_565), .B1(n_487), .B2(n_496), .Y(n_657) );
NAND3xp33_ASAP7_75t_L g658 ( .A(n_657), .B(n_499), .C(n_485), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_658), .A2(n_656), .B1(n_543), .B2(n_592), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_659), .A2(n_595), .B1(n_592), .B2(n_590), .Y(n_660) );
endmodule