module fake_jpeg_17786_n_83 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_83);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_83;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_5),
.B(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_0),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_28),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_15),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_13),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_34),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_23),
.B1(n_12),
.B2(n_13),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_24),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_1),
.B1(n_10),
.B2(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_4),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_16),
.B1(n_17),
.B2(n_1),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_37),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_41),
.B1(n_7),
.B2(n_44),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_24),
.C(n_39),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_63),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_29),
.B1(n_46),
.B2(n_4),
.Y(n_60)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_57),
.C(n_50),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_58),
.C(n_51),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_62),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_64),
.B(n_16),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_65),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_68),
.A2(n_64),
.B1(n_53),
.B2(n_37),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_61),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_72),
.Y(n_77)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_70),
.B(n_69),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_70),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_SL g81 ( 
.A(n_78),
.B(n_30),
.C(n_74),
.Y(n_81)
);

OAI31xp33_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_77),
.A3(n_71),
.B(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_80),
.B(n_81),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_30),
.Y(n_83)
);


endmodule