module fake_jpeg_17088_n_236 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_8),
.B(n_2),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

CKINVDCx6p67_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_34),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_26),
.B1(n_30),
.B2(n_18),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_45),
.A2(n_57),
.B1(n_62),
.B2(n_29),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_26),
.B1(n_30),
.B2(n_18),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_55),
.B1(n_59),
.B2(n_35),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_43),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_54),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_18),
.B(n_32),
.C(n_28),
.Y(n_49)
);

OAI32xp33_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_23),
.A3(n_19),
.B1(n_29),
.B2(n_33),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_30),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_27),
.B1(n_28),
.B2(n_32),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_34),
.B1(n_17),
.B2(n_21),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_29),
.B1(n_19),
.B2(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_13),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_1),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_61),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_17),
.B1(n_21),
.B2(n_20),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_1),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_61),
.Y(n_78)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_65),
.B(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_78),
.Y(n_92)
);

BUFx2_ASAP7_75t_SL g68 ( 
.A(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_68),
.Y(n_112)
);

AO22x1_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_35),
.B1(n_37),
.B2(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_22),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_71),
.B(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_22),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_72),
.B(n_81),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_77),
.Y(n_100)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_63),
.B(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_80),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_22),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_10),
.B(n_16),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_40),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_51),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_90),
.B(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_91),
.B(n_83),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_40),
.C(n_38),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_103),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_99),
.B(n_75),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_69),
.B1(n_3),
.B2(n_4),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_61),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_67),
.B(n_66),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_63),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_104),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_38),
.C(n_49),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_29),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_19),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_111),
.B(n_73),
.Y(n_122)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_96),
.A2(n_77),
.B1(n_86),
.B2(n_85),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_115),
.A2(n_120),
.B1(n_124),
.B2(n_130),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_126),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_118),
.B(n_122),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_109),
.B(n_82),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_119),
.B(n_125),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_112),
.A2(n_51),
.B1(n_64),
.B2(n_76),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_105),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_134),
.B(n_110),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_74),
.B1(n_69),
.B2(n_19),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_88),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_127),
.B(n_129),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_103),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_89),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_92),
.A2(n_52),
.B1(n_53),
.B2(n_6),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_97),
.A2(n_52),
.B1(n_53),
.B2(n_88),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_133),
.B1(n_93),
.B2(n_94),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_97),
.A2(n_52),
.B1(n_53),
.B2(n_24),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_24),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_115),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_141),
.B(n_143),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_95),
.B(n_92),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_137),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_142),
.B(n_156),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_99),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_150),
.C(n_155),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_102),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_117),
.Y(n_163)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_136),
.A2(n_92),
.B(n_98),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_160),
.B1(n_108),
.B2(n_33),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_104),
.C(n_98),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_107),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_156),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_171),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_139),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_129),
.B1(n_118),
.B2(n_133),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_164),
.A2(n_173),
.B1(n_141),
.B2(n_155),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_116),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_153),
.B(n_157),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_177),
.C(n_143),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_113),
.Y(n_169)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_146),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_172),
.B(n_147),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_148),
.A2(n_134),
.B1(n_125),
.B2(n_94),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_149),
.B1(n_146),
.B2(n_160),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_24),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_16),
.C(n_14),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_14),
.C(n_12),
.Y(n_182)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_187),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_169),
.B(n_140),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_183),
.B(n_188),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_179),
.C(n_167),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_191),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_166),
.A2(n_150),
.B1(n_138),
.B2(n_6),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_193),
.B1(n_162),
.B2(n_7),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_197),
.C(n_184),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_179),
.C(n_177),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_204),
.B1(n_193),
.B2(n_175),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_186),
.B(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_192),
.B(n_170),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_201),
.Y(n_213)
);

INVx11_ASAP7_75t_L g204 ( 
.A(n_194),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_167),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_209),
.C(n_211),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_168),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_199),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_191),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_202),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_215),
.C(n_203),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_206),
.A2(n_174),
.B1(n_185),
.B2(n_190),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_2),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_208),
.B(n_195),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_217),
.B(n_218),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_213),
.A2(n_206),
.B(n_205),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_220),
.A2(n_198),
.B(n_204),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_222),
.C(n_209),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_203),
.C(n_181),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_226),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_207),
.C(n_8),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_219),
.B(n_165),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_9),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_231),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_230),
.Y(n_232)
);

OAI21x1_ASAP7_75t_L g231 ( 
.A1(n_224),
.A2(n_7),
.B(n_8),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_234),
.A2(n_228),
.B(n_232),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_7),
.Y(n_236)
);


endmodule