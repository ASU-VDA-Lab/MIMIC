module real_jpeg_4935_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_0),
.A2(n_37),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_0),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_0),
.A2(n_248),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_0),
.A2(n_76),
.B1(n_248),
.B2(n_331),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_0),
.A2(n_132),
.B1(n_248),
.B2(n_428),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_1),
.A2(n_118),
.B1(n_195),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_1),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_1),
.B(n_270),
.C(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_1),
.B(n_114),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_1),
.B(n_177),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_1),
.B(n_90),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_1),
.B(n_341),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_2),
.A2(n_35),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_2),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_2),
.A2(n_77),
.B1(n_202),
.B2(n_266),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_2),
.A2(n_86),
.B1(n_178),
.B2(n_202),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_2),
.A2(n_202),
.B1(n_346),
.B2(n_348),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_3),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_3),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_3),
.Y(n_231)
);

INVx8_ASAP7_75t_L g319 ( 
.A(n_3),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_4),
.Y(n_151)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_4),
.Y(n_250)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_4),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_5),
.A2(n_112),
.B1(n_132),
.B2(n_134),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_5),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_5),
.A2(n_68),
.B1(n_134),
.B2(n_160),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_5),
.A2(n_134),
.B1(n_222),
.B2(n_226),
.Y(n_221)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g401 ( 
.A(n_6),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_7),
.A2(n_195),
.B1(n_288),
.B2(n_290),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_7),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_7),
.A2(n_290),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_7),
.A2(n_290),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_7),
.A2(n_34),
.B1(n_290),
.B2(n_456),
.Y(n_455)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_8),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_9),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_9),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_9),
.A2(n_34),
.B1(n_127),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_9),
.A2(n_127),
.B1(n_191),
.B2(n_194),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_9),
.A2(n_127),
.B1(n_277),
.B2(n_298),
.Y(n_413)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_11),
.A2(n_36),
.B1(n_58),
.B2(n_61),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_11),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_11),
.A2(n_61),
.B1(n_133),
.B2(n_167),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_11),
.A2(n_61),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_11),
.A2(n_61),
.B1(n_183),
.B2(n_277),
.Y(n_386)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_13),
.A2(n_36),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_13),
.A2(n_52),
.B1(n_240),
.B2(n_244),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_13),
.A2(n_52),
.B1(n_226),
.B2(n_353),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g431 ( 
.A1(n_13),
.A2(n_52),
.B1(n_432),
.B2(n_435),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_14),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_14),
.Y(n_186)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_14),
.Y(n_225)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_15),
.Y(n_104)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_17),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_18),
.A2(n_92),
.B1(n_94),
.B2(n_98),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_18),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_18),
.A2(n_98),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_18),
.A2(n_98),
.B1(n_183),
.B2(n_187),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_503),
.B(n_506),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_206),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_205),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_153),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_24),
.B(n_153),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_135),
.B2(n_136),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_62),
.C(n_99),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_27),
.A2(n_137),
.B1(n_138),
.B2(n_152),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_27),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_27),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_50),
.B1(n_55),
.B2(n_57),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_28),
.A2(n_55),
.B1(n_57),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_28),
.A2(n_247),
.B(n_251),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_28),
.A2(n_55),
.B1(n_247),
.B2(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_29),
.B(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_29),
.A2(n_420),
.B(n_424),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_40),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_41),
.B1(n_44),
.B2(n_48),
.Y(n_40)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g405 ( 
.A(n_35),
.Y(n_405)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_42),
.B(n_337),
.Y(n_402)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_45),
.Y(n_347)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_46),
.Y(n_343)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_47),
.Y(n_133)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_47),
.Y(n_338)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_49),
.Y(n_146)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_49),
.Y(n_169)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_49),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_51),
.B(n_56),
.Y(n_199)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_55),
.B(n_263),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_55),
.A2(n_200),
.B(n_455),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_56),
.B(n_201),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_62),
.A2(n_63),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_62),
.A2(n_63),
.B1(n_99),
.B2(n_100),
.Y(n_155)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_89),
.B(n_91),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_64),
.A2(n_262),
.B(n_264),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_64),
.A2(n_89),
.B1(n_287),
.B2(n_330),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_64),
.A2(n_264),
.B(n_330),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_64),
.A2(n_89),
.B1(n_431),
.B2(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_65),
.A2(n_90),
.B1(n_159),
.B2(n_162),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_65),
.A2(n_90),
.B1(n_159),
.B2(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_65),
.A2(n_90),
.B1(n_190),
.B2(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_65),
.B(n_265),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_79),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_71),
.B1(n_74),
.B2(n_76),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_68),
.B(n_269),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_69),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_69),
.Y(n_437)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_70),
.Y(n_237)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_70),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_70),
.Y(n_364)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_73),
.Y(n_270)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_79),
.A2(n_287),
.B(n_291),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_86),
.B2(n_88),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_85),
.Y(n_353)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_89),
.A2(n_291),
.B(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_90),
.B(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_93),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_122),
.B1(n_130),
.B2(n_131),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_101),
.A2(n_130),
.B1(n_131),
.B2(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_101),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_101),
.A2(n_130),
.B1(n_166),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_101),
.A2(n_130),
.B1(n_378),
.B2(n_427),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_114),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_105),
.B1(n_108),
.B2(n_112),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_107),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_107),
.Y(n_245)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_112),
.Y(n_380)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_114),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_114),
.A2(n_123),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

AOI22x1_ASAP7_75t_L g458 ( 
.A1(n_114),
.A2(n_164),
.B1(n_382),
.B2(n_459),
.Y(n_458)
);

AO22x2_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_114)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_117),
.Y(n_361)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_126),
.Y(n_348)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_130),
.B(n_345),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_130),
.A2(n_378),
.B(n_381),
.Y(n_377)
);

INVx6_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_147),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_144),
.Y(n_379)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_151),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_170),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_154),
.B(n_157),
.CI(n_170),
.CON(n_208),
.SN(n_208)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_157),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_163),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_158),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_164),
.A2(n_335),
.B(n_344),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_164),
.B(n_382),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_164),
.A2(n_344),
.B(n_475),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g395 ( 
.A1(n_167),
.A2(n_396),
.A3(n_399),
.B1(n_402),
.B2(n_403),
.Y(n_395)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B(n_198),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_189),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_172),
.A2(n_198),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_172),
.A2(n_189),
.B1(n_214),
.B2(n_446),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_181),
.B(n_182),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_173),
.A2(n_182),
.B1(n_221),
.B2(n_229),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_173),
.A2(n_275),
.B(n_280),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_173),
.A2(n_263),
.B(n_280),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_173),
.A2(n_408),
.B1(n_409),
.B2(n_412),
.Y(n_407)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_174),
.B(n_283),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_174),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_174),
.A2(n_176),
.B1(n_352),
.B2(n_386),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_174),
.A2(n_281),
.B1(n_413),
.B2(n_452),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

INVx3_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_177),
.Y(n_282)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_185),
.Y(n_276)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx8_ASAP7_75t_L g188 ( 
.A(n_186),
.Y(n_188)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_186),
.Y(n_308)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_187),
.Y(n_298)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_189),
.Y(n_446)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI32xp33_ASAP7_75t_L g354 ( 
.A1(n_192),
.A2(n_340),
.A3(n_355),
.B1(n_359),
.B2(n_362),
.Y(n_354)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_193),
.Y(n_289)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_198),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_252),
.B(n_502),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_208),
.B(n_209),
.Y(n_502)
);

BUFx24_ASAP7_75t_SL g510 ( 
.A(n_208),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.C(n_218),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_210),
.A2(n_211),
.B1(n_215),
.B2(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_215),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_218),
.B(n_461),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_238),
.C(n_246),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_219),
.B(n_444),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_232),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_220),
.B(n_232),
.Y(n_469)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_221),
.Y(n_452)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_225),
.Y(n_272)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_226),
.Y(n_304)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_229),
.A2(n_303),
.B(n_309),
.Y(n_302)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_233),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_234),
.Y(n_332)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_237),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_238),
.B(n_246),
.Y(n_444)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_239),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx5_ASAP7_75t_L g358 ( 
.A(n_245),
.Y(n_358)
);

INVx8_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_251),
.Y(n_424)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI311xp33_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_440),
.A3(n_478),
.B1(n_496),
.C1(n_497),
.Y(n_254)
);

AOI21x1_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_389),
.B(n_439),
.Y(n_255)
);

AO21x1_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_369),
.B(n_388),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_324),
.B(n_368),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_294),
.B(n_323),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_273),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_260),
.B(n_273),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_267),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_261),
.A2(n_267),
.B1(n_268),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_261),
.Y(n_321)
);

OAI21xp33_ASAP7_75t_SL g335 ( 
.A1(n_263),
.A2(n_336),
.B(n_339),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_263),
.B(n_404),
.Y(n_403)
);

OAI21xp33_ASAP7_75t_SL g420 ( 
.A1(n_263),
.A2(n_403),
.B(n_421),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_272),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_284),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_274),
.B(n_285),
.C(n_293),
.Y(n_325)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_282),
.A2(n_309),
.B(n_351),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_292),
.B2(n_293),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_312),
.B(n_322),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_301),
.B(n_311),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_310),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_310),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_320),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_320),
.Y(n_322)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx8_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_319),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_325),
.B(n_326),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_349),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_333),
.B2(n_334),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_329),
.B(n_333),
.C(n_349),
.Y(n_370)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_345),
.Y(n_382)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_354),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_350),
.B(n_354),
.Y(n_375)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx6_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx8_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx6_ASAP7_75t_L g367 ( 
.A(n_361),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_365),
.Y(n_362)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_370),
.B(n_371),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_373),
.B1(n_376),
.B2(n_387),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_375),
.C(n_387),
.Y(n_390)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_376),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_383),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_377),
.B(n_384),
.C(n_385),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_386),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_390),
.B(n_391),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_417),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_392)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_393),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_395),
.B1(n_406),
.B2(n_407),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_395),
.B(n_406),
.Y(n_473)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_398),
.Y(n_423)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx8_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_414),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_414),
.B(n_415),
.C(n_417),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_419),
.B1(n_425),
.B2(n_438),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_418),
.B(n_426),
.C(n_430),
.Y(n_487)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_425),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_430),
.Y(n_425)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_427),
.Y(n_475)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

NAND2xp33_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_463),
.Y(n_440)
);

A2O1A1Ixp33_ASAP7_75t_SL g497 ( 
.A1(n_441),
.A2(n_463),
.B(n_498),
.C(n_501),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_460),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_442),
.B(n_460),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_445),
.C(n_447),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_443),
.B(n_445),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_447),
.B(n_477),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_453),
.C(n_458),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_449),
.B(n_451),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_449),
.B(n_451),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_453),
.A2(n_454),
.B1(n_458),
.B2(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_458),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_476),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_464),
.B(n_476),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_469),
.C(n_470),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_465),
.A2(n_466),
.B1(n_469),
.B2(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_469),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_489),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_473),
.C(n_474),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_471),
.A2(n_472),
.B1(n_474),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_473),
.B(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_474),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_479),
.B(n_491),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_480),
.A2(n_499),
.B(n_500),
.Y(n_498)
);

NOR2x1_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_488),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_481),
.B(n_488),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_485),
.C(n_487),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_494),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_485),
.A2(n_486),
.B1(n_487),
.B2(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_487),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_492),
.B(n_493),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g507 ( 
.A(n_504),
.Y(n_507)
);

INVx13_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.Y(n_506)
);


endmodule