module fake_jpeg_27123_n_103 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx24_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_25),
.Y(n_28)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_27),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_11),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_11),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_19),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_27),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_22),
.B1(n_26),
.B2(n_16),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_46),
.B1(n_30),
.B2(n_29),
.Y(n_59)
);

BUFx24_ASAP7_75t_SL g37 ( 
.A(n_34),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_13),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_10),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_16),
.Y(n_45)
);

AO22x1_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_32),
.B1(n_33),
.B2(n_24),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_35),
.B(n_17),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_55),
.Y(n_63)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

OAI22x1_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_14),
.B1(n_20),
.B2(n_32),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_60),
.B(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVxp67_ASAP7_75t_SL g74 ( 
.A(n_67),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_41),
.C(n_29),
.Y(n_71)
);

A2O1A1O1Ixp25_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_47),
.B(n_56),
.C(n_55),
.D(n_50),
.Y(n_72)
);

AOI221xp5_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.C(n_4),
.Y(n_87)
);

OAI32xp33_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_56),
.A3(n_48),
.B1(n_59),
.B2(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_58),
.B(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_76),
.B(n_77),
.Y(n_82)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_14),
.C(n_20),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_62),
.C(n_66),
.Y(n_84)
);

AOI321xp33_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_68),
.A3(n_70),
.B1(n_65),
.B2(n_51),
.C(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_80),
.B(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_74),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_87),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_18),
.C(n_15),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_91),
.B(n_92),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_75),
.Y(n_92)
);

XNOR2x2_ASAP7_75t_SL g94 ( 
.A(n_88),
.B(n_15),
.Y(n_94)
);

HAxp5_ASAP7_75t_SL g95 ( 
.A(n_94),
.B(n_90),
.CON(n_95),
.SN(n_95)
);

AOI31xp33_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_4),
.A3(n_5),
.B(n_7),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_1),
.B(n_2),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_97)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_97),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_9),
.Y(n_99)
);

INVxp33_ASAP7_75t_SL g101 ( 
.A(n_99),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_100),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);


endmodule