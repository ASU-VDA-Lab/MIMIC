module fake_jpeg_20813_n_201 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_7),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_39),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_28),
.B1(n_29),
.B2(n_23),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_53),
.B1(n_36),
.B2(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_21),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_35),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_28),
.B1(n_29),
.B2(n_23),
.Y(n_53)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_24),
.B(n_20),
.C(n_22),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_27),
.B(n_30),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_41),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_49),
.B(n_20),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_60),
.B(n_67),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_36),
.B1(n_28),
.B2(n_35),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_71),
.B1(n_75),
.B2(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_70),
.Y(n_88)
);

BUFx4f_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_50),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_24),
.B1(n_21),
.B2(n_18),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_18),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_73),
.Y(n_89)
);

AOI32xp33_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_22),
.A3(n_23),
.B1(n_15),
.B2(n_27),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_35),
.B1(n_33),
.B2(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_27),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_19),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_90),
.B1(n_94),
.B2(n_99),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_84),
.B(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_43),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_43),
.B1(n_46),
.B2(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_56),
.B(n_13),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_97),
.Y(n_118)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_34),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_55),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_75),
.A2(n_46),
.B1(n_33),
.B2(n_31),
.Y(n_99)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_111),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_64),
.C(n_38),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_99),
.C(n_87),
.Y(n_129)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_76),
.B1(n_68),
.B2(n_46),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_107),
.B1(n_112),
.B2(n_113),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_33),
.B1(n_54),
.B2(n_48),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_121),
.Y(n_124)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_58),
.B1(n_66),
.B2(n_69),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_81),
.A2(n_69),
.B1(n_34),
.B2(n_61),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_91),
.B(n_98),
.Y(n_132)
);

AOI322xp5_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_12),
.A3(n_11),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_91),
.Y(n_134)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_89),
.A2(n_38),
.B1(n_19),
.B2(n_30),
.Y(n_119)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_94),
.A2(n_38),
.B1(n_30),
.B2(n_26),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_103),
.A2(n_94),
.B1(n_87),
.B2(n_79),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_83),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_128),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_88),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_138),
.C(n_120),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_134),
.Y(n_146)
);

AO21x2_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_78),
.B(n_98),
.Y(n_133)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_80),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_141),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_86),
.C(n_26),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_118),
.B(n_11),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_140),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_109),
.B(n_105),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_138),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_101),
.B(n_107),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_113),
.B1(n_111),
.B2(n_86),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_149),
.A2(n_123),
.B1(n_102),
.B2(n_106),
.Y(n_167)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

AOI22x1_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_129),
.B1(n_131),
.B2(n_125),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);

OAI321xp33_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_133),
.A3(n_127),
.B1(n_128),
.B2(n_139),
.C(n_131),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_159),
.A2(n_150),
.B1(n_143),
.B2(n_168),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_144),
.C(n_155),
.Y(n_174)
);

OAI322xp33_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_165),
.B(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_123),
.B1(n_2),
.B2(n_8),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_170),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_174),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_155),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_177),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_162),
.B(n_157),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_153),
.B(n_143),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_153),
.B(n_169),
.Y(n_179)
);

AO22x1_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_182),
.B1(n_171),
.B2(n_166),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_SL g182 ( 
.A1(n_178),
.A2(n_150),
.B(n_149),
.C(n_158),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_172),
.A2(n_163),
.B1(n_164),
.B2(n_160),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_185),
.B(n_167),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_174),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_187),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_175),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_189),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_182),
.C(n_180),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_193),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_188),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_194),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_198),
.B(n_8),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_1),
.Y(n_198)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_199),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_8),
.Y(n_201)
);


endmodule