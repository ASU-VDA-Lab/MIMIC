module fake_jpeg_17726_n_47 (n_3, n_2, n_1, n_0, n_4, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

HAxp5_ASAP7_75t_SL g6 ( 
.A(n_0),
.B(n_1),
.CON(n_6),
.SN(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_0),
.B(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_2),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_14),
.B(n_21),
.Y(n_24)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_16),
.B(n_8),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_6),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_9),
.C(n_12),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_7),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_19),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_23),
.A2(n_14),
.B(n_17),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_12),
.C(n_10),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_28),
.C(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_14),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_12),
.C(n_10),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_32),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_33),
.B1(n_35),
.B2(n_13),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_17),
.C(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_14),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_21),
.B1(n_15),
.B2(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_35),
.A2(n_15),
.B1(n_21),
.B2(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_40),
.Y(n_42)
);

AOI322xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_19),
.A3(n_8),
.B1(n_26),
.B2(n_13),
.C1(n_4),
.C2(n_5),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_36),
.C(n_37),
.Y(n_44)
);

NAND4xp25_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_45),
.C(n_42),
.D(n_36),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_38),
.Y(n_45)
);

AOI21x1_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_41),
.B(n_39),
.Y(n_47)
);


endmodule