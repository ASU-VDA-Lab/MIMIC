module fake_jpeg_17558_n_305 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_305);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_288;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_35),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_19),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_48),
.A2(n_25),
.B1(n_29),
.B2(n_35),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_55),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_21),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_54),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_63),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_36),
.B(n_19),
.C(n_34),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_SL g106 ( 
.A1(n_58),
.A2(n_39),
.B(n_27),
.Y(n_106)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_36),
.B1(n_29),
.B2(n_21),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_48),
.B1(n_53),
.B2(n_25),
.Y(n_88)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_33),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_72),
.Y(n_89)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_35),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_53),
.Y(n_83)
);

CKINVDCx12_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_34),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_75),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_80),
.Y(n_100)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_17),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_37),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_40),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_50),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_103),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_91),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_40),
.B1(n_53),
.B2(n_48),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_88),
.B1(n_92),
.B2(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_56),
.B(n_48),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_38),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_50),
.B1(n_39),
.B2(n_32),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_39),
.B1(n_32),
.B2(n_50),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_28),
.B(n_1),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_78),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_106),
.B1(n_108),
.B2(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_39),
.B1(n_17),
.B2(n_18),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_109),
.B1(n_16),
.B2(n_22),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_81),
.Y(n_130)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_38),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_67),
.A2(n_22),
.B1(n_24),
.B2(n_16),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_113),
.B(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_117),
.A2(n_108),
.B(n_83),
.Y(n_140)
);

BUFx16f_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_128),
.Y(n_144)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_124),
.B1(n_133),
.B2(n_103),
.Y(n_142)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_84),
.B(n_24),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_132),
.Y(n_153)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_131),
.Y(n_143)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_97),
.A2(n_77),
.B1(n_65),
.B2(n_64),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_88),
.B1(n_94),
.B2(n_90),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_92),
.B1(n_99),
.B2(n_89),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_104),
.Y(n_155)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_87),
.A3(n_84),
.B1(n_100),
.B2(n_103),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_127),
.A3(n_125),
.B1(n_120),
.B2(n_104),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_140),
.A2(n_151),
.B(n_162),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_145),
.B1(n_154),
.B2(n_159),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_100),
.B1(n_99),
.B2(n_108),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_116),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_114),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_126),
.A2(n_102),
.B(n_105),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_135),
.A2(n_57),
.B1(n_60),
.B2(n_59),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_152),
.A2(n_161),
.B1(n_69),
.B2(n_61),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_57),
.B1(n_64),
.B2(n_59),
.Y(n_154)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_112),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_30),
.B(n_26),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_158),
.A2(n_167),
.B(n_129),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_60),
.B1(n_85),
.B2(n_81),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_134),
.B1(n_118),
.B2(n_111),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_122),
.A2(n_86),
.B(n_104),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_117),
.B(n_76),
.C(n_52),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_165),
.C(n_28),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_110),
.B(n_28),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_115),
.A2(n_30),
.B(n_26),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_131),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_169),
.A2(n_166),
.B(n_163),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_173),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_174),
.A2(n_176),
.B(n_193),
.Y(n_221)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_149),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_79),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_146),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_188),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_137),
.A2(n_52),
.B1(n_74),
.B2(n_2),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_183),
.A2(n_189),
.B1(n_159),
.B2(n_151),
.Y(n_205)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_28),
.C(n_11),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_192),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_186),
.C(n_194),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_74),
.C(n_52),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_139),
.B(n_28),
.Y(n_187)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_23),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_74),
.B1(n_1),
.B2(n_2),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_161),
.A2(n_23),
.B1(n_20),
.B2(n_2),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_190),
.A2(n_198),
.B1(n_158),
.B2(n_167),
.Y(n_203)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_191),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_154),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_20),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_23),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_196),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_160),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_163),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_156),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_142),
.A2(n_20),
.B1(n_1),
.B2(n_3),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_185),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_183),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_172),
.B1(n_171),
.B2(n_168),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_200),
.A2(n_205),
.B1(n_196),
.B2(n_176),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_164),
.B(n_166),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_212),
.B(n_174),
.Y(n_231)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_152),
.Y(n_216)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_165),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_219),
.C(n_194),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_138),
.C(n_1),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_168),
.A2(n_138),
.B(n_3),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_220),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_178),
.Y(n_223)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_237),
.C(n_238),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_197),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_232),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_180),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_170),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_229),
.B(n_234),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_235),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_170),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_189),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_236),
.A2(n_208),
.B1(n_202),
.B2(n_216),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_190),
.C(n_187),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_195),
.C(n_173),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_198),
.C(n_192),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_219),
.C(n_200),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_240),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_245),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_250),
.C(n_256),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_208),
.B1(n_206),
.B2(n_204),
.Y(n_244)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_220),
.B(n_207),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_239),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_221),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_209),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_251),
.B(n_203),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_204),
.B1(n_202),
.B2(n_201),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_237),
.B1(n_231),
.B2(n_235),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_222),
.A2(n_201),
.B1(n_217),
.B2(n_205),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_255),
.A2(n_182),
.B1(n_191),
.B2(n_4),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_217),
.C(n_221),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_255),
.A2(n_230),
.B(n_226),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_263),
.B(n_267),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_210),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_261),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_210),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_262),
.B(n_264),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_228),
.B(n_223),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_269),
.C(n_253),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_256),
.B(n_213),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_269),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_9),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_260),
.A2(n_243),
.B1(n_246),
.B2(n_241),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_270),
.A2(n_275),
.B1(n_0),
.B2(n_5),
.Y(n_284)
);

OA21x2_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_253),
.B(n_252),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_276),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_9),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_252),
.C(n_3),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_11),
.C(n_13),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_263),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_10),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_277),
.A2(n_266),
.B(n_268),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_289),
.B(n_278),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_284),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_288),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_9),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_276),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_279),
.B(n_275),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_10),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_12),
.B(n_13),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_273),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_272),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_288),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_295),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_296),
.A2(n_298),
.B(n_294),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_290),
.C(n_297),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_291),
.B(n_270),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_301),
.A2(n_271),
.B(n_282),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_271),
.B(n_12),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_0),
.C(n_5),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_13),
.B(n_14),
.Y(n_305)
);


endmodule