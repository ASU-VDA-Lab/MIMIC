module real_aes_1116_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_789;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_0), .B(n_501), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_1), .A2(n_503), .B(n_504), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_2), .B(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_3), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_3), .A2(n_790), .B(n_794), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_4), .Y(n_795) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_5), .B(n_214), .Y(n_538) );
INVx1_ASAP7_75t_L g146 ( .A(n_6), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_7), .B(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_8), .B(n_214), .Y(n_587) );
INVx1_ASAP7_75t_L g184 ( .A(n_9), .Y(n_184) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_10), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_11), .Y(n_152) );
NAND2xp33_ASAP7_75t_L g579 ( .A(n_12), .B(n_211), .Y(n_579) );
INVx2_ASAP7_75t_L g128 ( .A(n_13), .Y(n_128) );
AOI221x1_ASAP7_75t_L g523 ( .A1(n_14), .A2(n_26), .B1(n_501), .B2(n_503), .C(n_524), .Y(n_523) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_15), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_16), .B(n_501), .Y(n_575) );
INVx1_ASAP7_75t_L g212 ( .A(n_17), .Y(n_212) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_18), .A2(n_181), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_19), .B(n_176), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_20), .B(n_214), .Y(n_512) );
AO21x1_ASAP7_75t_L g533 ( .A1(n_21), .A2(n_501), .B(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_SL g103 ( .A(n_22), .B(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g489 ( .A(n_22), .Y(n_489) );
INVx1_ASAP7_75t_L g209 ( .A(n_23), .Y(n_209) );
INVx1_ASAP7_75t_SL g196 ( .A(n_24), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_25), .B(n_139), .Y(n_254) );
AOI33xp33_ASAP7_75t_L g234 ( .A1(n_27), .A2(n_52), .A3(n_132), .B1(n_157), .B2(n_235), .B3(n_236), .Y(n_234) );
NAND2x1_ASAP7_75t_L g554 ( .A(n_28), .B(n_214), .Y(n_554) );
NAND2x1_ASAP7_75t_L g586 ( .A(n_29), .B(n_211), .Y(n_586) );
INVx1_ASAP7_75t_L g137 ( .A(n_30), .Y(n_137) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_31), .A2(n_86), .B(n_128), .Y(n_127) );
OR2x2_ASAP7_75t_L g178 ( .A(n_31), .B(n_86), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_32), .B(n_161), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_33), .B(n_211), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_34), .B(n_214), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_35), .B(n_211), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_36), .A2(n_503), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g145 ( .A(n_37), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g156 ( .A(n_37), .Y(n_156) );
AND2x2_ASAP7_75t_L g165 ( .A(n_37), .B(n_135), .Y(n_165) );
NOR3xp33_ASAP7_75t_L g105 ( .A(n_38), .B(n_106), .C(n_108), .Y(n_105) );
OR2x6_ASAP7_75t_L g487 ( .A(n_38), .B(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_39), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_40), .B(n_501), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_41), .B(n_161), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_42), .A2(n_126), .B1(n_203), .B2(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_43), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_44), .B(n_139), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_45), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_46), .B(n_211), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_47), .B(n_181), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_48), .B(n_139), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_49), .A2(n_503), .B(n_585), .Y(n_584) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_50), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_51), .B(n_211), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_53), .B(n_139), .Y(n_173) );
INVx1_ASAP7_75t_L g133 ( .A(n_54), .Y(n_133) );
INVx1_ASAP7_75t_L g141 ( .A(n_54), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_55), .Y(n_801) );
INVxp33_ASAP7_75t_L g815 ( .A(n_56), .Y(n_815) );
AND2x2_ASAP7_75t_L g175 ( .A(n_57), .B(n_176), .Y(n_175) );
AOI221xp5_ASAP7_75t_L g182 ( .A1(n_58), .A2(n_74), .B1(n_154), .B2(n_161), .C(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_59), .B(n_161), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_60), .B(n_214), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_61), .B(n_126), .Y(n_159) );
AOI21xp5_ASAP7_75t_SL g221 ( .A1(n_62), .A2(n_154), .B(n_222), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_63), .A2(n_503), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g206 ( .A(n_64), .Y(n_206) );
AO21x1_ASAP7_75t_L g535 ( .A1(n_65), .A2(n_503), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_66), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g172 ( .A(n_67), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_68), .B(n_501), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_69), .A2(n_154), .B(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g548 ( .A(n_70), .B(n_177), .Y(n_548) );
INVx1_ASAP7_75t_L g135 ( .A(n_71), .Y(n_135) );
INVx1_ASAP7_75t_L g143 ( .A(n_71), .Y(n_143) );
AND2x2_ASAP7_75t_L g589 ( .A(n_72), .B(n_125), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_73), .B(n_161), .Y(n_237) );
AND2x2_ASAP7_75t_L g198 ( .A(n_75), .B(n_125), .Y(n_198) );
INVx1_ASAP7_75t_L g207 ( .A(n_76), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_77), .A2(n_154), .B(n_195), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_78), .A2(n_154), .B(n_229), .C(n_253), .Y(n_252) );
OAI22xp33_ASAP7_75t_SL g809 ( .A1(n_79), .A2(n_490), .B1(n_792), .B2(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_79), .Y(n_810) );
INVx1_ASAP7_75t_L g104 ( .A(n_80), .Y(n_104) );
AND2x2_ASAP7_75t_L g498 ( .A(n_81), .B(n_125), .Y(n_498) );
AND2x2_ASAP7_75t_SL g219 ( .A(n_82), .B(n_125), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_83), .B(n_501), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_84), .A2(n_154), .B1(n_232), .B2(n_233), .Y(n_231) );
AND2x2_ASAP7_75t_L g534 ( .A(n_85), .B(n_203), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_87), .B(n_211), .Y(n_513) );
AND2x2_ASAP7_75t_L g557 ( .A(n_88), .B(n_125), .Y(n_557) );
INVx1_ASAP7_75t_L g223 ( .A(n_89), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_90), .B(n_214), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_91), .A2(n_503), .B(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_92), .B(n_211), .Y(n_525) );
AND2x2_ASAP7_75t_L g238 ( .A(n_93), .B(n_125), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_94), .B(n_214), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g129 ( .A1(n_95), .A2(n_130), .B(n_136), .C(n_144), .Y(n_129) );
BUFx2_ASAP7_75t_L g806 ( .A(n_96), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_97), .A2(n_503), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_98), .B(n_139), .Y(n_224) );
AOI21xp33_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_109), .B(n_814), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx3_ASAP7_75t_R g816 ( .A(n_101), .Y(n_816) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_105), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_104), .B(n_489), .Y(n_488) );
OR2x6_ASAP7_75t_SL g485 ( .A(n_108), .B(n_486), .Y(n_485) );
AND2x6_ASAP7_75t_SL g788 ( .A(n_108), .B(n_487), .Y(n_788) );
OR2x2_ASAP7_75t_L g798 ( .A(n_108), .B(n_487), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_108), .B(n_486), .Y(n_803) );
AO21x2_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_804), .B(n_807), .Y(n_109) );
OAI211xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_113), .B(n_789), .C(n_799), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
OAI22x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_483), .B1(n_490), .B2(n_785), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
OAI22xp5_ASAP7_75t_SL g790 ( .A1(n_116), .A2(n_791), .B1(n_792), .B2(n_793), .Y(n_790) );
NAND3x1_ASAP7_75t_L g116 ( .A(n_117), .B(n_362), .C(n_429), .Y(n_116) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_322), .Y(n_117) );
NOR3x1_ASAP7_75t_L g118 ( .A(n_119), .B(n_273), .C(n_302), .Y(n_118) );
OAI221xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_187), .B1(n_226), .B2(n_241), .C(n_258), .Y(n_119) );
A2O1A1Ixp33_ASAP7_75t_SL g436 ( .A1(n_120), .A2(n_200), .B(n_437), .C(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_121), .A2(n_408), .B1(n_411), .B2(n_413), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_121), .B(n_227), .Y(n_482) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_166), .Y(n_121) );
BUFx2_ASAP7_75t_L g401 ( .A(n_122), .Y(n_401) );
INVx1_ASAP7_75t_SL g414 ( .A(n_122), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_122), .B(n_269), .Y(n_456) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g239 ( .A(n_123), .B(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g284 ( .A(n_123), .B(n_180), .Y(n_284) );
INVx1_ASAP7_75t_L g295 ( .A(n_123), .Y(n_295) );
INVx2_ASAP7_75t_L g299 ( .A(n_123), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_123), .B(n_270), .Y(n_426) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_149), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_129), .B1(n_147), .B2(n_148), .Y(n_124) );
INVx3_ASAP7_75t_L g148 ( .A(n_125), .Y(n_148) );
INVx4_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_126), .B(n_151), .Y(n_150) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx4f_ASAP7_75t_L g181 ( .A(n_127), .Y(n_181) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_128), .B(n_178), .Y(n_177) );
AND2x4_ASAP7_75t_L g203 ( .A(n_128), .B(n_178), .Y(n_203) );
INVxp67_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_L g171 ( .A1(n_131), .A2(n_172), .B(n_173), .C(n_174), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_SL g183 ( .A1(n_131), .A2(n_174), .B(n_184), .C(n_185), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_SL g195 ( .A1(n_131), .A2(n_174), .B(n_196), .C(n_197), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g205 ( .A1(n_131), .A2(n_138), .B1(n_206), .B2(n_207), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_131), .A2(n_174), .B(n_223), .C(n_224), .Y(n_222) );
INVx2_ASAP7_75t_L g256 ( .A(n_131), .Y(n_256) );
OR2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_134), .Y(n_131) );
AND2x2_ASAP7_75t_L g162 ( .A(n_132), .B(n_163), .Y(n_162) );
INVxp33_ASAP7_75t_L g235 ( .A(n_132), .Y(n_235) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g158 ( .A(n_133), .B(n_146), .Y(n_158) );
AND2x4_ASAP7_75t_L g214 ( .A(n_133), .B(n_142), .Y(n_214) );
INVx3_ASAP7_75t_L g157 ( .A(n_134), .Y(n_157) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x6_ASAP7_75t_L g211 ( .A(n_135), .B(n_140), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g501 ( .A(n_139), .B(n_145), .Y(n_501) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx5_ASAP7_75t_L g174 ( .A(n_145), .Y(n_174) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_146), .Y(n_163) );
AO21x2_ASAP7_75t_L g167 ( .A1(n_148), .A2(n_168), .B(n_175), .Y(n_167) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_148), .A2(n_168), .B(n_175), .Y(n_270) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_148), .A2(n_542), .B(n_548), .Y(n_541) );
AO21x2_ASAP7_75t_L g550 ( .A1(n_148), .A2(n_551), .B(n_557), .Y(n_550) );
AO21x2_ASAP7_75t_L g563 ( .A1(n_148), .A2(n_551), .B(n_557), .Y(n_563) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_148), .A2(n_542), .B(n_548), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_153), .B1(n_159), .B2(n_160), .Y(n_149) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVxp67_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_155), .B(n_158), .Y(n_154) );
NOR2x1p5_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx1_ASAP7_75t_L g236 ( .A(n_157), .Y(n_236) );
AND2x6_ASAP7_75t_L g503 ( .A(n_158), .B(n_165), .Y(n_503) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_162), .B(n_164), .Y(n_161) );
INVx1_ASAP7_75t_L g249 ( .A(n_162), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_164), .Y(n_250) );
BUFx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g375 ( .A(n_166), .B(n_376), .Y(n_375) );
NOR2x1_ASAP7_75t_L g166 ( .A(n_167), .B(n_179), .Y(n_166) );
INVx2_ASAP7_75t_L g278 ( .A(n_167), .Y(n_278) );
AND2x2_ASAP7_75t_L g298 ( .A(n_167), .B(n_299), .Y(n_298) );
NOR2xp67_ASAP7_75t_L g423 ( .A(n_167), .B(n_299), .Y(n_423) );
AND2x2_ASAP7_75t_L g448 ( .A(n_167), .B(n_291), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_174), .B(n_203), .Y(n_215) );
INVx1_ASAP7_75t_L g232 ( .A(n_174), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_174), .A2(n_254), .B(n_255), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_174), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_174), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_174), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_174), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_174), .A2(n_545), .B(n_546), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_174), .A2(n_554), .B(n_555), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_174), .A2(n_578), .B(n_579), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_174), .A2(n_586), .B(n_587), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_176), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_176), .A2(n_500), .B(n_502), .Y(n_499) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_176), .A2(n_523), .B(n_527), .Y(n_522) );
OA21x2_ASAP7_75t_L g593 ( .A1(n_176), .A2(n_523), .B(n_527), .Y(n_593) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g240 ( .A(n_180), .Y(n_240) );
INVx1_ASAP7_75t_L g262 ( .A(n_180), .Y(n_262) );
INVxp67_ASAP7_75t_L g301 ( .A(n_180), .Y(n_301) );
AND2x4_ASAP7_75t_L g341 ( .A(n_180), .B(n_342), .Y(n_341) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_180), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_180), .B(n_292), .Y(n_427) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_186), .Y(n_180) );
INVx2_ASAP7_75t_SL g229 ( .A(n_181), .Y(n_229) );
INVx1_ASAP7_75t_SL g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_199), .Y(n_188) );
AND2x2_ASAP7_75t_L g315 ( .A(n_189), .B(n_287), .Y(n_315) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_190), .Y(n_243) );
AND2x2_ASAP7_75t_L g271 ( .A(n_190), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g282 ( .A(n_190), .Y(n_282) );
INVx1_ASAP7_75t_L g306 ( .A(n_190), .Y(n_306) );
AND2x2_ASAP7_75t_L g309 ( .A(n_190), .B(n_201), .Y(n_309) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_190), .Y(n_331) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_198), .Y(n_190) );
AO21x2_ASAP7_75t_L g582 ( .A1(n_191), .A2(n_583), .B(n_589), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
NOR2x1_ASAP7_75t_L g199 ( .A(n_200), .B(n_216), .Y(n_199) );
AND2x2_ASAP7_75t_L g296 ( .A(n_200), .B(n_218), .Y(n_296) );
NAND2x1_ASAP7_75t_L g329 ( .A(n_200), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g432 ( .A(n_200), .Y(n_432) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx3_ASAP7_75t_L g272 ( .A(n_201), .Y(n_272) );
AND2x2_ASAP7_75t_L g287 ( .A(n_201), .B(n_246), .Y(n_287) );
NOR2x1_ASAP7_75t_SL g356 ( .A(n_201), .B(n_218), .Y(n_356) );
AND2x4_ASAP7_75t_L g201 ( .A(n_202), .B(n_204), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_203), .A2(n_221), .B(n_225), .Y(n_220) );
INVx1_ASAP7_75t_SL g508 ( .A(n_203), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_203), .B(n_540), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_203), .A2(n_575), .B(n_576), .Y(n_574) );
OAI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_208), .B(n_215), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B1(n_212), .B2(n_213), .Y(n_208) );
INVxp67_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVxp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NOR2x1_ASAP7_75t_L g393 ( .A(n_216), .B(n_380), .Y(n_393) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g318 ( .A(n_217), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx4_ASAP7_75t_L g257 ( .A(n_218), .Y(n_257) );
AND2x4_ASAP7_75t_L g264 ( .A(n_218), .B(n_265), .Y(n_264) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_218), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_218), .B(n_281), .Y(n_381) );
AND2x2_ASAP7_75t_L g409 ( .A(n_218), .B(n_246), .Y(n_409) );
OR2x6_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
NAND2x1_ASAP7_75t_SL g226 ( .A(n_227), .B(n_239), .Y(n_226) );
OR2x2_ASAP7_75t_L g437 ( .A(n_227), .B(n_349), .Y(n_437) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x4_ASAP7_75t_L g277 ( .A(n_228), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g342 ( .A(n_228), .Y(n_342) );
AND2x2_ASAP7_75t_L g376 ( .A(n_228), .B(n_299), .Y(n_376) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_238), .Y(n_228) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_229), .A2(n_230), .B(n_238), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_231), .B(n_237), .Y(n_230) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx3_ASAP7_75t_L g349 ( .A(n_239), .Y(n_349) );
AND2x2_ASAP7_75t_L g357 ( .A(n_239), .B(n_290), .Y(n_357) );
AND2x2_ASAP7_75t_L g474 ( .A(n_239), .B(n_277), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g428 ( .A(n_243), .B(n_369), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_243), .B(n_268), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_244), .A2(n_305), .B(n_308), .Y(n_304) );
AND2x2_ASAP7_75t_L g374 ( .A(n_244), .B(n_280), .Y(n_374) );
INVx2_ASAP7_75t_SL g461 ( .A(n_244), .Y(n_461) );
AND2x4_ASAP7_75t_SL g244 ( .A(n_245), .B(n_257), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g265 ( .A(n_246), .Y(n_265) );
INVx2_ASAP7_75t_L g312 ( .A(n_246), .Y(n_312) );
AND2x4_ASAP7_75t_L g319 ( .A(n_246), .B(n_272), .Y(n_319) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_252), .Y(n_246) );
NOR3xp33_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .C(n_251), .Y(n_248) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_257), .Y(n_275) );
AND2x4_ASAP7_75t_L g351 ( .A(n_257), .B(n_265), .Y(n_351) );
OR2x2_ASAP7_75t_L g477 ( .A(n_257), .B(n_478), .Y(n_477) );
NAND4xp25_ASAP7_75t_L g258 ( .A(n_259), .B(n_263), .C(n_266), .D(n_271), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g324 ( .A(n_260), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g421 ( .A(n_260), .Y(n_421) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2x1p5_ASAP7_75t_L g321 ( .A(n_261), .B(n_269), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_261), .B(n_326), .Y(n_455) );
BUFx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_264), .B(n_280), .Y(n_333) );
INVx2_ASAP7_75t_L g435 ( .A(n_264), .Y(n_435) );
AND2x2_ASAP7_75t_SL g445 ( .A(n_264), .B(n_305), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_264), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g337 ( .A(n_268), .B(n_284), .Y(n_337) );
AND2x2_ASAP7_75t_L g405 ( .A(n_268), .B(n_341), .Y(n_405) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g290 ( .A(n_269), .B(n_291), .Y(n_290) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_270), .Y(n_344) );
AND2x2_ASAP7_75t_L g395 ( .A(n_270), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_270), .B(n_292), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_271), .B(n_435), .Y(n_442) );
INVx1_ASAP7_75t_SL g478 ( .A(n_271), .Y(n_478) );
INVx1_ASAP7_75t_L g307 ( .A(n_272), .Y(n_307) );
AND2x2_ASAP7_75t_L g369 ( .A(n_272), .B(n_312), .Y(n_369) );
OAI21xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_283), .B(n_285), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
AND2x2_ASAP7_75t_L g335 ( .A(n_277), .B(n_284), .Y(n_335) );
AND2x2_ASAP7_75t_L g443 ( .A(n_277), .B(n_294), .Y(n_443) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g317 ( .A(n_280), .Y(n_317) );
AND2x2_ASAP7_75t_L g350 ( .A(n_280), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g355 ( .A(n_280), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_280), .B(n_319), .Y(n_404) );
NOR3xp33_ASAP7_75t_L g454 ( .A(n_280), .B(n_455), .C(n_456), .Y(n_454) );
INVx3_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVxp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_289), .B1(n_296), .B2(n_297), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx2_ASAP7_75t_L g380 ( .A(n_287), .Y(n_380) );
AND2x2_ASAP7_75t_L g314 ( .A(n_288), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g336 ( .A(n_288), .B(n_309), .Y(n_336) );
AND2x2_ASAP7_75t_SL g368 ( .A(n_288), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
INVx1_ASAP7_75t_L g347 ( .A(n_290), .Y(n_347) );
AND2x2_ASAP7_75t_L g300 ( .A(n_291), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g326 ( .A(n_291), .Y(n_326) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g389 ( .A(n_295), .B(n_341), .Y(n_389) );
INVx1_ASAP7_75t_L g447 ( .A(n_295), .Y(n_447) );
INVx1_ASAP7_75t_L g303 ( .A(n_297), .Y(n_303) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
NAND2x1p5_ASAP7_75t_L g325 ( .A(n_298), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g434 ( .A(n_298), .B(n_341), .Y(n_434) );
AND2x2_ASAP7_75t_L g400 ( .A(n_300), .B(n_401), .Y(n_400) );
NAND2x1p5_ASAP7_75t_L g468 ( .A(n_300), .B(n_469), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B(n_313), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_305), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g361 ( .A(n_305), .B(n_310), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_305), .B(n_351), .Y(n_412) );
AND2x4_ASAP7_75t_SL g305 ( .A(n_306), .B(n_307), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_306), .B(n_369), .Y(n_399) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_306), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_308), .A2(n_335), .B1(n_336), .B2(n_337), .Y(n_334) );
AND2x2_ASAP7_75t_SL g308 ( .A(n_309), .B(n_310), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_309), .B(n_351), .Y(n_370) );
INVx1_ASAP7_75t_L g471 ( .A(n_309), .Y(n_471) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OAI21xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_316), .B(n_320), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_315), .B(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g452 ( .A(n_318), .Y(n_452) );
INVx4_ASAP7_75t_L g354 ( .A(n_319), .Y(n_354) );
INVxp33_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g382 ( .A(n_321), .B(n_383), .Y(n_382) );
NOR2x1_ASAP7_75t_L g322 ( .A(n_323), .B(n_338), .Y(n_322) );
OAI21xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_327), .B(n_334), .Y(n_323) );
INVx1_ASAP7_75t_L g372 ( .A(n_325), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_332), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g377 ( .A(n_329), .Y(n_377) );
INVx1_ASAP7_75t_L g410 ( .A(n_330), .Y(n_410) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_335), .A2(n_374), .B1(n_375), .B2(n_377), .Y(n_373) );
INVx1_ASAP7_75t_L g387 ( .A(n_336), .Y(n_387) );
NAND4xp25_ASAP7_75t_SL g338 ( .A(n_339), .B(n_345), .C(n_352), .D(n_358), .Y(n_338) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
INVx1_ASAP7_75t_L g360 ( .A(n_341), .Y(n_360) );
AND2x2_ASAP7_75t_L g472 ( .A(n_341), .B(n_469), .Y(n_472) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_350), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g479 ( .A(n_349), .B(n_416), .Y(n_479) );
INVx1_ASAP7_75t_L g476 ( .A(n_350), .Y(n_476) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_351), .Y(n_385) );
OAI21xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_355), .B(n_357), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_390), .Y(n_362) );
NOR3xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_378), .C(n_386), .Y(n_363) );
OAI21xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_371), .B(n_373), .Y(n_364) );
INVxp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_370), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_368), .A2(n_400), .B1(n_403), .B2(n_405), .Y(n_402) );
OAI22xp33_ASAP7_75t_L g378 ( .A1(n_371), .A2(n_379), .B1(n_382), .B2(n_384), .Y(n_378) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g383 ( .A(n_376), .Y(n_383) );
AND2x4_ASAP7_75t_L g394 ( .A(n_376), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_381), .Y(n_481) );
AOI31xp33_ASAP7_75t_L g480 ( .A1(n_384), .A2(n_457), .A3(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_406), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_392), .B(n_402), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B1(n_397), .B2(n_400), .Y(n_392) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_396), .Y(n_460) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_404), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_407), .B(n_417), .Y(n_406) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
AND2x2_ASAP7_75t_L g418 ( .A(n_409), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g457 ( .A(n_409), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g466 ( .A1(n_409), .A2(n_467), .B1(n_470), .B2(n_472), .Y(n_466) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_414), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_420), .B1(n_424), .B2(n_428), .Y(n_417) );
NOR2xp33_ASAP7_75t_SL g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVxp67_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx2_ASAP7_75t_SL g469 ( .A(n_426), .Y(n_469) );
INVx2_ASAP7_75t_L g450 ( .A(n_427), .Y(n_450) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_464), .Y(n_429) );
AOI211xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_436), .B(n_439), .C(n_453), .Y(n_430) );
OAI21xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B(n_435), .Y(n_431) );
INVx1_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g438 ( .A(n_435), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_440), .B(n_444), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_443), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_449), .B2(n_451), .Y(n_444) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
AND2x2_ASAP7_75t_L g449 ( .A(n_447), .B(n_450), .Y(n_449) );
AO22x1_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_457), .B1(n_458), .B2(n_462), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_475), .C(n_480), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_466), .B(n_473), .Y(n_465) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AOI21xp33_ASAP7_75t_R g475 ( .A1(n_476), .A2(n_477), .B(n_479), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_484), .Y(n_791) );
CKINVDCx11_ASAP7_75t_R g484 ( .A(n_485), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx3_ASAP7_75t_SL g792 ( .A(n_491), .Y(n_792) );
NOR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_672), .Y(n_491) );
AO211x2_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_517), .B(n_567), .C(n_640), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVxp67_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
AND3x2_ASAP7_75t_L g721 ( .A(n_495), .B(n_602), .C(n_618), .Y(n_721) );
AND2x4_ASAP7_75t_L g724 ( .A(n_495), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_507), .Y(n_495) );
NAND2x1p5_ASAP7_75t_L g580 ( .A(n_496), .B(n_581), .Y(n_580) );
INVx4_ASAP7_75t_L g633 ( .A(n_496), .Y(n_633) );
AND2x2_ASAP7_75t_SL g718 ( .A(n_496), .B(n_627), .Y(n_718) );
AND2x2_ASAP7_75t_L g761 ( .A(n_496), .B(n_582), .Y(n_761) );
INVx5_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g610 ( .A(n_497), .Y(n_610) );
AND2x2_ASAP7_75t_L g629 ( .A(n_497), .B(n_573), .Y(n_629) );
AND2x2_ASAP7_75t_L g647 ( .A(n_497), .B(n_582), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_497), .B(n_581), .Y(n_707) );
NOR2x1_ASAP7_75t_SL g734 ( .A(n_497), .B(n_507), .Y(n_734) );
OR2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_507), .B(n_573), .Y(n_572) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B(n_515), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_508), .B(n_516), .Y(n_515) );
AO21x2_ASAP7_75t_L g606 ( .A1(n_508), .A2(n_509), .B(n_515), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_514), .Y(n_509) );
AO21x1_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_549), .B(n_558), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_519), .A2(n_616), .B1(n_620), .B2(n_621), .Y(n_615) );
OR2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_528), .Y(n_519) );
AND2x2_ASAP7_75t_L g676 ( .A(n_520), .B(n_564), .Y(n_676) );
BUFx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x4_ASAP7_75t_L g609 ( .A(n_521), .B(n_592), .Y(n_609) );
AND2x2_ASAP7_75t_L g681 ( .A(n_521), .B(n_566), .Y(n_681) );
AND2x2_ASAP7_75t_L g700 ( .A(n_521), .B(n_666), .Y(n_700) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g559 ( .A(n_522), .Y(n_559) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_522), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_528), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g660 ( .A(n_529), .B(n_561), .Y(n_660) );
AND2x4_ASAP7_75t_L g529 ( .A(n_530), .B(n_541), .Y(n_529) );
AND2x2_ASAP7_75t_L g564 ( .A(n_530), .B(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g597 ( .A(n_530), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_SL g657 ( .A(n_530), .B(n_593), .Y(n_657) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g750 ( .A(n_531), .Y(n_750) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g592 ( .A(n_532), .Y(n_592) );
OAI21x1_ASAP7_75t_SL g532 ( .A1(n_533), .A2(n_535), .B(n_539), .Y(n_532) );
INVx1_ASAP7_75t_L g540 ( .A(n_534), .Y(n_540) );
INVx2_ASAP7_75t_L g598 ( .A(n_541), .Y(n_598) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_541), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_543), .B(n_547), .Y(n_542) );
INVx2_ASAP7_75t_L g594 ( .A(n_549), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_549), .B(n_726), .Y(n_752) );
AND2x2_ASAP7_75t_L g771 ( .A(n_549), .B(n_761), .Y(n_771) );
BUFx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x4_ASAP7_75t_SL g639 ( .A(n_550), .B(n_598), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_556), .Y(n_551) );
AND2x2_ASAP7_75t_SL g558 ( .A(n_559), .B(n_560), .Y(n_558) );
AND2x2_ASAP7_75t_L g638 ( .A(n_559), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_559), .B(n_608), .Y(n_643) );
INVx1_ASAP7_75t_SL g770 ( .A(n_559), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_560), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_564), .Y(n_560) );
INVx1_ASAP7_75t_L g596 ( .A(n_561), .Y(n_596) );
AND2x2_ASAP7_75t_L g782 ( .A(n_561), .B(n_783), .Y(n_782) );
BUFx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g658 ( .A(n_562), .B(n_565), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_562), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g712 ( .A(n_562), .B(n_566), .Y(n_712) );
AND2x2_ASAP7_75t_L g743 ( .A(n_562), .B(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g608 ( .A(n_563), .B(n_566), .Y(n_608) );
INVxp67_ASAP7_75t_L g625 ( .A(n_563), .Y(n_625) );
BUFx3_ASAP7_75t_L g666 ( .A(n_563), .Y(n_666) );
AND2x2_ASAP7_75t_L g686 ( .A(n_564), .B(n_687), .Y(n_686) );
NAND2xp33_ASAP7_75t_L g699 ( .A(n_564), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_565), .B(n_592), .Y(n_655) );
AND2x2_ASAP7_75t_L g744 ( .A(n_565), .B(n_593), .Y(n_744) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g671 ( .A(n_566), .B(n_593), .Y(n_671) );
OR3x1_ASAP7_75t_L g567 ( .A(n_568), .B(n_615), .C(n_630), .Y(n_567) );
OAI321xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_580), .A3(n_590), .B1(n_595), .B2(n_599), .C(n_607), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVxp67_ASAP7_75t_SL g646 ( .A(n_572), .Y(n_646) );
INVxp67_ASAP7_75t_SL g664 ( .A(n_572), .Y(n_664) );
OR2x2_ASAP7_75t_L g668 ( .A(n_572), .B(n_580), .Y(n_668) );
BUFx3_ASAP7_75t_L g602 ( .A(n_573), .Y(n_602) );
AND2x2_ASAP7_75t_L g619 ( .A(n_573), .B(n_605), .Y(n_619) );
INVx1_ASAP7_75t_L g636 ( .A(n_573), .Y(n_636) );
INVx2_ASAP7_75t_L g652 ( .A(n_573), .Y(n_652) );
OR2x2_ASAP7_75t_L g691 ( .A(n_573), .B(n_581), .Y(n_691) );
INVx2_ASAP7_75t_L g679 ( .A(n_580), .Y(n_679) );
AND2x2_ASAP7_75t_L g603 ( .A(n_581), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g618 ( .A(n_581), .Y(n_618) );
AND2x4_ASAP7_75t_L g627 ( .A(n_581), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_581), .B(n_604), .Y(n_650) );
AND2x2_ASAP7_75t_L g757 ( .A(n_581), .B(n_652), .Y(n_757) );
INVx4_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_582), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_588), .Y(n_583) );
INVx1_ASAP7_75t_L g644 ( .A(n_590), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_591), .B(n_594), .Y(n_590) );
AND2x2_ASAP7_75t_L g731 ( .A(n_591), .B(n_658), .Y(n_731) );
INVx1_ASAP7_75t_SL g748 ( .A(n_591), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_591), .B(n_724), .Y(n_777) );
AND2x4_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
OR2x2_ASAP7_75t_L g620 ( .A(n_592), .B(n_593), .Y(n_620) );
AND2x2_ASAP7_75t_L g713 ( .A(n_594), .B(n_609), .Y(n_713) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g736 ( .A(n_598), .B(n_609), .Y(n_736) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_600), .A2(n_749), .B1(n_754), .B2(n_756), .Y(n_753) );
AND2x4_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
AND2x2_ASAP7_75t_L g678 ( .A(n_601), .B(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g773 ( .A(n_601), .B(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g729 ( .A(n_602), .B(n_647), .Y(n_729) );
AND2x4_ASAP7_75t_L g683 ( .A(n_603), .B(n_629), .Y(n_683) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_605), .Y(n_781) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g614 ( .A(n_606), .Y(n_614) );
INVx1_ASAP7_75t_L g628 ( .A(n_606), .Y(n_628) );
NAND4xp25_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .C(n_610), .D(n_611), .Y(n_607) );
AND2x2_ASAP7_75t_L g765 ( .A(n_608), .B(n_750), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_608), .B(n_776), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_609), .B(n_685), .Y(n_684) );
OAI322xp33_ASAP7_75t_L g692 ( .A1(n_609), .A2(n_693), .A3(n_697), .B1(n_699), .B2(n_701), .C1(n_703), .C2(n_708), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_609), .B(n_658), .Y(n_708) );
INVx1_ASAP7_75t_L g776 ( .A(n_609), .Y(n_776) );
INVx2_ASAP7_75t_L g622 ( .A(n_610), .Y(n_622) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_613), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_614), .B(n_633), .Y(n_690) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_617), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g663 ( .A(n_618), .Y(n_663) );
AND2x2_ASAP7_75t_L g735 ( .A(n_618), .B(n_646), .Y(n_735) );
AOI31xp33_ASAP7_75t_L g621 ( .A1(n_619), .A2(n_622), .A3(n_623), .B(n_626), .Y(n_621) );
AND2x2_ASAP7_75t_L g632 ( .A(n_619), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g760 ( .A(n_619), .B(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_SL g767 ( .A(n_619), .B(n_647), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_619), .Y(n_768) );
INVx1_ASAP7_75t_SL g726 ( .A(n_620), .Y(n_726) );
NAND3xp33_ASAP7_75t_SL g754 ( .A(n_620), .B(n_748), .C(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g654 ( .A(n_625), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
AND2x2_ASAP7_75t_L g635 ( .A(n_627), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g696 ( .A(n_627), .Y(n_696) );
AOI322xp5_ASAP7_75t_L g778 ( .A1(n_627), .A2(n_657), .A3(n_660), .B1(n_779), .B2(n_780), .C1(n_782), .C2(n_784), .Y(n_778) );
AND2x2_ASAP7_75t_L g784 ( .A(n_627), .B(n_633), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_634), .B(n_637), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_633), .B(n_652), .Y(n_651) );
AND2x4_ASAP7_75t_L g779 ( .A(n_633), .B(n_666), .Y(n_779) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g705 ( .A(n_636), .Y(n_705) );
AND2x2_ASAP7_75t_L g733 ( .A(n_636), .B(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g780 ( .A(n_636), .B(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g685 ( .A(n_639), .Y(n_685) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
O2A1O1Ixp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_644), .B(n_645), .C(n_648), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
AND2x2_ASAP7_75t_L g702 ( .A(n_647), .B(n_652), .Y(n_702) );
OAI211xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_653), .B(n_659), .C(n_661), .Y(n_648) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_649), .A2(n_675), .B1(n_677), .B2(n_680), .C(n_682), .Y(n_674) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g694 ( .A(n_651), .Y(n_694) );
OR2x2_ASAP7_75t_L g714 ( .A(n_651), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .Y(n_653) );
INVx1_ASAP7_75t_L g759 ( .A(n_654), .Y(n_759) );
INVx1_ASAP7_75t_L g783 ( .A(n_655), .Y(n_783) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_657), .B(n_658), .Y(n_656) );
AND2x2_ASAP7_75t_L g665 ( .A(n_657), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_657), .B(n_727), .Y(n_739) );
INVx1_ASAP7_75t_L g719 ( .A(n_658), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_665), .B1(n_667), .B2(n_669), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_SL g727 ( .A(n_666), .Y(n_727) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND4xp75_ASAP7_75t_L g672 ( .A(n_673), .B(n_709), .C(n_737), .D(n_762), .Y(n_672) );
NOR2xp67_ASAP7_75t_L g673 ( .A(n_674), .B(n_692), .Y(n_673) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_SL g749 ( .A(n_681), .B(n_750), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B1(n_686), .B2(n_688), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_685), .B(n_748), .Y(n_747) );
INVx2_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
INVx2_ASAP7_75t_L g725 ( .A(n_691), .Y(n_725) );
OR2x2_ASAP7_75t_L g740 ( .A(n_691), .B(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g755 ( .A(n_700), .Y(n_755) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
OAI21xp5_ASAP7_75t_SL g746 ( .A1(n_702), .A2(n_747), .B(n_749), .Y(n_746) );
INVxp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NOR2x1_ASAP7_75t_L g709 ( .A(n_710), .B(n_722), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_714), .B1(n_717), .B2(n_719), .C(n_720), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
OAI21xp33_ASAP7_75t_L g758 ( .A1(n_712), .A2(n_759), .B(n_760), .Y(n_758) );
INVx3_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
OAI322xp33_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_726), .A3(n_727), .B1(n_728), .B2(n_730), .C1(n_732), .C2(n_736), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
NOR2x1_ASAP7_75t_L g732 ( .A(n_733), .B(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g745 ( .A(n_733), .Y(n_745) );
INVx1_ASAP7_75t_L g741 ( .A(n_734), .Y(n_741) );
AND2x2_ASAP7_75t_L g756 ( .A(n_734), .B(n_757), .Y(n_756) );
NOR2x1_ASAP7_75t_L g737 ( .A(n_738), .B(n_751), .Y(n_737) );
OAI221xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .B1(n_742), .B2(n_745), .C(n_746), .Y(n_738) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
OAI211xp5_ASAP7_75t_SL g751 ( .A1(n_745), .A2(n_752), .B(n_753), .C(n_758), .Y(n_751) );
INVx2_ASAP7_75t_SL g774 ( .A(n_761), .Y(n_774) );
NOR2x1_ASAP7_75t_L g762 ( .A(n_763), .B(n_772), .Y(n_762) );
OAI22xp33_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_766), .B1(n_768), .B2(n_769), .Y(n_763) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
OAI211xp5_ASAP7_75t_SL g772 ( .A1(n_773), .A2(n_775), .B(n_777), .C(n_778), .Y(n_772) );
CKINVDCx11_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
INVx3_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
CKINVDCx11_ASAP7_75t_R g793 ( .A(n_788), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
INVx3_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g807 ( .A1(n_799), .A2(n_808), .B(n_811), .Y(n_807) );
CKINVDCx14_ASAP7_75t_R g799 ( .A(n_800), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_802), .B(n_809), .Y(n_808) );
BUFx3_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_806), .Y(n_813) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_813), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
endmodule