module fake_netlist_6_1312_n_1756 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1756);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1756;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_52),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_69),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_79),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_140),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_36),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_81),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_22),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_25),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_137),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_108),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_27),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_130),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_136),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_89),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_41),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_26),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_5),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_14),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_80),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_99),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_135),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_29),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_53),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_49),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_124),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_134),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_83),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_10),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_105),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_147),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_57),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_90),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_176),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_61),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_16),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_28),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_1),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_22),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_169),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_17),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_92),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_138),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_70),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_65),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_168),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_2),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_111),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_3),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_66),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_71),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_133),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_16),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_10),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_74),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_77),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_119),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_60),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_172),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_161),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_91),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_43),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_45),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_72),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_35),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_114),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_164),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_170),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_167),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_67),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_18),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_103),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_53),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_97),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_31),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_13),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_155),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_13),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_45),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_139),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_93),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_131),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_128),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_41),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_162),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_40),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_143),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_50),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_110),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_43),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_148),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_62),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_102),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_37),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_171),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_42),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_177),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_178),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_26),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_18),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_100),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_23),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_84),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_29),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_113),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_68),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_14),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_52),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_34),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_123),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_175),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_5),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_49),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_33),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_106),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_87),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_42),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_4),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_55),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_1),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_21),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_126),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_116),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_158),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_44),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_27),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_141),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_144),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_48),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_21),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_58),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_34),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_39),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_11),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_0),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_150),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_104),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_24),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_156),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_3),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_31),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_149),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_28),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_142),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_39),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_101),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_24),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_12),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_120),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_78),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_85),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_95),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_117),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_73),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_12),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_154),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_96),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_51),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_118),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_82),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_23),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_64),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_165),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_54),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_88),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_59),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_32),
.Y(n_351)
);

BUFx10_ASAP7_75t_L g352 ( 
.A(n_19),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_7),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_151),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_115),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_76),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_180),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_180),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_269),
.B(n_0),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_193),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_213),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_221),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_222),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_194),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_188),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_188),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_188),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_188),
.Y(n_368)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_280),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_205),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_223),
.Y(n_371)
);

BUFx6f_ASAP7_75t_SL g372 ( 
.A(n_182),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_217),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_196),
.B(n_2),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_225),
.Y(n_375)
);

INVxp33_ASAP7_75t_SL g376 ( 
.A(n_187),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_191),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_231),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_276),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_233),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_238),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_247),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_249),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_263),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_320),
.B(n_245),
.Y(n_385)
);

NAND2xp33_ASAP7_75t_R g386 ( 
.A(n_179),
.B(n_4),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_188),
.Y(n_387)
);

BUFx6f_ASAP7_75t_SL g388 ( 
.A(n_182),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_320),
.B(n_6),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_276),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_199),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_270),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_187),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_199),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_272),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_274),
.Y(n_396)
);

BUFx2_ASAP7_75t_SL g397 ( 
.A(n_230),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_199),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_288),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_350),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_234),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_347),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_191),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_212),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_292),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_191),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_293),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_199),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_198),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_199),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_214),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_218),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_301),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_335),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_219),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_198),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_224),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_227),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_284),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_257),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_228),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_324),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_257),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_229),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_325),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_201),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_257),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_327),
.Y(n_428)
);

INVxp33_ASAP7_75t_SL g429 ( 
.A(n_201),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_329),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_332),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_339),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_232),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_342),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_257),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_257),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_314),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_R g438 ( 
.A(n_236),
.B(n_174),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g439 ( 
.A(n_207),
.B(n_6),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_284),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_314),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_314),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_335),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_284),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_239),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_360),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_365),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_366),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_390),
.B(n_245),
.Y(n_449)
);

CKINVDCx6p67_ASAP7_75t_R g450 ( 
.A(n_372),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_374),
.B(n_248),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_196),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_367),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_404),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_368),
.Y(n_455)
);

CKINVDCx9p33_ASAP7_75t_R g456 ( 
.A(n_359),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_364),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_362),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_R g459 ( 
.A(n_411),
.B(n_240),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_373),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_412),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_415),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_387),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_406),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_391),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_362),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_394),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_400),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_398),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_408),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_417),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_410),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_374),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_420),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_423),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_427),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_435),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_436),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_376),
.B(n_429),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_379),
.B(n_248),
.Y(n_480)
);

AND3x2_ASAP7_75t_L g481 ( 
.A(n_385),
.B(n_278),
.C(n_255),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_418),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_437),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_441),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_442),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_421),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_424),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_379),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_357),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_414),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_414),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_433),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_358),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_445),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_397),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_361),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_363),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_389),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_363),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_371),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_393),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_371),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_439),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_370),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_375),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_402),
.B(n_261),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_375),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_409),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_378),
.B(n_261),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_378),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_380),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_416),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_426),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_380),
.Y(n_514)
);

BUFx8_ASAP7_75t_L g515 ( 
.A(n_372),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_377),
.B(n_271),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_381),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_438),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_381),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_382),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_382),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_383),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g523 ( 
.A(n_451),
.B(n_271),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_473),
.B(n_281),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_446),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_473),
.B(n_383),
.Y(n_526)
);

AND2x2_ASAP7_75t_SL g527 ( 
.A(n_519),
.B(n_281),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_447),
.Y(n_528)
);

BUFx4f_ASAP7_75t_L g529 ( 
.A(n_450),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_491),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_509),
.B(n_504),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_491),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_447),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_491),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_490),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_479),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_488),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_488),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_490),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_490),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_489),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_447),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_504),
.B(n_384),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_SL g544 ( 
.A1(n_506),
.A2(n_440),
.B1(n_444),
.B2(n_403),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_513),
.B(n_419),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_498),
.A2(n_237),
.B1(n_314),
.B2(n_338),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_522),
.A2(n_401),
.B1(n_432),
.B2(n_431),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_490),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_473),
.B(n_384),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_483),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_483),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_483),
.Y(n_552)
);

AO22x2_ASAP7_75t_L g553 ( 
.A1(n_498),
.A2(n_237),
.B1(n_338),
.B2(n_348),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_473),
.B(n_392),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_519),
.B(n_256),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_513),
.B(n_464),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_482),
.Y(n_557)
);

BUFx4f_ASAP7_75t_L g558 ( 
.A(n_450),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_519),
.B(n_256),
.Y(n_559)
);

OR2x6_ASAP7_75t_L g560 ( 
.A(n_519),
.B(n_283),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_490),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_484),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_L g563 ( 
.A(n_514),
.B(n_392),
.Y(n_563)
);

AND3x2_ASAP7_75t_L g564 ( 
.A(n_458),
.B(n_246),
.C(n_220),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_513),
.B(n_395),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_490),
.B(n_259),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_451),
.B(n_256),
.Y(n_567)
);

BUFx4f_ASAP7_75t_L g568 ( 
.A(n_519),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_485),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_485),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_493),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_485),
.Y(n_572)
);

AO21x2_ASAP7_75t_L g573 ( 
.A1(n_514),
.A2(n_200),
.B(n_186),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_519),
.B(n_256),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_514),
.B(n_256),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_508),
.B(n_395),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_484),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_484),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_496),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_508),
.B(n_396),
.Y(n_580)
);

INVxp67_ASAP7_75t_SL g581 ( 
.A(n_451),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_518),
.B(n_451),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_472),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_496),
.Y(n_584)
);

OAI21xp33_ASAP7_75t_SL g585 ( 
.A1(n_449),
.A2(n_262),
.B(n_260),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_522),
.A2(n_434),
.B1(n_432),
.B2(n_431),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_517),
.B(n_396),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_452),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_487),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_501),
.B(n_399),
.Y(n_590)
);

BUFx6f_ASAP7_75t_SL g591 ( 
.A(n_512),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_472),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_518),
.B(n_399),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_512),
.B(n_405),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_485),
.Y(n_595)
);

INVx4_ASAP7_75t_SL g596 ( 
.A(n_485),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_485),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_517),
.B(n_405),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_448),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_448),
.Y(n_600)
);

AND2x2_ASAP7_75t_SL g601 ( 
.A(n_458),
.B(n_466),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_453),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_464),
.B(n_407),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_452),
.B(n_286),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_453),
.Y(n_605)
);

OAI21xp33_ASAP7_75t_SL g606 ( 
.A1(n_503),
.A2(n_297),
.B(n_296),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_503),
.B(n_407),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_455),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_455),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_463),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_463),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_502),
.B(n_413),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_502),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_465),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_502),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_465),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_499),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_516),
.B(n_298),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_467),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_501),
.B(n_413),
.Y(n_620)
);

INVx5_ASAP7_75t_L g621 ( 
.A(n_516),
.Y(n_621)
);

NAND2xp33_ASAP7_75t_R g622 ( 
.A(n_466),
.B(n_422),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_501),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_502),
.B(n_422),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_480),
.B(n_467),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_469),
.B(n_425),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_469),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_L g628 ( 
.A(n_501),
.B(n_425),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_511),
.B(n_428),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_470),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_501),
.B(n_305),
.Y(n_631)
);

OAI22xp33_ASAP7_75t_L g632 ( 
.A1(n_501),
.A2(n_369),
.B1(n_309),
.B2(n_302),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_511),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_516),
.A2(n_314),
.B1(n_313),
.B2(n_310),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_470),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_511),
.B(n_428),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_474),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_474),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_475),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_511),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_475),
.B(n_430),
.Y(n_641)
);

INVxp67_ASAP7_75t_SL g642 ( 
.A(n_476),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_476),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_516),
.B(n_430),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_497),
.B(n_319),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_477),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_477),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_478),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_500),
.A2(n_434),
.B1(n_386),
.B2(n_388),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_478),
.Y(n_650)
);

NOR2x1p5_ASAP7_75t_L g651 ( 
.A(n_505),
.B(n_208),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_497),
.B(n_345),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_459),
.B(n_495),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_481),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_520),
.B(n_507),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_510),
.B(n_203),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_520),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_521),
.B(n_208),
.Y(n_658)
);

NAND3xp33_ASAP7_75t_L g659 ( 
.A(n_515),
.B(n_302),
.C(n_209),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_L g660 ( 
.A(n_456),
.B(n_179),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_515),
.Y(n_661)
);

AND2x6_ASAP7_75t_L g662 ( 
.A(n_515),
.B(n_210),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_515),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_454),
.Y(n_664)
);

AND2x6_ASAP7_75t_L g665 ( 
.A(n_461),
.B(n_211),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_462),
.A2(n_311),
.B1(n_215),
.B2(n_216),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_471),
.B(n_352),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_457),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_486),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_460),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_492),
.B(n_226),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_531),
.B(n_185),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_SL g673 ( 
.A(n_666),
.B(n_291),
.C(n_331),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_527),
.B(n_258),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_581),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_581),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_531),
.B(n_235),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_527),
.A2(n_287),
.B1(n_356),
.B2(n_307),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_528),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_612),
.B(n_494),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_565),
.B(n_352),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_541),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_576),
.B(n_209),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_525),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_582),
.B(n_241),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_568),
.B(n_333),
.Y(n_686)
);

NOR2xp67_ASAP7_75t_L g687 ( 
.A(n_661),
.B(n_242),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_640),
.B(n_243),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_593),
.B(n_181),
.Y(n_689)
);

NAND2x1_ASAP7_75t_L g690 ( 
.A(n_523),
.B(n_254),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_670),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_670),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_546),
.A2(n_268),
.B1(n_351),
.B2(n_317),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_566),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_613),
.B(n_295),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_657),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_613),
.B(n_615),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_528),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_615),
.B(n_306),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_543),
.B(n_181),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_633),
.B(n_330),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_568),
.B(n_336),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_543),
.B(n_183),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_633),
.B(n_341),
.Y(n_704)
);

O2A1O1Ixp5_ASAP7_75t_L g705 ( 
.A1(n_524),
.A2(n_349),
.B(n_388),
.C(n_372),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_546),
.A2(n_184),
.B1(n_318),
.B2(n_322),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_607),
.B(n_526),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_642),
.B(n_244),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_566),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_642),
.B(n_250),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_625),
.B(n_251),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_533),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_554),
.A2(n_629),
.B1(n_612),
.B2(n_644),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_588),
.B(n_252),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_537),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_553),
.A2(n_353),
.B1(n_318),
.B2(n_304),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_588),
.B(n_253),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_548),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_533),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_549),
.B(n_183),
.Y(n_720)
);

AOI221xp5_ASAP7_75t_L g721 ( 
.A1(n_632),
.A2(n_304),
.B1(n_309),
.B2(n_316),
.C(n_353),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_602),
.B(n_264),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_553),
.A2(n_316),
.B1(n_322),
.B2(n_352),
.Y(n_723)
);

INVx8_ASAP7_75t_L g724 ( 
.A(n_665),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_657),
.B(n_468),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_538),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_602),
.B(n_265),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_530),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_614),
.B(n_266),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_614),
.B(n_267),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_623),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_616),
.B(n_273),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_524),
.A2(n_299),
.B(n_275),
.Y(n_733)
);

NAND3xp33_ASAP7_75t_L g734 ( 
.A(n_666),
.B(n_303),
.C(n_355),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_621),
.B(n_277),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_580),
.B(n_189),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_616),
.B(n_279),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_545),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_532),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_553),
.A2(n_182),
.B1(n_388),
.B2(n_354),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_539),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_554),
.B(n_282),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_617),
.Y(n_743)
);

O2A1O1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_606),
.A2(n_285),
.B(n_289),
.C(n_290),
.Y(n_744)
);

AND2x6_ASAP7_75t_SL g745 ( 
.A(n_664),
.B(n_7),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_621),
.B(n_294),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_621),
.B(n_300),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_587),
.B(n_189),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_534),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_634),
.A2(n_355),
.B1(n_354),
.B2(n_346),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_617),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_629),
.B(n_346),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_621),
.B(n_323),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_573),
.B(n_326),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_573),
.B(n_328),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_644),
.A2(n_334),
.B(n_343),
.C(n_340),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_634),
.A2(n_344),
.B1(n_190),
.B2(n_321),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_587),
.B(n_344),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_624),
.B(n_206),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_571),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_598),
.B(n_206),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_556),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_542),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_550),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_618),
.B(n_204),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_539),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_599),
.B(n_337),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_579),
.Y(n_768)
);

OAI221xp5_ASAP7_75t_L g769 ( 
.A1(n_585),
.A2(n_321),
.B1(n_315),
.B2(n_312),
.C(n_308),
.Y(n_769)
);

BUFx4f_ASAP7_75t_L g770 ( 
.A(n_665),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_598),
.B(n_202),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_584),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_608),
.Y(n_773)
);

OAI221xp5_ASAP7_75t_L g774 ( 
.A1(n_626),
.A2(n_315),
.B1(n_312),
.B2(n_308),
.C(n_303),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_658),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_655),
.B(n_204),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_609),
.B(n_202),
.Y(n_777)
);

INVx4_ASAP7_75t_L g778 ( 
.A(n_539),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_539),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_600),
.B(n_195),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_604),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_619),
.Y(n_782)
);

NOR2xp67_ASAP7_75t_L g783 ( 
.A(n_661),
.B(n_197),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_627),
.B(n_197),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_630),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_550),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_641),
.B(n_195),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_551),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_551),
.Y(n_789)
);

NAND3xp33_ASAP7_75t_L g790 ( 
.A(n_563),
.B(n_192),
.C(n_190),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_637),
.B(n_192),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_594),
.B(n_652),
.Y(n_792)
);

NAND3xp33_ASAP7_75t_L g793 ( 
.A(n_586),
.B(n_8),
.C(n_9),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_646),
.B(n_160),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_600),
.B(n_159),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_600),
.B(n_635),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_600),
.B(n_145),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_635),
.B(n_132),
.Y(n_798)
);

AND2x6_ASAP7_75t_SL g799 ( 
.A(n_669),
.B(n_8),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_635),
.B(n_129),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_635),
.B(n_127),
.Y(n_801)
);

NAND3xp33_ASAP7_75t_L g802 ( 
.A(n_660),
.B(n_9),
.C(n_11),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_L g803 ( 
.A(n_523),
.B(n_125),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_548),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_622),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_636),
.A2(n_122),
.B1(n_121),
.B2(n_112),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_560),
.B(n_15),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_647),
.B(n_109),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_605),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_636),
.B(n_15),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_647),
.B(n_107),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_656),
.B(n_17),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_656),
.B(n_19),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_665),
.A2(n_628),
.B1(n_590),
.B2(n_620),
.Y(n_814)
);

AO22x1_ASAP7_75t_L g815 ( 
.A1(n_654),
.A2(n_20),
.B1(n_25),
.B2(n_30),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_604),
.A2(n_20),
.B(n_30),
.C(n_32),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_560),
.B(n_33),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_647),
.B(n_98),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_618),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_647),
.B(n_94),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_560),
.A2(n_86),
.B1(n_75),
.B2(n_63),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_649),
.B(n_632),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_547),
.B(n_38),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_665),
.A2(n_56),
.B1(n_40),
.B2(n_44),
.Y(n_824)
);

BUFx6f_ASAP7_75t_SL g825 ( 
.A(n_601),
.Y(n_825)
);

INVx8_ASAP7_75t_L g826 ( 
.A(n_665),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_523),
.B(n_54),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_523),
.B(n_38),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_552),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_523),
.B(n_51),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_631),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_552),
.Y(n_832)
);

A2O1A1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_605),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_555),
.B(n_46),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_645),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_590),
.A2(n_47),
.B1(n_50),
.B2(n_620),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_555),
.B(n_574),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_631),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_697),
.A2(n_574),
.B(n_559),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_672),
.B(n_650),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_672),
.A2(n_700),
.B(n_703),
.C(n_707),
.Y(n_841)
);

AOI21x1_ASAP7_75t_L g842 ( 
.A1(n_695),
.A2(n_559),
.B(n_575),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_679),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_796),
.A2(n_535),
.B(n_540),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_713),
.A2(n_601),
.B1(n_575),
.B2(n_645),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_707),
.B(n_648),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_805),
.B(n_536),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_675),
.B(n_648),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_698),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_712),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_718),
.A2(n_535),
.B(n_540),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_718),
.A2(n_572),
.B(n_597),
.Y(n_852)
);

AOI21x1_ASAP7_75t_L g853 ( 
.A1(n_699),
.A2(n_595),
.B(n_583),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_701),
.A2(n_572),
.B(n_597),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_676),
.B(n_611),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_704),
.A2(n_570),
.B(n_569),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_700),
.B(n_536),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_677),
.B(n_611),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_684),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_703),
.A2(n_650),
.B(n_610),
.C(n_643),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_748),
.B(n_610),
.Y(n_861)
);

AOI21x1_ASAP7_75t_L g862 ( 
.A1(n_837),
.A2(n_595),
.B(n_583),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_748),
.B(n_668),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_696),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_691),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_758),
.B(n_638),
.Y(n_866)
);

A2O1A1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_810),
.A2(n_639),
.B(n_671),
.C(n_529),
.Y(n_867)
);

A2O1A1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_810),
.A2(n_671),
.B(n_529),
.C(n_558),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_719),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_778),
.A2(n_570),
.B(n_569),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_743),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_792),
.B(n_667),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_758),
.B(n_592),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_725),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_837),
.A2(n_561),
.B(n_578),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_761),
.B(n_577),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_812),
.A2(n_631),
.B1(n_567),
.B2(n_645),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_835),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_761),
.B(n_562),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_792),
.B(n_603),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_762),
.B(n_653),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_674),
.A2(n_561),
.B(n_578),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_682),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_674),
.A2(n_577),
.B(n_562),
.Y(n_884)
);

NOR2xp67_ASAP7_75t_L g885 ( 
.A(n_814),
.B(n_653),
.Y(n_885)
);

AOI21x1_ASAP7_75t_L g886 ( 
.A1(n_685),
.A2(n_702),
.B(n_754),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_778),
.A2(n_567),
.B(n_596),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_803),
.A2(n_567),
.B(n_596),
.Y(n_888)
);

NAND3xp33_ASAP7_75t_L g889 ( 
.A(n_693),
.B(n_813),
.C(n_812),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_720),
.A2(n_622),
.B1(n_651),
.B2(n_567),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_720),
.B(n_567),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_741),
.A2(n_596),
.B(n_544),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_741),
.A2(n_558),
.B(n_659),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_741),
.A2(n_663),
.B(n_589),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_741),
.A2(n_557),
.B(n_662),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_766),
.A2(n_662),
.B(n_564),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_775),
.B(n_591),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_755),
.A2(n_756),
.B(n_702),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_787),
.B(n_591),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_781),
.B(n_564),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_766),
.A2(n_662),
.B(n_779),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_766),
.A2(n_662),
.B(n_779),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_766),
.A2(n_662),
.B(n_779),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_773),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_689),
.B(n_787),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_681),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_782),
.Y(n_907)
);

OAI21x1_ASAP7_75t_L g908 ( 
.A1(n_763),
.A2(n_829),
.B(n_764),
.Y(n_908)
);

NAND2x1p5_ASAP7_75t_L g909 ( 
.A(n_770),
.B(n_694),
.Y(n_909)
);

AOI21x1_ASAP7_75t_L g910 ( 
.A1(n_688),
.A2(n_722),
.B(n_727),
.Y(n_910)
);

AOI21x1_ASAP7_75t_L g911 ( 
.A1(n_729),
.A2(n_737),
.B(n_730),
.Y(n_911)
);

NOR2xp67_ASAP7_75t_L g912 ( 
.A(n_790),
.B(n_738),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_779),
.A2(n_732),
.B(n_714),
.Y(n_913)
);

AOI21x1_ASAP7_75t_L g914 ( 
.A1(n_728),
.A2(n_739),
.B(n_749),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_776),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_717),
.A2(n_746),
.B(n_753),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_770),
.A2(n_709),
.B1(n_742),
.B2(n_822),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_813),
.A2(n_678),
.B(n_686),
.C(n_771),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_689),
.B(n_785),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_747),
.A2(n_686),
.B(n_711),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_797),
.A2(n_801),
.B(n_800),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_831),
.B(n_838),
.Y(n_922)
);

O2A1O1Ixp33_ASAP7_75t_SL g923 ( 
.A1(n_834),
.A2(n_808),
.B(n_798),
.C(n_795),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_811),
.A2(n_820),
.B(n_818),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_708),
.A2(n_710),
.B(n_767),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_786),
.B(n_788),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_680),
.B(n_771),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_765),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_789),
.B(n_832),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_836),
.A2(n_744),
.B(n_752),
.C(n_817),
.Y(n_930)
);

BUFx8_ASAP7_75t_L g931 ( 
.A(n_825),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_760),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_834),
.A2(n_823),
.B(n_816),
.C(n_819),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_804),
.A2(n_794),
.B(n_795),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_768),
.B(n_772),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_L g936 ( 
.A(n_673),
.B(n_721),
.C(n_734),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_780),
.A2(n_759),
.B(n_726),
.Y(n_937)
);

BUFx12f_ASAP7_75t_L g938 ( 
.A(n_751),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_715),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_765),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_804),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_804),
.A2(n_798),
.B(n_808),
.Y(n_942)
);

AOI21x1_ASAP7_75t_L g943 ( 
.A1(n_690),
.A2(n_735),
.B(n_780),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_692),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_693),
.A2(n_750),
.B1(n_757),
.B2(n_826),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_804),
.A2(n_735),
.B(n_830),
.Y(n_946)
);

BUFx8_ASAP7_75t_L g947 ( 
.A(n_825),
.Y(n_947)
);

OR2x6_ASAP7_75t_SL g948 ( 
.A(n_793),
.B(n_807),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_731),
.B(n_723),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_750),
.A2(n_757),
.B1(n_724),
.B2(n_826),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_723),
.B(n_716),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_724),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_724),
.A2(n_826),
.B1(n_806),
.B2(n_740),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_777),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_784),
.Y(n_955)
);

CKINVDCx10_ASAP7_75t_R g956 ( 
.A(n_745),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_827),
.A2(n_828),
.B(n_791),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_733),
.A2(n_821),
.B(n_705),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_687),
.A2(n_736),
.B(n_783),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_683),
.B(n_774),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_802),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_817),
.B(n_824),
.Y(n_962)
);

AOI33xp33_ASAP7_75t_L g963 ( 
.A1(n_706),
.A2(n_716),
.A3(n_740),
.B1(n_815),
.B2(n_799),
.B3(n_833),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_769),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_706),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_713),
.B(n_519),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_SL g967 ( 
.A1(n_674),
.A2(n_834),
.B(n_795),
.C(n_808),
.Y(n_967)
);

AND2x2_ASAP7_75t_SL g968 ( 
.A(n_693),
.B(n_601),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_697),
.A2(n_581),
.B(n_568),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_672),
.B(n_707),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_697),
.A2(n_581),
.B(n_568),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_672),
.A2(n_703),
.B(n_700),
.C(n_707),
.Y(n_972)
);

AND2x6_ASAP7_75t_L g973 ( 
.A(n_814),
.B(n_675),
.Y(n_973)
);

AOI22x1_ASAP7_75t_L g974 ( 
.A1(n_675),
.A2(n_615),
.B1(n_633),
.B2(n_613),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_672),
.B(n_707),
.Y(n_975)
);

BUFx4f_ASAP7_75t_L g976 ( 
.A(n_725),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_672),
.B(n_707),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_697),
.A2(n_581),
.B(n_568),
.Y(n_978)
);

BUFx2_ASAP7_75t_SL g979 ( 
.A(n_751),
.Y(n_979)
);

INVx5_ASAP7_75t_L g980 ( 
.A(n_724),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_713),
.B(n_519),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_672),
.B(n_805),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_672),
.B(n_805),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_697),
.A2(n_581),
.B(n_568),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_672),
.B(n_707),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_672),
.B(n_805),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_672),
.B(n_805),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_L g988 ( 
.A(n_673),
.B(n_672),
.C(n_700),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_679),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_697),
.A2(n_581),
.B(n_568),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_713),
.A2(n_672),
.B1(n_814),
.B2(n_676),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_809),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_672),
.B(n_707),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_672),
.B(n_707),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_781),
.B(n_831),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_804),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_672),
.B(n_805),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_804),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_697),
.A2(n_581),
.B(n_568),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_809),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_697),
.A2(n_581),
.B(n_568),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_697),
.A2(n_581),
.B(n_568),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_679),
.Y(n_1003)
);

INVx4_ASAP7_75t_L g1004 ( 
.A(n_804),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_713),
.A2(n_672),
.B1(n_814),
.B2(n_676),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_762),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_810),
.A2(n_672),
.B1(n_813),
.B2(n_812),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_672),
.A2(n_810),
.B(n_813),
.C(n_812),
.Y(n_1008)
);

AOI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_672),
.A2(n_810),
.B(n_703),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_809),
.Y(n_1010)
);

O2A1O1Ixp5_ASAP7_75t_L g1011 ( 
.A1(n_702),
.A2(n_672),
.B(n_686),
.C(n_674),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_809),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_672),
.B(n_805),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_672),
.B(n_707),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_713),
.B(n_519),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_713),
.B(n_519),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_672),
.B(n_805),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_713),
.B(n_519),
.Y(n_1018)
);

NOR3xp33_ASAP7_75t_L g1019 ( 
.A(n_673),
.B(n_672),
.C(n_700),
.Y(n_1019)
);

AOI21x1_ASAP7_75t_SL g1020 ( 
.A1(n_905),
.A2(n_985),
.B(n_970),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_878),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_975),
.B(n_977),
.Y(n_1022)
);

NAND2x1_ASAP7_75t_L g1023 ( 
.A(n_1004),
.B(n_952),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_862),
.A2(n_908),
.B(n_913),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_941),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_883),
.Y(n_1026)
);

AOI21xp33_ASAP7_75t_L g1027 ( 
.A1(n_1008),
.A2(n_1007),
.B(n_889),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_859),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_970),
.B(n_985),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_853),
.A2(n_902),
.B(n_901),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_944),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_841),
.A2(n_972),
.B(n_1009),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_969),
.A2(n_978),
.B(n_971),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_903),
.A2(n_934),
.B(n_844),
.Y(n_1034)
);

INVx2_ASAP7_75t_SL g1035 ( 
.A(n_874),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_984),
.A2(n_999),
.B(n_990),
.Y(n_1036)
);

AO31x2_ASAP7_75t_L g1037 ( 
.A1(n_991),
.A2(n_1005),
.A3(n_860),
.B(n_930),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_875),
.A2(n_942),
.B(n_851),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_1009),
.A2(n_993),
.B(n_994),
.C(n_1014),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_993),
.A2(n_994),
.B1(n_1014),
.B2(n_905),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_885),
.A2(n_1011),
.B(n_981),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_846),
.B(n_982),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_914),
.A2(n_852),
.B(n_921),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_941),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_924),
.A2(n_842),
.B(n_916),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_857),
.B(n_983),
.Y(n_1046)
);

AOI21x1_ASAP7_75t_SL g1047 ( 
.A1(n_891),
.A2(n_919),
.B(n_949),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_986),
.B(n_987),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_839),
.A2(n_870),
.B(n_911),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_854),
.A2(n_856),
.B(n_884),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_997),
.B(n_1013),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_849),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_880),
.B(n_872),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_863),
.B(n_1017),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_919),
.B(n_840),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_968),
.B(n_906),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_946),
.A2(n_882),
.B(n_943),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_840),
.B(n_846),
.Y(n_1058)
);

OR2x6_ASAP7_75t_L g1059 ( 
.A(n_979),
.B(n_938),
.Y(n_1059)
);

OA21x2_ASAP7_75t_L g1060 ( 
.A1(n_898),
.A2(n_957),
.B(n_876),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1001),
.A2(n_1002),
.B(n_925),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_923),
.A2(n_967),
.B(n_920),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_966),
.A2(n_1018),
.B(n_1016),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_899),
.B(n_915),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_910),
.A2(n_974),
.B(n_888),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_861),
.B(n_988),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1015),
.A2(n_918),
.B(n_879),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_1006),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_861),
.B(n_1019),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_886),
.A2(n_958),
.B(n_887),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_955),
.B(n_954),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_900),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_917),
.A2(n_879),
.B(n_876),
.Y(n_1073)
);

CKINVDCx8_ASAP7_75t_R g1074 ( 
.A(n_871),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_927),
.A2(n_960),
.B(n_933),
.C(n_945),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_941),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_926),
.A2(n_929),
.B(n_855),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_936),
.A2(n_951),
.B(n_845),
.C(n_937),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_973),
.A2(n_866),
.B(n_873),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_973),
.A2(n_866),
.B(n_873),
.Y(n_1080)
);

AOI21x1_ASAP7_75t_L g1081 ( 
.A1(n_891),
.A2(n_858),
.B(n_848),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_858),
.A2(n_848),
.B(n_855),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_931),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_900),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_973),
.B(n_965),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_850),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_953),
.A2(n_950),
.B(n_980),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_962),
.A2(n_912),
.B1(n_890),
.B2(n_881),
.Y(n_1088)
);

NAND2x1p5_ASAP7_75t_L g1089 ( 
.A(n_980),
.B(n_952),
.Y(n_1089)
);

NOR3xp33_ASAP7_75t_L g1090 ( 
.A(n_897),
.B(n_951),
.C(n_847),
.Y(n_1090)
);

AOI21x1_ASAP7_75t_L g1091 ( 
.A1(n_926),
.A2(n_929),
.B(n_1012),
.Y(n_1091)
);

AOI21xp33_ASAP7_75t_L g1092 ( 
.A1(n_962),
.A2(n_961),
.B(n_949),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_980),
.A2(n_935),
.B(n_959),
.Y(n_1093)
);

INVx5_ASAP7_75t_L g1094 ( 
.A(n_973),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_973),
.A2(n_964),
.B(n_867),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_922),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_935),
.A2(n_996),
.B(n_998),
.Y(n_1097)
);

O2A1O1Ixp5_ASAP7_75t_L g1098 ( 
.A1(n_868),
.A2(n_892),
.B(n_896),
.C(n_893),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_948),
.B(n_864),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_895),
.A2(n_998),
.B(n_996),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_865),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_869),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_992),
.A2(n_1010),
.B(n_1000),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_904),
.B(n_907),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1004),
.A2(n_1003),
.B(n_989),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_976),
.B(n_877),
.Y(n_1106)
);

AO31x2_ASAP7_75t_L g1107 ( 
.A1(n_932),
.A2(n_939),
.A3(n_894),
.B(n_963),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_976),
.B(n_940),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_909),
.A2(n_928),
.B(n_922),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_909),
.A2(n_995),
.B(n_947),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_995),
.A2(n_931),
.B(n_947),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_956),
.B(n_1007),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_SL g1113 ( 
.A1(n_1008),
.A2(n_933),
.B(n_892),
.Y(n_1113)
);

AO21x2_ASAP7_75t_L g1114 ( 
.A1(n_1009),
.A2(n_898),
.B(n_841),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_941),
.Y(n_1115)
);

AOI221xp5_ASAP7_75t_SL g1116 ( 
.A1(n_1008),
.A2(n_1007),
.B1(n_841),
.B2(n_972),
.C(n_977),
.Y(n_1116)
);

NAND3xp33_ASAP7_75t_SL g1117 ( 
.A(n_988),
.B(n_1019),
.C(n_1007),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_841),
.A2(n_972),
.B(n_1008),
.C(n_1009),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_862),
.A2(n_908),
.B(n_913),
.Y(n_1119)
);

AO21x1_ASAP7_75t_L g1120 ( 
.A1(n_1009),
.A2(n_1008),
.B(n_985),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_928),
.B(n_940),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_975),
.B(n_977),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_975),
.B(n_977),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_975),
.B(n_977),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_975),
.B(n_977),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_862),
.A2(n_908),
.B(n_913),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_975),
.B(n_977),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_843),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_880),
.B(n_872),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1007),
.B(n_905),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_843),
.Y(n_1131)
);

OAI21xp33_ASAP7_75t_L g1132 ( 
.A1(n_1007),
.A2(n_672),
.B(n_693),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_969),
.A2(n_568),
.B(n_581),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_975),
.B(n_977),
.Y(n_1134)
);

INVxp67_ASAP7_75t_SL g1135 ( 
.A(n_941),
.Y(n_1135)
);

NOR2xp67_ASAP7_75t_SL g1136 ( 
.A(n_980),
.B(n_979),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_862),
.A2(n_908),
.B(n_913),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_975),
.B(n_977),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_975),
.B(n_977),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_859),
.Y(n_1140)
);

INVx4_ASAP7_75t_L g1141 ( 
.A(n_941),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_944),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_970),
.A2(n_993),
.B1(n_994),
.B2(n_985),
.Y(n_1143)
);

OAI22x1_ASAP7_75t_L g1144 ( 
.A1(n_889),
.A2(n_857),
.B1(n_822),
.B2(n_863),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_941),
.Y(n_1145)
);

AOI21xp33_ASAP7_75t_L g1146 ( 
.A1(n_1008),
.A2(n_1007),
.B(n_889),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_944),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_975),
.B(n_977),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_975),
.B(n_977),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_988),
.A2(n_1019),
.B1(n_672),
.B2(n_977),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_969),
.A2(n_568),
.B(n_581),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_841),
.A2(n_972),
.B(n_1008),
.Y(n_1152)
);

AO32x2_ASAP7_75t_L g1153 ( 
.A1(n_991),
.A2(n_1005),
.A3(n_945),
.B1(n_845),
.B2(n_953),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_944),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_841),
.A2(n_972),
.B(n_1008),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_880),
.B(n_872),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_841),
.A2(n_972),
.B(n_1008),
.C(n_1009),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_862),
.A2(n_908),
.B(n_913),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_862),
.A2(n_908),
.B(n_913),
.Y(n_1159)
);

NAND2xp33_ASAP7_75t_L g1160 ( 
.A(n_841),
.B(n_972),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_975),
.B(n_977),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_975),
.B(n_977),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_980),
.B(n_952),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_975),
.B(n_977),
.Y(n_1164)
);

OAI22x1_ASAP7_75t_L g1165 ( 
.A1(n_889),
.A2(n_857),
.B1(n_822),
.B2(n_863),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_841),
.A2(n_972),
.B(n_1008),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_862),
.A2(n_908),
.B(n_913),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_841),
.A2(n_972),
.B(n_1008),
.Y(n_1168)
);

INVx5_ASAP7_75t_L g1169 ( 
.A(n_1025),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1026),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_1021),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_1142),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1053),
.B(n_1129),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_1142),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1156),
.B(n_1054),
.Y(n_1175)
);

NOR2xp67_ASAP7_75t_L g1176 ( 
.A(n_1028),
.B(n_1140),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1110),
.B(n_1109),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1134),
.B(n_1149),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1061),
.A2(n_1160),
.B(n_1062),
.Y(n_1179)
);

AOI221xp5_ASAP7_75t_L g1180 ( 
.A1(n_1132),
.A2(n_1146),
.B1(n_1027),
.B2(n_1143),
.C(n_1040),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1143),
.B(n_1029),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1040),
.B(n_1039),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1121),
.B(n_1096),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1056),
.B(n_1046),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1064),
.B(n_1072),
.Y(n_1185)
);

NAND4xp25_ASAP7_75t_L g1186 ( 
.A(n_1099),
.B(n_1071),
.C(n_1112),
.D(n_1084),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1031),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1022),
.B(n_1122),
.Y(n_1188)
);

BUFx12f_ASAP7_75t_L g1189 ( 
.A(n_1059),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_1154),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1022),
.B(n_1122),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1074),
.Y(n_1192)
);

CKINVDCx8_ASAP7_75t_R g1193 ( 
.A(n_1147),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1121),
.B(n_1096),
.Y(n_1194)
);

BUFx12f_ASAP7_75t_L g1195 ( 
.A(n_1059),
.Y(n_1195)
);

CKINVDCx11_ASAP7_75t_R g1196 ( 
.A(n_1083),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1123),
.B(n_1124),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1117),
.A2(n_1146),
.B1(n_1027),
.B2(n_1166),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1123),
.B(n_1124),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1125),
.B(n_1127),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1125),
.B(n_1127),
.Y(n_1201)
);

INVx5_ASAP7_75t_L g1202 ( 
.A(n_1025),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1138),
.B(n_1139),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1148),
.B(n_1161),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1096),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1138),
.B(n_1139),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1162),
.B(n_1164),
.Y(n_1207)
);

AOI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1081),
.A2(n_1091),
.B(n_1087),
.Y(n_1208)
);

AOI222xp33_ASAP7_75t_L g1209 ( 
.A1(n_1152),
.A2(n_1166),
.B1(n_1155),
.B2(n_1168),
.C1(n_1130),
.C2(n_1032),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1152),
.A2(n_1168),
.B1(n_1155),
.B2(n_1120),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1150),
.B(n_1162),
.Y(n_1211)
);

AOI211xp5_ASAP7_75t_L g1212 ( 
.A1(n_1075),
.A2(n_1078),
.B(n_1157),
.C(n_1118),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1101),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1033),
.A2(n_1036),
.B(n_1073),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1035),
.B(n_1108),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1104),
.Y(n_1216)
);

NOR2xp67_ASAP7_75t_L g1217 ( 
.A(n_1144),
.B(n_1165),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1032),
.A2(n_1106),
.B1(n_1090),
.B2(n_1092),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1107),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1088),
.A2(n_1116),
.B1(n_1069),
.B2(n_1066),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1052),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1164),
.B(n_1055),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1048),
.B(n_1051),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_SL g1224 ( 
.A1(n_1094),
.A2(n_1114),
.B1(n_1113),
.B2(n_1095),
.Y(n_1224)
);

CKINVDCx12_ASAP7_75t_R g1225 ( 
.A(n_1059),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1066),
.A2(n_1069),
.B(n_1042),
.C(n_1092),
.Y(n_1226)
);

BUFx12f_ASAP7_75t_L g1227 ( 
.A(n_1025),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1044),
.Y(n_1228)
);

BUFx2_ASAP7_75t_SL g1229 ( 
.A(n_1044),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1114),
.A2(n_1085),
.B1(n_1095),
.B2(n_1079),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1082),
.A2(n_1151),
.B(n_1133),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1086),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1107),
.B(n_1102),
.Y(n_1233)
);

OR2x6_ASAP7_75t_L g1234 ( 
.A(n_1111),
.B(n_1163),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1042),
.B(n_1058),
.Y(n_1235)
);

CKINVDCx6p67_ASAP7_75t_R g1236 ( 
.A(n_1044),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1128),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_1085),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1131),
.B(n_1094),
.Y(n_1239)
);

INVx2_ASAP7_75t_SL g1240 ( 
.A(n_1115),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1145),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1145),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1079),
.A2(n_1080),
.B1(n_1094),
.B2(n_1067),
.Y(n_1243)
);

OR2x6_ASAP7_75t_L g1244 ( 
.A(n_1089),
.B(n_1163),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1080),
.A2(n_1094),
.B1(n_1103),
.B2(n_1041),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1067),
.A2(n_1041),
.B(n_1063),
.C(n_1098),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1089),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1103),
.Y(n_1248)
);

BUFx12f_ASAP7_75t_L g1249 ( 
.A(n_1141),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1077),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1076),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1135),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_SL g1253 ( 
.A1(n_1060),
.A2(n_1093),
.B(n_1097),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_1141),
.B(n_1023),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1060),
.A2(n_1105),
.B(n_1153),
.C(n_1020),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1037),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1100),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1045),
.A2(n_1050),
.B(n_1049),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1030),
.Y(n_1259)
);

OAI21xp33_ASAP7_75t_L g1260 ( 
.A1(n_1153),
.A2(n_1057),
.B(n_1038),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1034),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1024),
.B(n_1126),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1119),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1043),
.B(n_1137),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1158),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1065),
.B(n_1159),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1167),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1047),
.B(n_1053),
.Y(n_1268)
);

O2A1O1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1132),
.A2(n_841),
.B(n_972),
.C(n_1009),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1110),
.B(n_1109),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1110),
.B(n_1109),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1132),
.A2(n_841),
.B(n_972),
.C(n_1008),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1154),
.Y(n_1273)
);

A2O1A1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1132),
.A2(n_841),
.B(n_972),
.C(n_1008),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1134),
.B(n_1149),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1061),
.A2(n_568),
.B(n_1160),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1068),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1028),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1134),
.B(n_1149),
.Y(n_1279)
);

CKINVDCx20_ASAP7_75t_R g1280 ( 
.A(n_1074),
.Y(n_1280)
);

NAND2x1p5_ASAP7_75t_L g1281 ( 
.A(n_1136),
.B(n_1004),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1053),
.B(n_1129),
.Y(n_1282)
);

NAND2x1p5_ASAP7_75t_L g1283 ( 
.A(n_1136),
.B(n_1004),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1025),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1132),
.A2(n_841),
.B(n_972),
.C(n_1008),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1134),
.B(n_1149),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1053),
.B(n_1129),
.Y(n_1287)
);

BUFx4f_ASAP7_75t_L g1288 ( 
.A(n_1059),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1132),
.A2(n_841),
.B(n_972),
.C(n_1009),
.Y(n_1289)
);

OR2x2_ASAP7_75t_SL g1290 ( 
.A(n_1117),
.B(n_673),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1134),
.B(n_1149),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1134),
.B(n_1149),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1061),
.A2(n_568),
.B(n_1160),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1053),
.B(n_1129),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1134),
.B(n_1149),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1110),
.B(n_1109),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1154),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1154),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1030),
.A2(n_1070),
.B(n_1024),
.Y(n_1299)
);

CKINVDCx16_ASAP7_75t_R g1300 ( 
.A(n_1083),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1053),
.B(n_1129),
.Y(n_1301)
);

BUFx2_ASAP7_75t_R g1302 ( 
.A(n_1278),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_SL g1303 ( 
.A1(n_1198),
.A2(n_1209),
.B(n_1269),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1178),
.A2(n_1291),
.B1(n_1295),
.B2(n_1286),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1299),
.A2(n_1258),
.B(n_1179),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1178),
.A2(n_1292),
.B1(n_1275),
.B2(n_1286),
.Y(n_1306)
);

BUFx4f_ASAP7_75t_SL g1307 ( 
.A(n_1280),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1196),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1275),
.A2(n_1292),
.B1(n_1291),
.B2(n_1279),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_SL g1310 ( 
.A(n_1273),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1211),
.A2(n_1209),
.B1(n_1180),
.B2(n_1279),
.Y(n_1311)
);

INVxp67_ASAP7_75t_SL g1312 ( 
.A(n_1277),
.Y(n_1312)
);

CKINVDCx11_ASAP7_75t_R g1313 ( 
.A(n_1193),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1295),
.A2(n_1184),
.B1(n_1204),
.B2(n_1288),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1180),
.A2(n_1210),
.B1(n_1218),
.B2(n_1220),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_SL g1316 ( 
.A1(n_1288),
.A2(n_1206),
.B1(n_1207),
.B2(n_1191),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1233),
.Y(n_1317)
);

OA21x2_ASAP7_75t_L g1318 ( 
.A1(n_1179),
.A2(n_1214),
.B(n_1231),
.Y(n_1318)
);

CKINVDCx11_ASAP7_75t_R g1319 ( 
.A(n_1300),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1169),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1259),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1177),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1177),
.Y(n_1323)
);

INVx1_ASAP7_75t_SL g1324 ( 
.A(n_1172),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_1172),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1258),
.A2(n_1231),
.B(n_1214),
.Y(n_1326)
);

CKINVDCx11_ASAP7_75t_R g1327 ( 
.A(n_1189),
.Y(n_1327)
);

OR2x6_ASAP7_75t_SL g1328 ( 
.A(n_1192),
.B(n_1223),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1276),
.A2(n_1293),
.B(n_1266),
.Y(n_1329)
);

AO21x1_ASAP7_75t_L g1330 ( 
.A1(n_1269),
.A2(n_1289),
.B(n_1212),
.Y(n_1330)
);

AO21x1_ASAP7_75t_L g1331 ( 
.A1(n_1289),
.A2(n_1181),
.B(n_1226),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1175),
.B(n_1173),
.Y(n_1332)
);

AO21x2_ASAP7_75t_L g1333 ( 
.A1(n_1276),
.A2(n_1293),
.B(n_1266),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1185),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1282),
.B(n_1301),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1182),
.A2(n_1217),
.B1(n_1181),
.B2(n_1191),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1171),
.Y(n_1337)
);

OAI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1188),
.A2(n_1206),
.B1(n_1200),
.B2(n_1199),
.Y(n_1338)
);

AOI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1208),
.A2(n_1182),
.B(n_1262),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1188),
.A2(n_1199),
.B1(n_1200),
.B2(n_1207),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1197),
.A2(n_1203),
.B1(n_1201),
.B2(n_1186),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1197),
.B(n_1201),
.Y(n_1342)
);

OA21x2_ASAP7_75t_L g1343 ( 
.A1(n_1246),
.A2(n_1260),
.B(n_1243),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1203),
.A2(n_1222),
.B1(n_1235),
.B2(n_1216),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1287),
.B(n_1294),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1239),
.B(n_1270),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1297),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1222),
.A2(n_1235),
.B1(n_1248),
.B2(n_1268),
.Y(n_1348)
);

INVx2_ASAP7_75t_SL g1349 ( 
.A(n_1298),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1290),
.A2(n_1238),
.B1(n_1272),
.B2(n_1274),
.Y(n_1350)
);

INVx1_ASAP7_75t_SL g1351 ( 
.A(n_1174),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1226),
.B(n_1285),
.Y(n_1352)
);

AOI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1263),
.A2(n_1257),
.B(n_1267),
.Y(n_1353)
);

OAI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1245),
.A2(n_1234),
.B1(n_1232),
.B2(n_1237),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1221),
.Y(n_1355)
);

BUFx12f_ASAP7_75t_L g1356 ( 
.A(n_1195),
.Y(n_1356)
);

INVxp67_ASAP7_75t_SL g1357 ( 
.A(n_1252),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1250),
.A2(n_1255),
.B(n_1253),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1256),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1219),
.Y(n_1360)
);

AOI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1264),
.A2(n_1296),
.B(n_1271),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_SL g1362 ( 
.A1(n_1281),
.A2(n_1283),
.B(n_1239),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1213),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1202),
.B(n_1296),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1224),
.A2(n_1215),
.B1(n_1230),
.B2(n_1187),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1224),
.A2(n_1215),
.B1(n_1234),
.B2(n_1183),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1183),
.B(n_1194),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1194),
.B(n_1190),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1205),
.B(n_1176),
.Y(n_1369)
);

CKINVDCx11_ASAP7_75t_R g1370 ( 
.A(n_1249),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1270),
.B(n_1271),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1284),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_SL g1373 ( 
.A1(n_1247),
.A2(n_1251),
.B1(n_1254),
.B2(n_1229),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1284),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1284),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1281),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1234),
.B(n_1242),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1244),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1228),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1240),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1241),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1236),
.Y(n_1382)
);

CKINVDCx8_ASAP7_75t_R g1383 ( 
.A(n_1244),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1225),
.A2(n_1261),
.B1(n_1265),
.B2(n_1264),
.Y(n_1384)
);

INVx2_ASAP7_75t_SL g1385 ( 
.A(n_1261),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1277),
.Y(n_1386)
);

BUFx2_ASAP7_75t_SL g1387 ( 
.A(n_1280),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1178),
.A2(n_968),
.B1(n_601),
.B2(n_825),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1198),
.A2(n_972),
.B(n_841),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1178),
.A2(n_977),
.B1(n_975),
.B2(n_970),
.Y(n_1390)
);

BUFx10_ASAP7_75t_L g1391 ( 
.A(n_1278),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1172),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1198),
.A2(n_1132),
.B1(n_968),
.B2(n_889),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1170),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1196),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_1172),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1227),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1175),
.B(n_1173),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1198),
.A2(n_1132),
.B1(n_968),
.B2(n_889),
.Y(n_1399)
);

BUFx2_ASAP7_75t_R g1400 ( 
.A(n_1278),
.Y(n_1400)
);

CKINVDCx11_ASAP7_75t_R g1401 ( 
.A(n_1196),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1178),
.A2(n_977),
.B1(n_975),
.B2(n_970),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1383),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1361),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1389),
.A2(n_1311),
.B(n_1393),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1350),
.A2(n_1315),
.B1(n_1393),
.B2(n_1399),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1317),
.B(n_1343),
.Y(n_1407)
);

OAI21xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1315),
.A2(n_1311),
.B(n_1352),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1371),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1305),
.A2(n_1329),
.B(n_1326),
.Y(n_1410)
);

AO31x2_ASAP7_75t_L g1411 ( 
.A1(n_1331),
.A2(n_1330),
.A3(n_1360),
.B(n_1359),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1318),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1343),
.B(n_1348),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1348),
.B(n_1343),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1332),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1353),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1371),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1371),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1365),
.B(n_1303),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1358),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1386),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1322),
.B(n_1323),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1358),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1339),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1383),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1318),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1333),
.Y(n_1427)
);

INVxp67_ASAP7_75t_L g1428 ( 
.A(n_1335),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1322),
.B(n_1323),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1323),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1398),
.B(n_1345),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1304),
.B(n_1306),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1399),
.A2(n_1336),
.B(n_1344),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1307),
.B(n_1334),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1340),
.B(n_1336),
.Y(n_1435)
);

INVxp67_ASAP7_75t_L g1436 ( 
.A(n_1363),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1344),
.B(n_1342),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1321),
.Y(n_1438)
);

AO21x2_ASAP7_75t_L g1439 ( 
.A1(n_1354),
.A2(n_1309),
.B(n_1338),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1346),
.B(n_1341),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1341),
.B(n_1309),
.Y(n_1441)
);

CKINVDCx11_ASAP7_75t_R g1442 ( 
.A(n_1401),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1312),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_1324),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1325),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1394),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1338),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1355),
.A2(n_1385),
.B(n_1366),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1378),
.Y(n_1449)
);

OR2x6_ASAP7_75t_L g1450 ( 
.A(n_1362),
.B(n_1364),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1378),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1354),
.Y(n_1452)
);

OA21x2_ASAP7_75t_L g1453 ( 
.A1(n_1377),
.A2(n_1357),
.B(n_1376),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1364),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1384),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1316),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1314),
.B(n_1367),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1390),
.B(n_1402),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1351),
.B(n_1392),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1388),
.B(n_1396),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1337),
.B(n_1368),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1379),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1328),
.B(n_1369),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1453),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1437),
.B(n_1373),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1453),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1437),
.B(n_1374),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1407),
.B(n_1375),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1407),
.B(n_1372),
.Y(n_1469)
);

INVx4_ASAP7_75t_L g1470 ( 
.A(n_1450),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1413),
.B(n_1380),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1413),
.B(n_1381),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1414),
.B(n_1387),
.Y(n_1473)
);

INVx4_ASAP7_75t_L g1474 ( 
.A(n_1450),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1414),
.B(n_1347),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1405),
.A2(n_1319),
.B1(n_1327),
.B2(n_1310),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1443),
.Y(n_1477)
);

AOI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1406),
.A2(n_1310),
.B1(n_1356),
.B2(n_1319),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1432),
.B(n_1391),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1453),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1453),
.B(n_1349),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1422),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1447),
.B(n_1320),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1431),
.B(n_1307),
.Y(n_1484)
);

OR2x6_ASAP7_75t_L g1485 ( 
.A(n_1450),
.B(n_1404),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1416),
.B(n_1382),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1420),
.B(n_1397),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1447),
.B(n_1458),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1423),
.B(n_1427),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_SL g1490 ( 
.A1(n_1408),
.A2(n_1395),
.B1(n_1308),
.B2(n_1356),
.Y(n_1490)
);

OAI21xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1419),
.A2(n_1302),
.B(n_1400),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1438),
.Y(n_1492)
);

AOI221xp5_ASAP7_75t_L g1493 ( 
.A1(n_1408),
.A2(n_1397),
.B1(n_1308),
.B2(n_1395),
.C(n_1401),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1429),
.B(n_1327),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1430),
.B(n_1424),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1438),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1412),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1477),
.B(n_1421),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1490),
.A2(n_1419),
.B1(n_1441),
.B2(n_1456),
.Y(n_1499)
);

AOI221xp5_ASAP7_75t_L g1500 ( 
.A1(n_1493),
.A2(n_1456),
.B1(n_1436),
.B2(n_1460),
.C(n_1428),
.Y(n_1500)
);

OAI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1490),
.A2(n_1463),
.B(n_1435),
.Y(n_1501)
);

AND2x2_ASAP7_75t_SL g1502 ( 
.A(n_1470),
.B(n_1433),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1467),
.B(n_1435),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1472),
.B(n_1448),
.Y(n_1504)
);

OAI21xp5_ASAP7_75t_SL g1505 ( 
.A1(n_1493),
.A2(n_1460),
.B(n_1457),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1478),
.A2(n_1457),
.B(n_1455),
.Y(n_1506)
);

NOR3xp33_ASAP7_75t_L g1507 ( 
.A(n_1479),
.B(n_1434),
.C(n_1442),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1496),
.Y(n_1508)
);

NAND3xp33_ASAP7_75t_L g1509 ( 
.A(n_1473),
.B(n_1452),
.C(n_1440),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1471),
.B(n_1488),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1465),
.B(n_1409),
.Y(n_1511)
);

NAND3xp33_ASAP7_75t_L g1512 ( 
.A(n_1478),
.B(n_1440),
.C(n_1451),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1472),
.B(n_1448),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1465),
.B(n_1409),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1484),
.B(n_1415),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_L g1516 ( 
.A(n_1475),
.B(n_1451),
.C(n_1449),
.Y(n_1516)
);

AND2x2_ASAP7_75t_SL g1517 ( 
.A(n_1470),
.B(n_1433),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1468),
.B(n_1439),
.Y(n_1518)
);

OAI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1476),
.A2(n_1425),
.B1(n_1403),
.B2(n_1461),
.C(n_1444),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1491),
.A2(n_1425),
.B1(n_1403),
.B2(n_1433),
.Y(n_1520)
);

NAND3xp33_ASAP7_75t_L g1521 ( 
.A(n_1481),
.B(n_1451),
.C(n_1449),
.Y(n_1521)
);

NAND4xp25_ASAP7_75t_L g1522 ( 
.A(n_1486),
.B(n_1461),
.C(n_1459),
.D(n_1445),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1482),
.B(n_1411),
.Y(n_1523)
);

NAND3xp33_ASAP7_75t_L g1524 ( 
.A(n_1481),
.B(n_1454),
.C(n_1433),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1491),
.A2(n_1418),
.B(n_1417),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1466),
.Y(n_1526)
);

OA21x2_ASAP7_75t_L g1527 ( 
.A1(n_1480),
.A2(n_1410),
.B(n_1426),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1468),
.B(n_1439),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1469),
.B(n_1439),
.Y(n_1529)
);

OAI21xp5_ASAP7_75t_SL g1530 ( 
.A1(n_1494),
.A2(n_1417),
.B(n_1418),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1494),
.B(n_1459),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1469),
.B(n_1411),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1469),
.B(n_1411),
.Y(n_1533)
);

INVx2_ASAP7_75t_SL g1534 ( 
.A(n_1492),
.Y(n_1534)
);

OAI221xp5_ASAP7_75t_SL g1535 ( 
.A1(n_1485),
.A2(n_1425),
.B1(n_1403),
.B2(n_1462),
.C(n_1446),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1521),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1508),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1504),
.B(n_1513),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1526),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1527),
.Y(n_1540)
);

OR2x6_ASAP7_75t_L g1541 ( 
.A(n_1530),
.B(n_1485),
.Y(n_1541)
);

INVx4_ASAP7_75t_L g1542 ( 
.A(n_1502),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1523),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1502),
.B(n_1464),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1502),
.B(n_1464),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1517),
.B(n_1485),
.Y(n_1546)
);

AOI211xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1499),
.A2(n_1483),
.B(n_1494),
.C(n_1487),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1532),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1532),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1518),
.B(n_1480),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1533),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1517),
.B(n_1485),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1517),
.B(n_1489),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1528),
.B(n_1496),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1533),
.Y(n_1555)
);

NOR2xp67_ASAP7_75t_SL g1556 ( 
.A(n_1505),
.B(n_1470),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1534),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1529),
.B(n_1497),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1527),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1510),
.B(n_1495),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1550),
.B(n_1524),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1537),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1548),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1536),
.B(n_1503),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1553),
.B(n_1511),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1548),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1540),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1550),
.B(n_1498),
.Y(n_1568)
);

NAND2x1p5_ASAP7_75t_L g1569 ( 
.A(n_1556),
.B(n_1470),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1553),
.B(n_1511),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1549),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1553),
.B(n_1514),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1551),
.B(n_1538),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1560),
.B(n_1522),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1538),
.B(n_1531),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1557),
.Y(n_1576)
);

NAND2x1_ASAP7_75t_L g1577 ( 
.A(n_1542),
.B(n_1474),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1542),
.B(n_1474),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1540),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1555),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1558),
.Y(n_1581)
);

INVx2_ASAP7_75t_SL g1582 ( 
.A(n_1539),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1546),
.B(n_1516),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1542),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1546),
.B(n_1474),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_1537),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1539),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1567),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1573),
.B(n_1542),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1563),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1584),
.B(n_1541),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1573),
.B(n_1543),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_SL g1593 ( 
.A(n_1569),
.B(n_1556),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1576),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1561),
.B(n_1550),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1576),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1561),
.B(n_1554),
.Y(n_1597)
);

INVx3_ASAP7_75t_SL g1598 ( 
.A(n_1582),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1577),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1567),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1567),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1579),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1584),
.B(n_1543),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1579),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1584),
.B(n_1543),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1562),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1584),
.B(n_1544),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1566),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1577),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1579),
.Y(n_1610)
);

INVx1_ASAP7_75t_SL g1611 ( 
.A(n_1582),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1583),
.B(n_1544),
.Y(n_1612)
);

INVx2_ASAP7_75t_SL g1613 ( 
.A(n_1587),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1568),
.B(n_1554),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1568),
.B(n_1554),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1571),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1583),
.B(n_1544),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1574),
.B(n_1370),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1583),
.B(n_1545),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1583),
.B(n_1545),
.Y(n_1620)
);

AOI32xp33_ASAP7_75t_L g1621 ( 
.A1(n_1586),
.A2(n_1547),
.A3(n_1500),
.B1(n_1520),
.B2(n_1507),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1580),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1606),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1622),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1598),
.Y(n_1625)
);

INVx1_ASAP7_75t_SL g1626 ( 
.A(n_1606),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1621),
.B(n_1564),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1595),
.B(n_1564),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1621),
.B(n_1565),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1622),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1613),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1613),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1613),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1589),
.B(n_1585),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1618),
.A2(n_1556),
.B1(n_1585),
.B2(n_1546),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1595),
.B(n_1565),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1598),
.A2(n_1506),
.B1(n_1569),
.B2(n_1525),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1597),
.B(n_1370),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1598),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1595),
.B(n_1581),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1611),
.B(n_1570),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1589),
.B(n_1585),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1616),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1616),
.Y(n_1644)
);

AOI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1593),
.A2(n_1501),
.B1(n_1519),
.B2(n_1512),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1592),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1590),
.Y(n_1647)
);

OAI21x1_ASAP7_75t_L g1648 ( 
.A1(n_1599),
.A2(n_1569),
.B(n_1559),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1611),
.B(n_1570),
.Y(n_1649)
);

INVx1_ASAP7_75t_SL g1650 ( 
.A(n_1594),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1593),
.B(n_1585),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1612),
.B(n_1572),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1612),
.B(n_1572),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1594),
.A2(n_1541),
.B1(n_1535),
.B2(n_1509),
.Y(n_1654)
);

NAND2xp33_ASAP7_75t_L g1655 ( 
.A(n_1596),
.B(n_1587),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1591),
.A2(n_1552),
.B1(n_1578),
.B2(n_1541),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1612),
.B(n_1575),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1625),
.B(n_1589),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1625),
.B(n_1592),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1624),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1645),
.A2(n_1591),
.B1(n_1578),
.B2(n_1617),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1645),
.A2(n_1541),
.B1(n_1596),
.B2(n_1609),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1631),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1623),
.B(n_1617),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1634),
.B(n_1592),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1624),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1630),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1626),
.Y(n_1668)
);

NAND3xp33_ASAP7_75t_SL g1669 ( 
.A(n_1627),
.B(n_1547),
.C(n_1597),
.Y(n_1669)
);

O2A1O1Ixp33_ASAP7_75t_L g1670 ( 
.A1(n_1655),
.A2(n_1609),
.B(n_1599),
.C(n_1617),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1630),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1647),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1647),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1643),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1631),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1634),
.B(n_1619),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1643),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1650),
.B(n_1619),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1642),
.B(n_1619),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1642),
.B(n_1620),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1632),
.Y(n_1681)
);

OAI22xp33_ASAP7_75t_SL g1682 ( 
.A1(n_1629),
.A2(n_1609),
.B1(n_1599),
.B2(n_1614),
.Y(n_1682)
);

AOI21xp33_ASAP7_75t_SL g1683 ( 
.A1(n_1651),
.A2(n_1599),
.B(n_1614),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1668),
.B(n_1639),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1664),
.B(n_1638),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1659),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1659),
.B(n_1655),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1658),
.B(n_1641),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1660),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1678),
.B(n_1657),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1669),
.B(n_1636),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1676),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1662),
.A2(n_1637),
.B1(n_1654),
.B2(n_1635),
.Y(n_1693)
);

BUFx3_ASAP7_75t_L g1694 ( 
.A(n_1658),
.Y(n_1694)
);

NAND2xp33_ASAP7_75t_SL g1695 ( 
.A(n_1676),
.B(n_1628),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1660),
.Y(n_1696)
);

INVxp67_ASAP7_75t_L g1697 ( 
.A(n_1663),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1666),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1665),
.B(n_1679),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1665),
.B(n_1679),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1680),
.B(n_1649),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1682),
.B(n_1652),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1680),
.B(n_1646),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1695),
.A2(n_1670),
.B(n_1683),
.Y(n_1704)
);

OAI211xp5_ASAP7_75t_L g1705 ( 
.A1(n_1702),
.A2(n_1661),
.B(n_1667),
.C(n_1666),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1702),
.A2(n_1675),
.B(n_1663),
.Y(n_1706)
);

NAND2xp33_ASAP7_75t_R g1707 ( 
.A(n_1686),
.B(n_1684),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1687),
.A2(n_1681),
.B(n_1675),
.Y(n_1708)
);

OAI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1693),
.A2(n_1656),
.B1(n_1628),
.B2(n_1646),
.C(n_1681),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1685),
.B(n_1653),
.Y(n_1710)
);

NAND3xp33_ASAP7_75t_SL g1711 ( 
.A(n_1691),
.B(n_1685),
.C(n_1688),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1694),
.B(n_1620),
.Y(n_1712)
);

AOI222xp33_ASAP7_75t_L g1713 ( 
.A1(n_1690),
.A2(n_1677),
.B1(n_1674),
.B2(n_1671),
.C1(n_1667),
.C2(n_1673),
.Y(n_1713)
);

AOI31xp33_ASAP7_75t_L g1714 ( 
.A1(n_1697),
.A2(n_1674),
.A3(n_1677),
.B(n_1671),
.Y(n_1714)
);

INVxp67_ASAP7_75t_SL g1715 ( 
.A(n_1697),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1712),
.B(n_1692),
.Y(n_1716)
);

NOR2x1_ASAP7_75t_L g1717 ( 
.A(n_1711),
.B(n_1689),
.Y(n_1717)
);

AOI211x1_ASAP7_75t_L g1718 ( 
.A1(n_1705),
.A2(n_1704),
.B(n_1706),
.C(n_1709),
.Y(n_1718)
);

NOR2xp67_ASAP7_75t_L g1719 ( 
.A(n_1708),
.B(n_1633),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1710),
.B(n_1699),
.Y(n_1720)
);

AOI211x1_ASAP7_75t_L g1721 ( 
.A1(n_1714),
.A2(n_1700),
.B(n_1701),
.C(n_1703),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1715),
.B(n_1696),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1707),
.A2(n_1632),
.B1(n_1591),
.B2(n_1698),
.Y(n_1723)
);

NAND4xp25_ASAP7_75t_L g1724 ( 
.A(n_1713),
.B(n_1672),
.C(n_1644),
.D(n_1640),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1711),
.B(n_1640),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1723),
.B(n_1620),
.Y(n_1726)
);

AND4x1_ASAP7_75t_L g1727 ( 
.A(n_1717),
.B(n_1644),
.C(n_1313),
.D(n_1603),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1719),
.B(n_1607),
.Y(n_1728)
);

O2A1O1Ixp33_ASAP7_75t_L g1729 ( 
.A1(n_1725),
.A2(n_1591),
.B(n_1603),
.C(n_1605),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1720),
.B(n_1716),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1726),
.B(n_1722),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1730),
.B(n_1718),
.Y(n_1732)
);

NOR2x1_ASAP7_75t_L g1733 ( 
.A(n_1728),
.B(n_1724),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1729),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1727),
.Y(n_1735)
);

NOR3xp33_ASAP7_75t_L g1736 ( 
.A(n_1730),
.B(n_1313),
.C(n_1721),
.Y(n_1736)
);

NOR3xp33_ASAP7_75t_L g1737 ( 
.A(n_1735),
.B(n_1648),
.C(n_1515),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1731),
.B(n_1591),
.Y(n_1738)
);

NAND4xp25_ASAP7_75t_L g1739 ( 
.A(n_1736),
.B(n_1607),
.C(n_1603),
.D(n_1605),
.Y(n_1739)
);

NAND3xp33_ASAP7_75t_SL g1740 ( 
.A(n_1732),
.B(n_1605),
.C(n_1615),
.Y(n_1740)
);

NOR2x1_ASAP7_75t_L g1741 ( 
.A(n_1733),
.B(n_1590),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1738),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1741),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1737),
.A2(n_1734),
.B1(n_1615),
.B2(n_1608),
.Y(n_1744)
);

INVxp67_ASAP7_75t_L g1745 ( 
.A(n_1743),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1745),
.B(n_1742),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1746),
.A2(n_1740),
.B1(n_1739),
.B2(n_1744),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1746),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1748),
.A2(n_1648),
.B(n_1600),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1747),
.A2(n_1600),
.B1(n_1602),
.B2(n_1601),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1750),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1749),
.Y(n_1752)
);

OAI21xp33_ASAP7_75t_SL g1753 ( 
.A1(n_1752),
.A2(n_1600),
.B(n_1588),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1753),
.A2(n_1751),
.B1(n_1588),
.B2(n_1601),
.Y(n_1754)
);

AOI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1754),
.A2(n_1602),
.B1(n_1601),
.B2(n_1604),
.C(n_1610),
.Y(n_1755)
);

AOI211xp5_ASAP7_75t_L g1756 ( 
.A1(n_1755),
.A2(n_1604),
.B(n_1610),
.C(n_1602),
.Y(n_1756)
);


endmodule