module fake_jpeg_23754_n_133 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_133);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_1),
.Y(n_63)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_28),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_24),
.B1(n_14),
.B2(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_42),
.Y(n_49)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_16),
.C(n_28),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_63),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_59),
.B(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_25),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_19),
.C(n_22),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_21),
.B1(n_15),
.B2(n_24),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_39),
.B1(n_14),
.B2(n_31),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_29),
.B(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_2),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_67),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_62),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_71),
.B(n_79),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_47),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_42),
.B(n_34),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_42),
.B1(n_3),
.B2(n_4),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_55),
.B1(n_45),
.B2(n_48),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_58),
.B1(n_63),
.B2(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_54),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_81),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_6),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_90),
.Y(n_97)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_89),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_59),
.C(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_65),
.B(n_44),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_92),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_43),
.C(n_62),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_68),
.C(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_75),
.B(n_13),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_79),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_65),
.Y(n_98)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_99),
.B(n_106),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_70),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_83),
.C(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_70),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_105),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_64),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_77),
.B(n_73),
.Y(n_106)
);

NAND5xp2_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_87),
.C(n_91),
.D(n_83),
.E(n_86),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_112),
.B(n_98),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_93),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_111),
.Y(n_121)
);

NOR2x1p5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_74),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_73),
.B1(n_74),
.B2(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_115),
.B(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_117),
.B(n_120),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_118),
.A2(n_108),
.B1(n_114),
.B2(n_109),
.Y(n_123)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_99),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_119),
.A2(n_118),
.B(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_126),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_124),
.B(n_125),
.Y(n_127)
);

AOI321xp33_ASAP7_75t_L g125 ( 
.A1(n_119),
.A2(n_109),
.A3(n_114),
.B1(n_92),
.B2(n_74),
.C(n_13),
.Y(n_125)
);

AOI321xp33_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_6),
.A3(n_8),
.B1(n_10),
.B2(n_12),
.C(n_82),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_107),
.Y(n_129)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_121),
.B(n_10),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_131),
.Y(n_132)
);

AOI21x1_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_127),
.B(n_128),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_12),
.Y(n_133)
);


endmodule