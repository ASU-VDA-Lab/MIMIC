module fake_jpeg_3760_n_291 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_291);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx24_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_2),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_16),
.B1(n_13),
.B2(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_16),
.B1(n_22),
.B2(n_25),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_48),
.B1(n_24),
.B2(n_13),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_35),
.B1(n_23),
.B2(n_18),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_22),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_20),
.B1(n_26),
.B2(n_25),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_20),
.C(n_26),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_20),
.B1(n_24),
.B2(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_28),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_57),
.B(n_23),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_15),
.Y(n_97)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_69),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

AO22x2_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_35),
.B1(n_33),
.B2(n_28),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_47),
.B1(n_53),
.B2(n_52),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_36),
.B1(n_43),
.B2(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_18),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_13),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_73),
.Y(n_92)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_75),
.B(n_50),
.Y(n_79)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_51),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_80),
.Y(n_109)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_81),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_85),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_58),
.B(n_50),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_94),
.B1(n_68),
.B2(n_61),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_15),
.B(n_21),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_73),
.B(n_59),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_56),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_64),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_68),
.A2(n_47),
.B1(n_43),
.B2(n_40),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_96),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_62),
.B1(n_72),
.B2(n_40),
.Y(n_115)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_102),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_68),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_110),
.Y(n_144)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_116),
.B1(n_97),
.B2(n_92),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_59),
.B(n_68),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_106),
.A2(n_112),
.B(n_97),
.Y(n_124)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_57),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_28),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_81),
.C(n_84),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_60),
.B1(n_15),
.B2(n_74),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_64),
.B1(n_46),
.B2(n_63),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_88),
.A2(n_36),
.B1(n_76),
.B2(n_17),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_120),
.A2(n_76),
.B1(n_98),
.B2(n_87),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_124),
.A2(n_143),
.B(n_27),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_126),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_106),
.B(n_108),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_130),
.B(n_141),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_97),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_127),
.B1(n_133),
.B2(n_143),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_103),
.Y(n_132)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_94),
.B1(n_31),
.B2(n_83),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_138),
.C(n_139),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_117),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_0),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_80),
.B1(n_82),
.B2(n_96),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_93),
.B1(n_31),
.B2(n_72),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_110),
.C(n_113),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_102),
.C(n_107),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_31),
.B(n_33),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_103),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_105),
.Y(n_149)
);

NOR2x1_ASAP7_75t_R g143 ( 
.A(n_116),
.B(n_33),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_78),
.B1(n_67),
.B2(n_95),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_118),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_150),
.C(n_152),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_124),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_156),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_148),
.A2(n_151),
.B1(n_153),
.B2(n_162),
.Y(n_189)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_120),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_131),
.A2(n_100),
.B1(n_111),
.B2(n_121),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_99),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_133),
.A2(n_105),
.B1(n_74),
.B2(n_67),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_103),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_168),
.Y(n_173)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_157),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_17),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_139),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_132),
.B1(n_123),
.B2(n_91),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_78),
.B1(n_27),
.B2(n_60),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_60),
.B1(n_17),
.B2(n_95),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_163),
.A2(n_128),
.B1(n_141),
.B2(n_125),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_91),
.C(n_17),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_170),
.C(n_132),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_128),
.A2(n_27),
.B1(n_17),
.B2(n_95),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_191)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_21),
.B(n_91),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_21),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_179),
.B1(n_3),
.B2(n_4),
.Y(n_210)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_153),
.A2(n_137),
.B1(n_129),
.B2(n_123),
.Y(n_175)
);

OA21x2_ASAP7_75t_L g208 ( 
.A1(n_175),
.A2(n_156),
.B(n_4),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_129),
.Y(n_176)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_181),
.Y(n_198)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_164),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_147),
.B(n_21),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_183),
.B(n_3),
.Y(n_209)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_186),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_165),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_190),
.C(n_194),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_140),
.C(n_1),
.Y(n_190)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_159),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_3),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_0),
.C(n_2),
.Y(n_194)
);

INVxp33_ASAP7_75t_SL g195 ( 
.A(n_175),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_195),
.A2(n_208),
.B(n_213),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_197),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_150),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_206),
.C(n_211),
.Y(n_215)
);

NAND3xp33_ASAP7_75t_SL g201 ( 
.A(n_175),
.B(n_169),
.C(n_170),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_201),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_205),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_171),
.B(n_161),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_161),
.Y(n_206)
);

FAx1_ASAP7_75t_SL g231 ( 
.A(n_209),
.B(n_194),
.CI(n_191),
.CON(n_231),
.SN(n_231)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_212),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_12),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_192),
.B1(n_185),
.B2(n_174),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_218),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_189),
.B(n_182),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_227),
.B(n_228),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_184),
.C(n_190),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_223),
.C(n_207),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_184),
.C(n_187),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_207),
.B(n_171),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_230),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_203),
.A2(n_188),
.B(n_173),
.Y(n_227)
);

FAx1_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_183),
.CI(n_189),
.CON(n_228),
.SN(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_173),
.B(n_172),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_229),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_208),
.B(n_202),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_231),
.B(n_211),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_12),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_231),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_233),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_237),
.C(n_240),
.Y(n_259)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_209),
.C(n_6),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_230),
.B(n_217),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_11),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_243),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_7),
.C(n_8),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_11),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_219),
.B(n_7),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_225),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_8),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_225),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_8),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_247),
.B(n_226),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_228),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_256),
.C(n_258),
.Y(n_267)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_252),
.B(n_253),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_227),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_231),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_229),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_235),
.A2(n_220),
.B(n_218),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_221),
.C(n_228),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_8),
.C(n_9),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_249),
.B(n_238),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_263),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_237),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_243),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_265),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_239),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_240),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_270),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_271),
.A2(n_259),
.B(n_248),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_267),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_272),
.A2(n_274),
.B(n_275),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g274 ( 
.A1(n_270),
.A2(n_250),
.B(n_255),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_257),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_262),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_269),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_277),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_269),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_282),
.A2(n_284),
.B(n_261),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_283),
.A2(n_278),
.B(n_280),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_273),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_285),
.A2(n_286),
.B(n_281),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_279),
.C(n_253),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_9),
.C(n_10),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_289),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_10),
.B(n_272),
.Y(n_291)
);


endmodule