module real_aes_10392_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_552;
wire n_590;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_360;
wire n_859;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_315;
wire n_1161;
wire n_686;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_837;
wire n_829;
wire n_1030;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_333;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1162;
wire n_762;
wire n_325;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1050;
wire n_426;
wire n_1134;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_714;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1033;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_644;
wire n_1150;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_974;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1198;
wire n_304;
wire n_993;
wire n_819;
wire n_737;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_269;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_338;
wire n_698;
wire n_371;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_340;
wire n_483;
wire n_1280;
wire n_729;
wire n_394;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_0), .A2(n_220), .B1(n_656), .B2(n_780), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_0), .A2(n_220), .B1(n_545), .B2(n_820), .Y(n_1270) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_1), .A2(n_13), .B1(n_378), .B2(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g419 ( .A(n_1), .Y(n_419) );
INVx1_ASAP7_75t_L g865 ( .A(n_2), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_2), .A2(n_136), .B1(n_599), .B2(n_824), .Y(n_875) );
AO221x1_ASAP7_75t_L g1044 ( .A1(n_3), .A2(n_151), .B1(n_991), .B2(n_1045), .C(n_1047), .Y(n_1044) );
INVxp67_ASAP7_75t_SL g713 ( .A(n_4), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_4), .A2(n_22), .B1(n_553), .B2(n_612), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_5), .A2(n_10), .B1(n_383), .B2(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g891 ( .A(n_5), .Y(n_891) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_6), .Y(n_262) );
INVx1_ASAP7_75t_L g372 ( .A(n_6), .Y(n_372) );
INVx1_ASAP7_75t_L g326 ( .A(n_7), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g1036 ( .A1(n_8), .A2(n_107), .B1(n_991), .B2(n_1016), .Y(n_1036) );
AOI22xp33_ASAP7_75t_SL g772 ( .A1(n_9), .A2(n_197), .B1(n_342), .B2(n_729), .Y(n_772) );
AOI22xp33_ASAP7_75t_SL g782 ( .A1(n_9), .A2(n_197), .B1(n_386), .B2(n_562), .Y(n_782) );
INVx1_ASAP7_75t_L g892 ( .A(n_10), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_11), .A2(n_39), .B1(n_624), .B2(n_626), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_11), .A2(n_39), .B1(n_629), .B2(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g518 ( .A(n_12), .Y(n_518) );
INVx1_ASAP7_75t_L g409 ( .A(n_13), .Y(n_409) );
INVx1_ASAP7_75t_L g590 ( .A(n_14), .Y(n_590) );
INVxp33_ASAP7_75t_SL g649 ( .A(n_15), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_15), .A2(n_240), .B1(n_547), .B2(n_669), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_16), .A2(n_171), .B1(n_342), .B2(n_729), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_16), .A2(n_171), .B1(n_386), .B2(n_576), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_17), .A2(n_237), .B1(n_386), .B2(n_562), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_17), .A2(n_237), .B1(n_430), .B2(n_434), .Y(n_986) );
INVx1_ASAP7_75t_L g702 ( .A(n_18), .Y(n_702) );
CKINVDCx5p33_ASAP7_75t_R g859 ( .A(n_19), .Y(n_859) );
AO221x2_ASAP7_75t_L g1067 ( .A1(n_20), .A2(n_161), .B1(n_1045), .B2(n_1068), .C(n_1070), .Y(n_1067) );
INVx1_ASAP7_75t_L g863 ( .A(n_21), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_21), .A2(n_245), .B1(n_612), .B2(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g712 ( .A(n_22), .Y(n_712) );
INVx1_ASAP7_75t_L g751 ( .A(n_23), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_23), .A2(n_120), .B1(n_718), .B2(n_774), .Y(n_777) );
INVx1_ASAP7_75t_L g1210 ( .A(n_24), .Y(n_1210) );
AOI22xp33_ASAP7_75t_L g1234 ( .A1(n_24), .A2(n_179), .B1(n_1235), .B2(n_1236), .Y(n_1234) );
INVx2_ASAP7_75t_L g284 ( .A(n_25), .Y(n_284) );
INVx1_ASAP7_75t_L g697 ( .A(n_26), .Y(n_697) );
INVxp33_ASAP7_75t_SL g529 ( .A(n_27), .Y(n_529) );
AOI22xp5_ASAP7_75t_SL g571 ( .A1(n_27), .A2(n_62), .B1(n_572), .B2(n_576), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_28), .A2(n_209), .B1(n_729), .B2(n_909), .Y(n_908) );
INVxp67_ASAP7_75t_SL g938 ( .A(n_28), .Y(n_938) );
INVx1_ASAP7_75t_L g808 ( .A(n_29), .Y(n_808) );
AOI22xp33_ASAP7_75t_SL g823 ( .A1(n_29), .A2(n_200), .B1(n_718), .B2(n_824), .Y(n_823) );
BUFx2_ASAP7_75t_L g331 ( .A(n_30), .Y(n_331) );
INVx1_ASAP7_75t_L g368 ( .A(n_30), .Y(n_368) );
BUFx2_ASAP7_75t_L g403 ( .A(n_30), .Y(n_403) );
AO22x1_ASAP7_75t_L g510 ( .A1(n_31), .A2(n_511), .B1(n_512), .B2(n_581), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_31), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_32), .A2(n_177), .B1(n_918), .B2(n_919), .Y(n_917) );
OAI211xp5_ASAP7_75t_SL g923 ( .A1(n_32), .A2(n_426), .B(n_924), .C(n_927), .Y(n_923) );
INVx1_ASAP7_75t_L g654 ( .A(n_33), .Y(n_654) );
AOI22xp33_ASAP7_75t_SL g670 ( .A1(n_33), .A2(n_68), .B1(n_346), .B2(n_671), .Y(n_670) );
AOI22xp33_ASAP7_75t_SL g1267 ( .A1(n_34), .A2(n_101), .B1(n_562), .B2(n_1268), .Y(n_1267) );
INVxp67_ASAP7_75t_L g1277 ( .A(n_34), .Y(n_1277) );
AOI22xp33_ASAP7_75t_SL g345 ( .A1(n_35), .A2(n_199), .B1(n_346), .B2(n_350), .Y(n_345) );
AOI22xp33_ASAP7_75t_SL g374 ( .A1(n_35), .A2(n_199), .B1(n_375), .B2(n_378), .Y(n_374) );
INVx1_ASAP7_75t_L g593 ( .A(n_36), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_36), .A2(n_92), .B1(n_599), .B2(n_615), .Y(n_614) );
AOI22xp33_ASAP7_75t_SL g539 ( .A1(n_37), .A2(n_163), .B1(n_540), .B2(n_543), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_37), .A2(n_163), .B1(n_567), .B2(n_570), .Y(n_566) );
INVx1_ASAP7_75t_L g595 ( .A(n_38), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_38), .A2(n_145), .B1(n_469), .B2(n_470), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_40), .A2(n_169), .B1(n_599), .B2(n_774), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_40), .A2(n_169), .B1(n_656), .B2(n_913), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_41), .A2(n_50), .B1(n_612), .B2(n_619), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_41), .A2(n_50), .B1(n_565), .B2(n_632), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_42), .A2(n_146), .B1(n_665), .B2(n_666), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_42), .A2(n_146), .B1(n_497), .B2(n_676), .Y(n_675) );
INVxp67_ASAP7_75t_L g473 ( .A(n_43), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_43), .A2(n_118), .B1(n_504), .B2(n_505), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_44), .A2(n_244), .B1(n_335), .B2(n_1218), .Y(n_1217) );
AOI22xp33_ASAP7_75t_SL g1225 ( .A1(n_44), .A2(n_244), .B1(n_1226), .B2(n_1227), .Y(n_1225) );
INVx1_ASAP7_75t_L g754 ( .A(n_45), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_45), .A2(n_226), .B1(n_342), .B2(n_549), .Y(n_776) );
OAI211xp5_ASAP7_75t_L g309 ( .A1(n_46), .A2(n_310), .B(n_313), .C(n_318), .Y(n_309) );
AOI22xp33_ASAP7_75t_SL g364 ( .A1(n_46), .A2(n_198), .B1(n_347), .B2(n_350), .Y(n_364) );
INVx1_ASAP7_75t_L g701 ( .A(n_47), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_47), .A2(n_182), .B1(n_615), .B2(n_718), .Y(n_733) );
INVx1_ASAP7_75t_L g1048 ( .A(n_48), .Y(n_1048) );
INVx1_ASAP7_75t_L g1197 ( .A(n_49), .Y(n_1197) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_49), .A2(n_143), .B1(n_547), .B2(n_669), .Y(n_1219) );
INVx1_ASAP7_75t_L g657 ( .A(n_51), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_51), .A2(n_213), .B1(n_469), .B2(n_686), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_52), .A2(n_170), .B1(n_335), .B2(n_340), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_52), .A2(n_170), .B1(n_381), .B2(n_384), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_53), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g1266 ( .A1(n_54), .A2(n_221), .B1(n_913), .B2(n_919), .Y(n_1266) );
INVxp33_ASAP7_75t_L g1279 ( .A(n_54), .Y(n_1279) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_55), .A2(n_129), .B1(n_346), .B2(n_556), .Y(n_663) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_55), .A2(n_129), .B1(n_378), .B2(n_393), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_56), .A2(n_204), .B1(n_599), .B2(n_820), .Y(n_910) );
INVx1_ASAP7_75t_L g934 ( .A(n_56), .Y(n_934) );
INVx1_ASAP7_75t_L g532 ( .A(n_57), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_57), .A2(n_138), .B1(n_567), .B2(n_579), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_58), .A2(n_82), .B1(n_280), .B2(n_295), .Y(n_948) );
INVx1_ASAP7_75t_L g965 ( .A(n_58), .Y(n_965) );
INVx1_ASAP7_75t_L g1202 ( .A(n_59), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g1220 ( .A1(n_59), .A2(n_105), .B1(n_543), .B2(n_1221), .Y(n_1220) );
INVx1_ASAP7_75t_L g453 ( .A(n_60), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_60), .A2(n_75), .B1(n_350), .B2(n_481), .Y(n_490) );
OAI22xp33_ASAP7_75t_L g954 ( .A1(n_61), .A2(n_228), .B1(n_290), .B2(n_303), .Y(n_954) );
AOI221xp5_ASAP7_75t_L g961 ( .A1(n_61), .A2(n_228), .B1(n_547), .B2(n_962), .C(n_964), .Y(n_961) );
INVxp33_ASAP7_75t_SL g530 ( .A(n_62), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_63), .A2(n_233), .B1(n_656), .B2(n_780), .Y(n_881) );
INVx1_ASAP7_75t_L g887 ( .A(n_63), .Y(n_887) );
INVx1_ASAP7_75t_L g1049 ( .A(n_64), .Y(n_1049) );
INVx1_ASAP7_75t_L g450 ( .A(n_65), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g1243 ( .A1(n_66), .A2(n_1244), .B1(n_1245), .B2(n_1280), .Y(n_1243) );
CKINVDCx5p33_ASAP7_75t_R g1244 ( .A(n_66), .Y(n_1244) );
INVxp67_ASAP7_75t_SL g606 ( .A(n_67), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_67), .A2(n_144), .B1(n_504), .B2(n_572), .Y(n_638) );
INVxp33_ASAP7_75t_SL g647 ( .A(n_68), .Y(n_647) );
AOI22xp33_ASAP7_75t_SL g818 ( .A1(n_69), .A2(n_242), .B1(n_342), .B2(n_729), .Y(n_818) );
AOI22xp33_ASAP7_75t_SL g827 ( .A1(n_69), .A2(n_242), .B1(n_383), .B2(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g769 ( .A(n_70), .Y(n_769) );
AOI22xp33_ASAP7_75t_SL g785 ( .A1(n_70), .A2(n_81), .B1(n_562), .B2(n_745), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_71), .A2(n_149), .B1(n_718), .B2(n_774), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_71), .A2(n_149), .B1(n_656), .B2(n_780), .Y(n_779) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_72), .A2(n_96), .B1(n_710), .B2(n_759), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_72), .A2(n_96), .B1(n_470), .B2(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g722 ( .A(n_73), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_73), .A2(n_93), .B1(n_562), .B2(n_745), .Y(n_744) );
AO221x1_ASAP7_75t_L g1025 ( .A1(n_74), .A2(n_113), .B1(n_991), .B2(n_1016), .C(n_1026), .Y(n_1025) );
AOI222xp33_ASAP7_75t_L g1190 ( .A1(n_74), .A2(n_1191), .B1(n_1237), .B2(n_1242), .C1(n_1281), .C2(n_1285), .Y(n_1190) );
XNOR2x2_ASAP7_75t_L g1192 ( .A(n_74), .B(n_1193), .Y(n_1192) );
INVxp33_ASAP7_75t_SL g445 ( .A(n_75), .Y(n_445) );
INVx1_ASAP7_75t_L g1073 ( .A(n_76), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_77), .A2(n_206), .B1(n_547), .B2(n_550), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_77), .A2(n_206), .B1(n_561), .B2(n_563), .Y(n_560) );
INVx1_ASAP7_75t_L g525 ( .A(n_78), .Y(n_525) );
INVxp33_ASAP7_75t_SL g588 ( .A(n_79), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_79), .A2(n_158), .B1(n_612), .B2(n_613), .Y(n_611) );
AO22x2_ASAP7_75t_L g791 ( .A1(n_80), .A2(n_792), .B1(n_834), .B2(n_835), .Y(n_791) );
INVxp67_ASAP7_75t_L g834 ( .A(n_80), .Y(n_834) );
INVx1_ASAP7_75t_L g767 ( .A(n_81), .Y(n_767) );
INVx1_ASAP7_75t_L g985 ( .A(n_82), .Y(n_985) );
AO221x1_ASAP7_75t_L g1019 ( .A1(n_83), .A2(n_156), .B1(n_991), .B2(n_1016), .C(n_1020), .Y(n_1019) );
INVx1_ASAP7_75t_L g941 ( .A(n_84), .Y(n_941) );
INVx1_ASAP7_75t_L g329 ( .A(n_85), .Y(n_329) );
INVx1_ASAP7_75t_L g929 ( .A(n_86), .Y(n_929) );
INVx1_ASAP7_75t_L g1253 ( .A(n_87), .Y(n_1253) );
OAI22xp5_ASAP7_75t_L g1274 ( .A1(n_87), .A2(n_88), .B1(n_469), .B2(n_686), .Y(n_1274) );
INVx1_ASAP7_75t_L g1254 ( .A(n_88), .Y(n_1254) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_89), .A2(n_178), .B1(n_707), .B2(n_710), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_89), .A2(n_178), .B1(n_469), .B2(n_470), .Y(n_719) );
INVx1_ASAP7_75t_L g958 ( .A(n_90), .Y(n_958) );
INVxp67_ASAP7_75t_SL g465 ( .A(n_91), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_91), .A2(n_128), .B1(n_493), .B2(n_502), .Y(n_501) );
INVxp33_ASAP7_75t_SL g587 ( .A(n_92), .Y(n_587) );
INVxp67_ASAP7_75t_L g724 ( .A(n_93), .Y(n_724) );
INVx1_ASAP7_75t_L g867 ( .A(n_94), .Y(n_867) );
OAI22xp33_ASAP7_75t_L g889 ( .A1(n_94), .A2(n_174), .B1(n_686), .B2(n_801), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_95), .A2(n_140), .B1(n_383), .B2(n_565), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_95), .A2(n_140), .B1(n_430), .B2(n_434), .Y(n_922) );
INVx1_ASAP7_75t_L g795 ( .A(n_97), .Y(n_795) );
AOI22xp33_ASAP7_75t_SL g833 ( .A1(n_97), .A2(n_208), .B1(n_562), .B2(n_745), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_98), .A2(n_192), .B1(n_466), .B2(n_820), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_98), .A2(n_192), .B1(n_456), .B2(n_502), .Y(n_826) );
INVxp33_ASAP7_75t_SL g515 ( .A(n_99), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_99), .A2(n_246), .B1(n_540), .B2(n_556), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_100), .A2(n_202), .B1(n_991), .B2(n_1016), .Y(n_1041) );
INVxp33_ASAP7_75t_L g1276 ( .A(n_101), .Y(n_1276) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_102), .A2(n_214), .B1(n_384), .B2(n_396), .Y(n_681) );
INVxp67_ASAP7_75t_SL g689 ( .A(n_102), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_103), .A2(n_217), .B1(n_342), .B2(n_729), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_103), .A2(n_217), .B1(n_565), .B2(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g1028 ( .A(n_104), .Y(n_1028) );
INVx1_ASAP7_75t_L g1196 ( .A(n_105), .Y(n_1196) );
INVx1_ASAP7_75t_L g254 ( .A(n_106), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_108), .A2(n_162), .B1(n_396), .B2(n_399), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_108), .A2(n_162), .B1(n_430), .B2(n_434), .Y(n_429) );
INVx1_ASAP7_75t_L g766 ( .A(n_109), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_109), .A2(n_190), .B1(n_456), .B2(n_780), .Y(n_784) );
AOI221xp5_ASAP7_75t_L g956 ( .A1(n_110), .A2(n_193), .B1(n_665), .B2(n_669), .C(n_957), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_110), .A2(n_193), .B1(n_562), .B2(n_745), .Y(n_975) );
INVx1_ASAP7_75t_L g953 ( .A(n_111), .Y(n_953) );
AOI22xp5_ASAP7_75t_L g1005 ( .A1(n_112), .A2(n_184), .B1(n_1006), .B2(n_1012), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_114), .A2(n_177), .B1(n_263), .B2(n_423), .Y(n_930) );
OAI22xp33_ASAP7_75t_L g940 ( .A1(n_114), .A2(n_204), .B1(n_280), .B2(n_295), .Y(n_940) );
INVx1_ASAP7_75t_L g1027 ( .A(n_115), .Y(n_1027) );
XNOR2xp5_ASAP7_75t_L g276 ( .A(n_116), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g522 ( .A(n_117), .Y(n_522) );
INVxp67_ASAP7_75t_L g474 ( .A(n_118), .Y(n_474) );
AOI22xp33_ASAP7_75t_SL g678 ( .A1(n_119), .A2(n_236), .B1(n_630), .B2(n_679), .Y(n_678) );
INVxp67_ASAP7_75t_SL g684 ( .A(n_119), .Y(n_684) );
INVx1_ASAP7_75t_L g757 ( .A(n_120), .Y(n_757) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_121), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g1015 ( .A1(n_122), .A2(n_166), .B1(n_991), .B2(n_1016), .Y(n_1015) );
AOI22xp5_ASAP7_75t_L g1042 ( .A1(n_123), .A2(n_247), .B1(n_1006), .B2(n_1012), .Y(n_1042) );
INVx1_ASAP7_75t_L g1207 ( .A(n_124), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_124), .A2(n_189), .B1(n_1230), .B2(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1256 ( .A(n_125), .Y(n_1256) );
INVxp67_ASAP7_75t_SL g459 ( .A(n_126), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_126), .A2(n_248), .B1(n_469), .B2(n_470), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g1260 ( .A1(n_127), .A2(n_134), .B1(n_745), .B2(n_1261), .Y(n_1260) );
AOI22xp33_ASAP7_75t_SL g1269 ( .A1(n_127), .A2(n_134), .B1(n_342), .B2(n_729), .Y(n_1269) );
INVxp67_ASAP7_75t_SL g462 ( .A(n_128), .Y(n_462) );
CKINVDCx14_ASAP7_75t_R g945 ( .A(n_130), .Y(n_945) );
INVx1_ASAP7_75t_L g651 ( .A(n_131), .Y(n_651) );
INVx1_ASAP7_75t_L g952 ( .A(n_132), .Y(n_952) );
INVx1_ASAP7_75t_L g1071 ( .A(n_133), .Y(n_1071) );
INVxp33_ASAP7_75t_SL g1249 ( .A(n_135), .Y(n_1249) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_135), .A2(n_150), .B1(n_545), .B2(n_774), .Y(n_1264) );
INVx1_ASAP7_75t_L g862 ( .A(n_136), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g294 ( .A1(n_137), .A2(n_223), .B1(n_295), .B2(n_303), .Y(n_294) );
INVxp33_ASAP7_75t_SL g421 ( .A(n_137), .Y(n_421) );
INVxp33_ASAP7_75t_SL g535 ( .A(n_138), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_139), .A2(n_147), .B1(n_729), .B2(n_905), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_139), .A2(n_147), .B1(n_398), .B2(n_828), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g279 ( .A1(n_141), .A2(n_198), .B1(n_280), .B2(n_290), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_141), .A2(n_223), .B1(n_335), .B2(n_361), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g1199 ( .A(n_142), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_143), .Y(n_1200) );
INVxp33_ASAP7_75t_L g604 ( .A(n_144), .Y(n_604) );
INVx1_ASAP7_75t_L g594 ( .A(n_145), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_148), .A2(n_165), .B1(n_346), .B2(n_556), .Y(n_1216) );
AOI22xp33_ASAP7_75t_SL g1229 ( .A1(n_148), .A2(n_165), .B1(n_679), .B2(n_1230), .Y(n_1229) );
INVxp67_ASAP7_75t_SL g1252 ( .A(n_150), .Y(n_1252) );
INVxp33_ASAP7_75t_SL g448 ( .A(n_152), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g486 ( .A1(n_152), .A2(n_229), .B1(n_478), .B2(n_487), .Y(n_486) );
INVxp33_ASAP7_75t_SL g1257 ( .A(n_153), .Y(n_1257) );
AOI22xp33_ASAP7_75t_SL g1263 ( .A1(n_153), .A2(n_167), .B1(n_342), .B2(n_729), .Y(n_1263) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_154), .A2(n_224), .B1(n_545), .B2(n_820), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_154), .A2(n_224), .B1(n_656), .B2(n_780), .Y(n_877) );
XNOR2xp5_ASAP7_75t_L g440 ( .A(n_155), .B(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_157), .Y(n_256) );
AND3x2_ASAP7_75t_L g995 ( .A(n_157), .B(n_254), .C(n_996), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_157), .B(n_254), .Y(n_1011) );
INVxp33_ASAP7_75t_SL g591 ( .A(n_158), .Y(n_591) );
INVxp33_ASAP7_75t_SL g608 ( .A(n_159), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_159), .A2(n_207), .B1(n_629), .B2(n_630), .Y(n_637) );
INVx2_ASAP7_75t_L g267 ( .A(n_160), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_164), .A2(n_211), .B1(n_361), .B2(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_164), .A2(n_211), .B1(n_496), .B2(n_497), .Y(n_495) );
INVxp33_ASAP7_75t_SL g1250 ( .A(n_167), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_168), .A2(n_175), .B1(n_481), .B2(n_483), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_168), .A2(n_175), .B1(n_375), .B2(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g996 ( .A(n_172), .Y(n_996) );
INVx1_ASAP7_75t_L g1203 ( .A(n_173), .Y(n_1203) );
OAI22xp5_ASAP7_75t_L g1208 ( .A1(n_173), .A2(n_201), .B1(n_469), .B2(n_470), .Y(n_1208) );
INVx1_ASAP7_75t_L g866 ( .A(n_174), .Y(n_866) );
INVx1_ASAP7_75t_L g814 ( .A(n_176), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_176), .A2(n_216), .B1(n_550), .B2(n_612), .Y(n_822) );
INVx1_ASAP7_75t_L g1211 ( .A(n_179), .Y(n_1211) );
CKINVDCx5p33_ASAP7_75t_R g752 ( .A(n_180), .Y(n_752) );
INVx1_ASAP7_75t_L g978 ( .A(n_181), .Y(n_978) );
INVx1_ASAP7_75t_L g705 ( .A(n_182), .Y(n_705) );
INVx1_ASAP7_75t_L g269 ( .A(n_183), .Y(n_269) );
INVx2_ASAP7_75t_L g371 ( .A(n_183), .Y(n_371) );
XOR2x2_ASAP7_75t_L g643 ( .A(n_184), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g716 ( .A(n_185), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_185), .A2(n_234), .B1(n_456), .B2(n_502), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_186), .A2(n_215), .B1(n_466), .B2(n_615), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_186), .A2(n_215), .B1(n_738), .B2(n_739), .Y(n_737) );
XNOR2xp5_ASAP7_75t_L g747 ( .A(n_187), .B(n_748), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g1035 ( .A1(n_187), .A2(n_203), .B1(n_1006), .B2(n_1012), .Y(n_1035) );
OAI211xp5_ASAP7_75t_L g949 ( .A1(n_188), .A2(n_313), .B(n_950), .C(n_951), .Y(n_949) );
INVx1_ASAP7_75t_L g968 ( .A(n_188), .Y(n_968) );
INVx1_ASAP7_75t_L g1213 ( .A(n_189), .Y(n_1213) );
INVx1_ASAP7_75t_L g762 ( .A(n_190), .Y(n_762) );
INVx1_ASAP7_75t_L g798 ( .A(n_191), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_191), .A2(n_241), .B1(n_739), .B2(n_832), .Y(n_831) );
OAI211xp5_ASAP7_75t_L g838 ( .A1(n_191), .A2(n_426), .B(n_839), .C(n_844), .Y(n_838) );
INVx1_ASAP7_75t_L g1021 ( .A(n_194), .Y(n_1021) );
XNOR2xp5_ASAP7_75t_L g855 ( .A(n_195), .B(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g960 ( .A(n_196), .Y(n_960) );
INVx1_ASAP7_75t_L g812 ( .A(n_200), .Y(n_812) );
OAI211xp5_ASAP7_75t_L g849 ( .A1(n_200), .A2(n_313), .B(n_850), .C(n_852), .Y(n_849) );
INVx1_ASAP7_75t_L g1204 ( .A(n_201), .Y(n_1204) );
INVxp33_ASAP7_75t_SL g519 ( .A(n_205), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_205), .A2(n_225), .B1(n_547), .B2(n_553), .Y(n_552) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_207), .Y(n_601) );
INVx1_ASAP7_75t_L g796 ( .A(n_208), .Y(n_796) );
INVx1_ASAP7_75t_L g939 ( .A(n_209), .Y(n_939) );
INVx1_ASAP7_75t_L g323 ( .A(n_210), .Y(n_323) );
XOR2x2_ASAP7_75t_L g583 ( .A(n_212), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g659 ( .A(n_213), .Y(n_659) );
INVxp33_ASAP7_75t_SL g688 ( .A(n_214), .Y(n_688) );
INVx1_ASAP7_75t_L g809 ( .A(n_216), .Y(n_809) );
INVx1_ASAP7_75t_L g928 ( .A(n_218), .Y(n_928) );
INVx1_ASAP7_75t_L g994 ( .A(n_219), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_219), .B(n_1009), .Y(n_1014) );
INVxp67_ASAP7_75t_SL g1273 ( .A(n_221), .Y(n_1273) );
CKINVDCx5p33_ASAP7_75t_R g802 ( .A(n_222), .Y(n_802) );
INVxp33_ASAP7_75t_SL g516 ( .A(n_225), .Y(n_516) );
INVx1_ASAP7_75t_L g755 ( .A(n_226), .Y(n_755) );
AO22x1_ASAP7_75t_L g1061 ( .A1(n_227), .A2(n_232), .B1(n_1016), .B2(n_1062), .Y(n_1061) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_229), .Y(n_451) );
INVx2_ASAP7_75t_L g266 ( .A(n_230), .Y(n_266) );
AO22x1_ASAP7_75t_L g1063 ( .A1(n_231), .A2(n_235), .B1(n_1006), .B2(n_1012), .Y(n_1063) );
INVx1_ASAP7_75t_L g894 ( .A(n_233), .Y(n_894) );
INVxp33_ASAP7_75t_L g721 ( .A(n_234), .Y(n_721) );
INVxp33_ASAP7_75t_SL g691 ( .A(n_236), .Y(n_691) );
INVx1_ASAP7_75t_L g287 ( .A(n_238), .Y(n_287) );
BUFx3_ASAP7_75t_L g293 ( .A(n_238), .Y(n_293) );
INVx1_ASAP7_75t_L g289 ( .A(n_239), .Y(n_289) );
BUFx3_ASAP7_75t_L g302 ( .A(n_239), .Y(n_302) );
INVxp67_ASAP7_75t_SL g652 ( .A(n_240), .Y(n_652) );
INVx1_ASAP7_75t_L g804 ( .A(n_241), .Y(n_804) );
INVx1_ASAP7_75t_L g979 ( .A(n_243), .Y(n_979) );
INVx1_ASAP7_75t_L g860 ( .A(n_245), .Y(n_860) );
INVx1_ASAP7_75t_L g521 ( .A(n_246), .Y(n_521) );
INVxp67_ASAP7_75t_SL g457 ( .A(n_248), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_270), .B(n_988), .Y(n_249) );
BUFx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_252), .B(n_257), .Y(n_251) );
AND2x4_ASAP7_75t_L g1241 ( .A(n_252), .B(n_258), .Y(n_1241) );
NOR2xp33_ASAP7_75t_SL g252 ( .A(n_253), .B(n_255), .Y(n_252) );
INVx1_ASAP7_75t_SL g1284 ( .A(n_253), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_253), .B(n_255), .Y(n_1289) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_255), .B(n_1284), .Y(n_1283) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_263), .Y(n_258) );
INVxp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OR2x6_ASAP7_75t_L g439 ( .A(n_260), .B(n_403), .Y(n_439) );
OR2x2_ASAP7_75t_L g725 ( .A(n_260), .B(n_403), .Y(n_725) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g358 ( .A(n_261), .B(n_269), .Y(n_358) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx8_ASAP7_75t_L g420 ( .A(n_263), .Y(n_420) );
OR2x6_ASAP7_75t_L g263 ( .A(n_264), .B(n_268), .Y(n_263) );
OR2x6_ASAP7_75t_L g423 ( .A(n_264), .B(n_424), .Y(n_423) );
HB1xp67_ASAP7_75t_L g959 ( .A(n_264), .Y(n_959) );
INVx2_ASAP7_75t_SL g967 ( .A(n_264), .Y(n_967) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_L g337 ( .A(n_266), .Y(n_337) );
AND2x4_ASAP7_75t_L g343 ( .A(n_266), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g349 ( .A(n_266), .B(n_267), .Y(n_349) );
INVx1_ASAP7_75t_L g354 ( .A(n_266), .Y(n_354) );
INVx1_ASAP7_75t_L g415 ( .A(n_266), .Y(n_415) );
INVx1_ASAP7_75t_L g339 ( .A(n_267), .Y(n_339) );
INVx2_ASAP7_75t_L g344 ( .A(n_267), .Y(n_344) );
INVx1_ASAP7_75t_L g411 ( .A(n_267), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_267), .B(n_337), .Y(n_433) );
INVx1_ASAP7_75t_L g843 ( .A(n_267), .Y(n_843) );
AND2x4_ASAP7_75t_L g410 ( .A(n_268), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g470 ( .A(n_269), .B(n_414), .Y(n_470) );
OR2x2_ASAP7_75t_L g686 ( .A(n_269), .B(n_414), .Y(n_686) );
OAI22xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B1(n_786), .B2(n_787), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B1(n_640), .B2(n_641), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
XNOR2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_508), .Y(n_274) );
XOR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_440), .Y(n_275) );
NAND3x1_ASAP7_75t_L g277 ( .A(n_278), .B(n_332), .C(n_406), .Y(n_277) );
OAI31xp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_294), .A3(n_309), .B(n_327), .Y(n_278) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_285), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x6_ASAP7_75t_L g291 ( .A(n_282), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g315 ( .A(n_282), .Y(n_315) );
AND2x2_ASAP7_75t_L g704 ( .A(n_282), .B(n_656), .Y(n_704) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x6_ASAP7_75t_L g324 ( .A(n_283), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_284), .Y(n_298) );
INVx1_ASAP7_75t_L g306 ( .A(n_284), .Y(n_306) );
AND2x2_ASAP7_75t_L g390 ( .A(n_284), .B(n_329), .Y(n_390) );
INVx2_ASAP7_75t_L g405 ( .A(n_284), .Y(n_405) );
INVx2_ASAP7_75t_L g972 ( .A(n_285), .Y(n_972) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
AND2x2_ASAP7_75t_L g312 ( .A(n_286), .B(n_288), .Y(n_312) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g308 ( .A(n_287), .B(n_302), .Y(n_308) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_L g292 ( .A(n_289), .B(n_293), .Y(n_292) );
CKINVDCx6p67_ASAP7_75t_R g290 ( .A(n_291), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_291), .A2(n_445), .B1(n_446), .B2(n_448), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_291), .A2(n_446), .B1(n_515), .B2(n_516), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_291), .A2(n_446), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_291), .A2(n_647), .B1(n_648), .B2(n_649), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_291), .A2(n_304), .B1(n_712), .B2(n_713), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_291), .A2(n_304), .B1(n_754), .B2(n_755), .Y(n_753) );
AOI22xp5_ASAP7_75t_SL g807 ( .A1(n_291), .A2(n_648), .B1(n_808), .B2(n_809), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g861 ( .A1(n_291), .A2(n_446), .B1(n_862), .B2(n_863), .Y(n_861) );
AOI22xp5_ASAP7_75t_L g937 ( .A1(n_291), .A2(n_304), .B1(n_938), .B2(n_939), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_291), .A2(n_648), .B1(n_1196), .B2(n_1197), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_291), .A2(n_446), .B1(n_1249), .B2(n_1250), .Y(n_1248) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_292), .Y(n_383) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_292), .Y(n_398) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_292), .Y(n_496) );
BUFx3_ASAP7_75t_L g562 ( .A(n_292), .Y(n_562) );
INVx2_ASAP7_75t_SL g577 ( .A(n_292), .Y(n_577) );
BUFx2_ASAP7_75t_L g632 ( .A(n_292), .Y(n_632) );
BUFx6f_ASAP7_75t_L g1261 ( .A(n_292), .Y(n_1261) );
INVx2_ASAP7_75t_L g300 ( .A(n_293), .Y(n_300) );
AND2x2_ASAP7_75t_L g317 ( .A(n_293), .B(n_302), .Y(n_317) );
INVx4_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_296), .A2(n_304), .B1(n_450), .B2(n_451), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_296), .A2(n_304), .B1(n_518), .B2(n_519), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_296), .A2(n_304), .B1(n_590), .B2(n_591), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_296), .A2(n_304), .B1(n_651), .B2(n_652), .Y(n_650) );
AOI22xp5_ASAP7_75t_SL g700 ( .A1(n_296), .A2(n_446), .B1(n_701), .B2(n_702), .Y(n_700) );
AOI22xp5_ASAP7_75t_SL g750 ( .A1(n_296), .A2(n_648), .B1(n_751), .B2(n_752), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_296), .A2(n_304), .B1(n_805), .B2(n_814), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_296), .A2(n_304), .B1(n_859), .B2(n_860), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_296), .A2(n_304), .B1(n_1199), .B2(n_1200), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_296), .A2(n_304), .B1(n_1256), .B2(n_1257), .Y(n_1255) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
AND2x4_ASAP7_75t_L g319 ( .A(n_297), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_SL g458 ( .A(n_297), .B(n_320), .Y(n_458) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx6_ASAP7_75t_L g377 ( .A(n_299), .Y(n_377) );
BUFx2_ASAP7_75t_L g502 ( .A(n_299), .Y(n_502) );
INVx2_ASAP7_75t_L g781 ( .A(n_299), .Y(n_781) );
AND2x4_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g325 ( .A(n_300), .Y(n_325) );
INVx1_ASAP7_75t_L g322 ( .A(n_301), .Y(n_322) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx4_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x6_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
AND2x4_ASAP7_75t_L g446 ( .A(n_305), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g648 ( .A(n_305), .B(n_447), .Y(n_648) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g708 ( .A(n_306), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g506 ( .A(n_307), .Y(n_506) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_307), .Y(n_565) );
BUFx6f_ASAP7_75t_L g745 ( .A(n_307), .Y(n_745) );
INVx1_ASAP7_75t_L g884 ( .A(n_307), .Y(n_884) );
INVx2_ASAP7_75t_L g1228 ( .A(n_307), .Y(n_1228) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_308), .Y(n_386) );
INVx1_ASAP7_75t_L g400 ( .A(n_308), .Y(n_400) );
INVx2_ASAP7_75t_L g575 ( .A(n_308), .Y(n_575) );
INVx1_ASAP7_75t_L g829 ( .A(n_308), .Y(n_829) );
INVx2_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g851 ( .A(n_312), .Y(n_851) );
INVx2_ASAP7_75t_L g974 ( .A(n_312), .Y(n_974) );
NAND4xp25_ASAP7_75t_SL g443 ( .A(n_313), .B(n_444), .C(n_449), .D(n_452), .Y(n_443) );
NAND4xp25_ASAP7_75t_L g585 ( .A(n_313), .B(n_586), .C(n_589), .D(n_592), .Y(n_585) );
NAND3xp33_ASAP7_75t_SL g932 ( .A(n_313), .B(n_933), .C(n_937), .Y(n_932) );
NAND4xp25_ASAP7_75t_L g1247 ( .A(n_313), .B(n_1248), .C(n_1251), .D(n_1255), .Y(n_1247) );
CKINVDCx8_ASAP7_75t_R g313 ( .A(n_314), .Y(n_313) );
INVx5_ASAP7_75t_L g526 ( .A(n_314), .Y(n_526) );
AND2x4_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_316), .Y(n_494) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_316), .Y(n_656) );
INVx1_ASAP7_75t_L g740 ( .A(n_316), .Y(n_740) );
INVx2_ASAP7_75t_L g920 ( .A(n_316), .Y(n_920) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_317), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g318 ( .A1(n_319), .A2(n_323), .B1(n_324), .B2(n_326), .Y(n_318) );
INVx1_ASAP7_75t_L g524 ( .A(n_319), .Y(n_524) );
BUFx4f_ASAP7_75t_L g658 ( .A(n_319), .Y(n_658) );
AOI22xp33_ASAP7_75t_SL g852 ( .A1(n_319), .A2(n_324), .B1(n_799), .B2(n_802), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_319), .A2(n_324), .B1(n_952), .B2(n_953), .Y(n_951) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g709 ( .A(n_321), .Y(n_709) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AOI222xp33_ASAP7_75t_L g408 ( .A1(n_323), .A2(n_326), .B1(n_352), .B2(n_409), .C1(n_410), .C2(n_412), .Y(n_408) );
AOI222xp33_ASAP7_75t_L g452 ( .A1(n_324), .A2(n_453), .B1(n_454), .B2(n_457), .C1(n_458), .C2(n_459), .Y(n_452) );
AOI222xp33_ASAP7_75t_L g520 ( .A1(n_324), .A2(n_378), .B1(n_521), .B2(n_522), .C1(n_523), .C2(n_525), .Y(n_520) );
AOI222xp33_ASAP7_75t_L g592 ( .A1(n_324), .A2(n_458), .B1(n_493), .B2(n_593), .C1(n_594), .C2(n_595), .Y(n_592) );
AOI222xp33_ASAP7_75t_L g653 ( .A1(n_324), .A2(n_654), .B1(n_655), .B2(n_657), .C1(n_658), .C2(n_659), .Y(n_653) );
INVx3_ASAP7_75t_L g710 ( .A(n_324), .Y(n_710) );
AOI222xp33_ASAP7_75t_L g810 ( .A1(n_324), .A2(n_658), .B1(n_799), .B2(n_802), .C1(n_811), .C2(n_812), .Y(n_810) );
AOI222xp33_ASAP7_75t_L g864 ( .A1(n_324), .A2(n_378), .B1(n_458), .B2(n_865), .C1(n_866), .C2(n_867), .Y(n_864) );
AOI222xp33_ASAP7_75t_L g933 ( .A1(n_324), .A2(n_708), .B1(n_928), .B2(n_929), .C1(n_934), .C2(n_935), .Y(n_933) );
AOI222xp33_ASAP7_75t_L g1201 ( .A1(n_324), .A2(n_523), .B1(n_630), .B2(n_1202), .C1(n_1203), .C2(n_1204), .Y(n_1201) );
AOI222xp33_ASAP7_75t_L g1251 ( .A1(n_324), .A2(n_458), .B1(n_579), .B2(n_1252), .C1(n_1253), .C2(n_1254), .Y(n_1251) );
AOI211xp5_ASAP7_75t_L g698 ( .A1(n_327), .A2(n_699), .B(n_714), .C(n_726), .Y(n_698) );
AOI211xp5_ASAP7_75t_L g748 ( .A1(n_327), .A2(n_749), .B(n_760), .C(n_770), .Y(n_748) );
AOI211xp5_ASAP7_75t_L g856 ( .A1(n_327), .A2(n_857), .B(n_868), .C(n_885), .Y(n_856) );
OAI21xp5_ASAP7_75t_SL g931 ( .A1(n_327), .A2(n_932), .B(n_940), .Y(n_931) );
OAI31xp33_ASAP7_75t_L g947 ( .A1(n_327), .A2(n_948), .A3(n_949), .B(n_954), .Y(n_947) );
AOI211x1_ASAP7_75t_L g1246 ( .A1(n_327), .A2(n_1247), .B(n_1258), .C(n_1271), .Y(n_1246) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
AND2x4_ASAP7_75t_L g442 ( .A(n_328), .B(n_330), .Y(n_442) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g404 ( .A(n_329), .B(n_405), .Y(n_404) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g357 ( .A(n_331), .Y(n_357) );
AND4x1_ASAP7_75t_L g332 ( .A(n_333), .B(n_359), .C(n_373), .D(n_391), .Y(n_332) );
NAND3xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_345), .C(n_355), .Y(n_333) );
BUFx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x4_ASAP7_75t_L g472 ( .A(n_336), .B(n_424), .Y(n_472) );
INVx1_ASAP7_75t_L g479 ( .A(n_336), .Y(n_479) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_336), .Y(n_549) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_336), .Y(n_612) );
BUFx2_ASAP7_75t_L g665 ( .A(n_336), .Y(n_665) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_336), .Y(n_729) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_SL g1218 ( .A(n_341), .Y(n_1218) );
INVx4_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_SL g667 ( .A(n_342), .Y(n_667) );
BUFx3_ASAP7_75t_L g669 ( .A(n_342), .Y(n_669) );
INVx2_ASAP7_75t_SL g963 ( .A(n_342), .Y(n_963) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx3_ASAP7_75t_L g363 ( .A(n_343), .Y(n_363) );
INVx1_ASAP7_75t_L g437 ( .A(n_343), .Y(n_437) );
INVx1_ASAP7_75t_L g622 ( .A(n_343), .Y(n_622) );
AND2x4_ASAP7_75t_L g353 ( .A(n_344), .B(n_354), .Y(n_353) );
BUFx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_SL g482 ( .A(n_348), .Y(n_482) );
INVx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_349), .Y(n_542) );
AOI222xp33_ASAP7_75t_L g531 ( .A1(n_350), .A2(n_410), .B1(n_522), .B2(n_525), .C1(n_532), .C2(n_533), .Y(n_531) );
AOI211xp5_ASAP7_75t_L g761 ( .A1(n_350), .A2(n_427), .B(n_762), .C(n_763), .Y(n_761) );
AOI211xp5_ASAP7_75t_L g1206 ( .A1(n_350), .A2(n_427), .B(n_1207), .C(n_1208), .Y(n_1206) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g626 ( .A(n_351), .Y(n_626) );
INVx2_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
BUFx2_ASAP7_75t_L g483 ( .A(n_352), .Y(n_483) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g427 ( .A(n_353), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g467 ( .A(n_353), .Y(n_467) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_353), .Y(n_545) );
BUFx3_ASAP7_75t_L g600 ( .A(n_353), .Y(n_600) );
BUFx2_ASAP7_75t_L g673 ( .A(n_353), .Y(n_673) );
BUFx3_ASAP7_75t_L g718 ( .A(n_353), .Y(n_718) );
BUFx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AOI33xp33_ASAP7_75t_L g662 ( .A1(n_356), .A2(n_557), .A3(n_663), .B1(n_664), .B2(n_668), .B3(n_670), .Y(n_662) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
OR2x2_ASAP7_75t_L g388 ( .A(n_357), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g484 ( .A(n_357), .B(n_358), .Y(n_484) );
OR2x6_ASAP7_75t_L g499 ( .A(n_357), .B(n_389), .Y(n_499) );
OR2x2_ASAP7_75t_L g634 ( .A(n_357), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g734 ( .A(n_357), .B(n_735), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_364), .C(n_365), .Y(n_359) );
BUFx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx3_ASAP7_75t_L g489 ( .A(n_363), .Y(n_489) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_363), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g485 ( .A(n_365), .B(n_486), .C(n_490), .Y(n_485) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_365), .B(n_611), .C(n_614), .Y(n_610) );
INVx5_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx6_ASAP7_75t_L g557 ( .A(n_366), .Y(n_557) );
OR2x6_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g735 ( .A(n_369), .Y(n_735) );
NAND2x1p5_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
INVx1_ASAP7_75t_L g417 ( .A(n_370), .Y(n_417) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g425 ( .A(n_371), .Y(n_425) );
NAND3xp33_ASAP7_75t_L g373 ( .A(n_374), .B(n_380), .C(n_387), .Y(n_373) );
INVx4_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g629 ( .A(n_376), .Y(n_629) );
INVx1_ASAP7_75t_L g832 ( .A(n_376), .Y(n_832) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_377), .Y(n_394) );
INVx2_ASAP7_75t_L g447 ( .A(n_377), .Y(n_447) );
INVx2_ASAP7_75t_L g569 ( .A(n_377), .Y(n_569) );
INVx2_ASAP7_75t_L g680 ( .A(n_377), .Y(n_680) );
INVx1_ASAP7_75t_L g738 ( .A(n_377), .Y(n_738) );
INVx1_ASAP7_75t_L g918 ( .A(n_377), .Y(n_918) );
BUFx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_379), .Y(n_456) );
INVx1_ASAP7_75t_L g580 ( .A(n_379), .Y(n_580) );
BUFx4f_ASAP7_75t_L g630 ( .A(n_379), .Y(n_630) );
INVx1_ASAP7_75t_L g936 ( .A(n_379), .Y(n_936) );
INVx2_ASAP7_75t_SL g1231 ( .A(n_379), .Y(n_1231) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx3_ASAP7_75t_L g1226 ( .A(n_383), .Y(n_1226) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_386), .Y(n_497) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
OAI22xp5_ASAP7_75t_SL g969 ( .A1(n_388), .A2(n_970), .B1(n_976), .B2(n_977), .Y(n_969) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g635 ( .A(n_390), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_395), .C(n_401), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g676 ( .A(n_397), .Y(n_676) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g1236 ( .A(n_400), .Y(n_1236) );
AOI33xp33_ASAP7_75t_L g674 ( .A1(n_401), .A2(n_559), .A3(n_675), .B1(n_677), .B2(n_678), .B3(n_681), .Y(n_674) );
AOI33xp33_ASAP7_75t_L g1223 ( .A1(n_401), .A2(n_1224), .A3(n_1225), .B1(n_1229), .B2(n_1232), .B3(n_1234), .Y(n_1223) );
BUFx4f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx4f_ASAP7_75t_L g507 ( .A(n_402), .Y(n_507) );
AOI33xp33_ASAP7_75t_L g558 ( .A1(n_402), .A2(n_559), .A3(n_560), .B1(n_566), .B2(n_571), .B3(n_578), .Y(n_558) );
INVx4_ASAP7_75t_L g976 ( .A(n_402), .Y(n_976) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
AND2x4_ASAP7_75t_L g639 ( .A(n_403), .B(n_404), .Y(n_639) );
OAI21xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_429), .B(n_438), .Y(n_406) );
NAND3xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_418), .C(n_426), .Y(n_407) );
INVx2_ASAP7_75t_L g469 ( .A(n_410), .Y(n_469) );
INVx2_ASAP7_75t_L g764 ( .A(n_410), .Y(n_764) );
INVx2_ASAP7_75t_L g801 ( .A(n_410), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_410), .A2(n_533), .B1(n_928), .B2(n_929), .Y(n_927) );
AOI222xp33_ASAP7_75t_L g983 ( .A1(n_410), .A2(n_533), .B1(n_717), .B2(n_952), .C1(n_953), .C2(n_979), .Y(n_983) );
AOI222xp33_ASAP7_75t_L g797 ( .A1(n_412), .A2(n_599), .B1(n_798), .B2(n_799), .C1(n_800), .C2(n_802), .Y(n_797) );
AND2x4_ASAP7_75t_L g412 ( .A(n_413), .B(n_416), .Y(n_412) );
AND2x4_ASAP7_75t_L g533 ( .A(n_413), .B(n_416), .Y(n_533) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g842 ( .A(n_415), .B(n_843), .Y(n_842) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g428 ( .A(n_417), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B1(n_421), .B2(n_422), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_420), .A2(n_450), .B1(n_462), .B2(n_463), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_420), .A2(n_463), .B1(n_518), .B2(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_420), .A2(n_463), .B1(n_590), .B2(n_608), .Y(n_607) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_420), .A2(n_422), .B1(n_651), .B2(n_691), .Y(n_690) );
AOI22xp33_ASAP7_75t_SL g720 ( .A1(n_420), .A2(n_472), .B1(n_721), .B2(n_722), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_420), .A2(n_472), .B1(n_766), .B2(n_767), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_420), .A2(n_422), .B1(n_804), .B2(n_805), .Y(n_803) );
AOI22xp33_ASAP7_75t_SL g893 ( .A1(n_420), .A2(n_422), .B1(n_859), .B2(n_894), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_420), .A2(n_422), .B1(n_978), .B2(n_985), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g1212 ( .A1(n_420), .A2(n_422), .B1(n_1199), .B2(n_1213), .Y(n_1212) );
AOI22xp33_ASAP7_75t_SL g1278 ( .A1(n_420), .A2(n_463), .B1(n_1256), .B2(n_1279), .Y(n_1278) );
INVx4_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx5_ASAP7_75t_L g463 ( .A(n_423), .Y(n_463) );
INVx1_ASAP7_75t_L g431 ( .A(n_424), .Y(n_431) );
AND2x4_ASAP7_75t_L g435 ( .A(n_424), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g605 ( .A(n_424), .B(n_436), .Y(n_605) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND4xp25_ASAP7_75t_SL g527 ( .A(n_426), .B(n_528), .C(n_531), .D(n_534), .Y(n_527) );
NAND4xp25_ASAP7_75t_L g793 ( .A(n_426), .B(n_794), .C(n_797), .D(n_803), .Y(n_793) );
NAND3xp33_ASAP7_75t_L g982 ( .A(n_426), .B(n_983), .C(n_984), .Y(n_982) );
CKINVDCx11_ASAP7_75t_R g426 ( .A(n_427), .Y(n_426) );
AOI211xp5_ASAP7_75t_L g464 ( .A1(n_427), .A2(n_465), .B(n_466), .C(n_468), .Y(n_464) );
AOI211xp5_ASAP7_75t_L g597 ( .A1(n_427), .A2(n_598), .B(n_601), .C(n_602), .Y(n_597) );
AOI211xp5_ASAP7_75t_SL g683 ( .A1(n_427), .A2(n_466), .B(n_684), .C(n_685), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g715 ( .A1(n_427), .A2(n_716), .B(n_717), .C(n_719), .Y(n_715) );
AOI211xp5_ASAP7_75t_L g886 ( .A1(n_427), .A2(n_887), .B(n_888), .C(n_889), .Y(n_886) );
AOI211xp5_ASAP7_75t_L g1272 ( .A1(n_427), .A2(n_888), .B(n_1273), .C(n_1274), .Y(n_1272) );
OR2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
BUFx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx5_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
AOI22xp5_ASAP7_75t_SL g471 ( .A1(n_435), .A2(n_472), .B1(n_473), .B2(n_474), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_435), .A2(n_472), .B1(n_529), .B2(n_530), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_435), .A2(n_472), .B1(n_688), .B2(n_689), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_435), .A2(n_463), .B1(n_702), .B2(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_435), .A2(n_463), .B1(n_752), .B2(n_769), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_435), .A2(n_472), .B1(n_795), .B2(n_796), .Y(n_794) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_437), .Y(n_554) );
AOI221xp5_ASAP7_75t_L g512 ( .A1(n_438), .A2(n_442), .B1(n_513), .B2(n_527), .C(n_536), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g584 ( .A1(n_438), .A2(n_442), .B1(n_585), .B2(n_596), .C(n_609), .Y(n_584) );
AOI221x1_ASAP7_75t_L g792 ( .A1(n_438), .A2(n_660), .B1(n_793), .B2(n_806), .C(n_815), .Y(n_792) );
OAI31xp33_ASAP7_75t_L g836 ( .A1(n_438), .A2(n_837), .A3(n_838), .B(n_846), .Y(n_836) );
OAI31xp33_ASAP7_75t_SL g921 ( .A1(n_438), .A2(n_922), .A3(n_923), .B(n_930), .Y(n_921) );
OAI21xp5_ASAP7_75t_L g981 ( .A1(n_438), .A2(n_982), .B(n_986), .Y(n_981) );
CKINVDCx16_ASAP7_75t_R g438 ( .A(n_439), .Y(n_438) );
AOI31xp33_ASAP7_75t_L g460 ( .A1(n_439), .A2(n_461), .A3(n_464), .B(n_471), .Y(n_460) );
AOI31xp33_ASAP7_75t_L g682 ( .A1(n_439), .A2(n_683), .A3(n_687), .B(n_690), .Y(n_682) );
AOI31xp33_ASAP7_75t_L g885 ( .A1(n_439), .A2(n_886), .A3(n_890), .B(n_893), .Y(n_885) );
AOI31xp33_ASAP7_75t_L g1205 ( .A1(n_439), .A2(n_1206), .A3(n_1209), .B(n_1212), .Y(n_1205) );
AO211x2_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_443), .B(n_460), .C(n_475), .Y(n_441) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_442), .Y(n_660) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g570 ( .A(n_455), .Y(n_570) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_472), .A2(n_604), .B1(n_605), .B2(n_606), .Y(n_603) );
AOI22xp33_ASAP7_75t_SL g890 ( .A1(n_472), .A2(n_605), .B1(n_891), .B2(n_892), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_472), .A2(n_605), .B1(n_1210), .B2(n_1211), .Y(n_1209) );
AOI22xp33_ASAP7_75t_SL g1275 ( .A1(n_472), .A2(n_605), .B1(n_1276), .B2(n_1277), .Y(n_1275) );
NAND4xp25_ASAP7_75t_L g475 ( .A(n_476), .B(n_485), .C(n_491), .D(n_500), .Y(n_475) );
NAND3xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_480), .C(n_484), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g625 ( .A(n_482), .Y(n_625) );
BUFx3_ASAP7_75t_L g538 ( .A(n_484), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g617 ( .A(n_484), .B(n_618), .C(n_623), .Y(n_617) );
NAND3xp33_ASAP7_75t_L g727 ( .A(n_484), .B(n_728), .C(n_730), .Y(n_727) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_484), .B(n_772), .C(n_773), .Y(n_771) );
NAND3xp33_ASAP7_75t_L g817 ( .A(n_484), .B(n_818), .C(n_819), .Y(n_817) );
NAND3xp33_ASAP7_75t_L g869 ( .A(n_484), .B(n_870), .C(n_871), .Y(n_869) );
NAND3xp33_ASAP7_75t_L g903 ( .A(n_484), .B(n_904), .C(n_906), .Y(n_903) );
AOI33xp33_ASAP7_75t_L g1265 ( .A1(n_484), .A2(n_639), .A3(n_1266), .B1(n_1267), .B2(n_1269), .B3(n_1270), .Y(n_1265) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_495), .C(n_498), .Y(n_491) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx4f_ASAP7_75t_L g504 ( .A(n_496), .Y(n_504) );
BUFx2_ASAP7_75t_L g1235 ( .A(n_496), .Y(n_1235) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_499), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g1224 ( .A(n_499), .Y(n_1224) );
NAND3xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .C(n_507), .Y(n_500) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B1(n_582), .B2(n_583), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g581 ( .A(n_512), .Y(n_581) );
NAND4xp25_ASAP7_75t_L g513 ( .A(n_514), .B(n_517), .C(n_520), .D(n_526), .Y(n_513) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND4xp25_ASAP7_75t_SL g645 ( .A(n_526), .B(n_646), .C(n_650), .D(n_653), .Y(n_645) );
NAND4xp25_ASAP7_75t_L g699 ( .A(n_526), .B(n_700), .C(n_703), .D(n_711), .Y(n_699) );
NAND4xp25_ASAP7_75t_L g749 ( .A(n_526), .B(n_750), .C(n_753), .D(n_756), .Y(n_749) );
NAND4xp25_ASAP7_75t_L g806 ( .A(n_526), .B(n_807), .C(n_810), .D(n_813), .Y(n_806) );
NAND4xp25_ASAP7_75t_L g857 ( .A(n_526), .B(n_858), .C(n_861), .D(n_864), .Y(n_857) );
NAND4xp25_ASAP7_75t_SL g1194 ( .A(n_526), .B(n_1195), .C(n_1198), .D(n_1201), .Y(n_1194) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_533), .A2(n_799), .B1(n_802), .B2(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_558), .Y(n_536) );
AOI33xp33_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_539), .A3(n_546), .B1(n_552), .B2(n_555), .B3(n_557), .Y(n_537) );
AOI221xp5_ASAP7_75t_L g955 ( .A1(n_538), .A2(n_557), .B1(n_956), .B2(n_961), .C(n_969), .Y(n_955) );
AOI33xp33_ASAP7_75t_L g1215 ( .A1(n_538), .A2(n_557), .A3(n_1216), .B1(n_1217), .B2(n_1219), .B3(n_1220), .Y(n_1215) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g1222 ( .A(n_541), .Y(n_1222) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx3_ASAP7_75t_L g616 ( .A(n_542), .Y(n_616) );
BUFx2_ASAP7_75t_L g824 ( .A(n_542), .Y(n_824) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_SL g556 ( .A(n_544), .Y(n_556) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
BUFx6f_ASAP7_75t_L g888 ( .A(n_545), .Y(n_888) );
INVx3_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
INVx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g613 ( .A(n_551), .Y(n_613) );
INVx2_ASAP7_75t_SL g874 ( .A(n_551), .Y(n_874) );
INVx2_ASAP7_75t_L g905 ( .A(n_551), .Y(n_905) );
INVx2_ASAP7_75t_L g909 ( .A(n_551), .Y(n_909) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND3xp33_ASAP7_75t_L g907 ( .A(n_557), .B(n_908), .C(n_910), .Y(n_907) );
BUFx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
BUFx2_ASAP7_75t_L g1268 ( .A(n_574), .Y(n_1268) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g879 ( .A(n_577), .Y(n_879) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND3xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_603), .C(n_607), .Y(n_596) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND4xp25_ASAP7_75t_L g609 ( .A(n_610), .B(n_617), .C(n_627), .D(n_636), .Y(n_609) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g774 ( .A(n_616), .Y(n_774) );
INVx2_ASAP7_75t_SL g820 ( .A(n_616), .Y(n_820) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_631), .C(n_633), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g736 ( .A(n_633), .B(n_737), .C(n_741), .Y(n_736) );
NAND3xp33_ASAP7_75t_L g778 ( .A(n_633), .B(n_779), .C(n_782), .Y(n_778) );
NAND3xp33_ASAP7_75t_L g825 ( .A(n_633), .B(n_826), .C(n_827), .Y(n_825) );
NAND3xp33_ASAP7_75t_L g876 ( .A(n_633), .B(n_877), .C(n_878), .Y(n_876) );
NAND3xp33_ASAP7_75t_L g911 ( .A(n_633), .B(n_912), .C(n_914), .Y(n_911) );
AOI33xp33_ASAP7_75t_L g1259 ( .A1(n_633), .A2(n_734), .A3(n_1260), .B1(n_1262), .B2(n_1263), .B3(n_1264), .Y(n_1259) );
INVx3_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .C(n_639), .Y(n_636) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_639), .B(n_743), .C(n_744), .Y(n_742) );
NAND3xp33_ASAP7_75t_L g783 ( .A(n_639), .B(n_784), .C(n_785), .Y(n_783) );
NAND3xp33_ASAP7_75t_L g830 ( .A(n_639), .B(n_831), .C(n_833), .Y(n_830) );
NAND3xp33_ASAP7_75t_L g880 ( .A(n_639), .B(n_881), .C(n_882), .Y(n_880) );
NAND3xp33_ASAP7_75t_L g915 ( .A(n_639), .B(n_916), .C(n_917), .Y(n_915) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
XNOR2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_692), .Y(n_641) );
INVx2_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
AOI211xp5_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_660), .B(n_661), .C(n_682), .Y(n_644) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_656), .Y(n_811) );
OAI31xp33_ASAP7_75t_L g847 ( .A1(n_660), .A2(n_848), .A3(n_849), .B(n_853), .Y(n_847) );
AOI211x1_ASAP7_75t_L g1193 ( .A1(n_660), .A2(n_1194), .B(n_1205), .C(n_1214), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_674), .Y(n_661) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
BUFx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_746), .B2(n_747), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
XNOR2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B(n_706), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_704), .A2(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g950 ( .A(n_704), .Y(n_950) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g759 ( .A(n_708), .Y(n_759) );
AOI31xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_720), .A3(n_723), .B(n_725), .Y(n_714) );
BUFx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AOI31xp33_ASAP7_75t_L g760 ( .A1(n_725), .A2(n_761), .A3(n_765), .B(n_768), .Y(n_760) );
AOI31xp33_ASAP7_75t_L g1271 ( .A1(n_725), .A2(n_1272), .A3(n_1275), .B(n_1278), .Y(n_1271) );
NAND4xp25_ASAP7_75t_L g726 ( .A(n_727), .B(n_731), .C(n_736), .D(n_742), .Y(n_726) );
NAND3xp33_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .C(n_734), .Y(n_731) );
NAND3xp33_ASAP7_75t_L g775 ( .A(n_734), .B(n_776), .C(n_777), .Y(n_775) );
NAND3xp33_ASAP7_75t_L g821 ( .A(n_734), .B(n_822), .C(n_823), .Y(n_821) );
NAND3xp33_ASAP7_75t_L g872 ( .A(n_734), .B(n_873), .C(n_875), .Y(n_872) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g845 ( .A(n_764), .Y(n_845) );
NAND4xp25_ASAP7_75t_L g770 ( .A(n_771), .B(n_775), .C(n_778), .D(n_783), .Y(n_770) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_SL g913 ( .A(n_781), .Y(n_913) );
INVx1_ASAP7_75t_L g1233 ( .A(n_781), .Y(n_1233) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_895), .B1(n_896), .B2(n_987), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
HB1xp67_ASAP7_75t_L g987 ( .A(n_789), .Y(n_987) );
AO22x2_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_791), .B1(n_854), .B2(n_855), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g846 ( .A(n_794), .Y(n_846) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g837 ( .A(n_803), .Y(n_837) );
INVxp67_ASAP7_75t_L g848 ( .A(n_807), .Y(n_848) );
INVxp67_ASAP7_75t_L g853 ( .A(n_813), .Y(n_853) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NAND3xp33_ASAP7_75t_L g835 ( .A(n_816), .B(n_836), .C(n_847), .Y(n_835) );
AND4x1_ASAP7_75t_L g816 ( .A(n_817), .B(n_821), .C(n_825), .D(n_830), .Y(n_816) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
OAI22xp33_ASAP7_75t_L g957 ( .A1(n_841), .A2(n_958), .B1(n_959), .B2(n_960), .Y(n_957) );
OAI22xp33_ASAP7_75t_SL g964 ( .A1(n_841), .A2(n_965), .B1(n_966), .B2(n_968), .Y(n_964) );
INVx3_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_L g926 ( .A(n_842), .Y(n_926) );
HB1xp67_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
NAND4xp25_ASAP7_75t_L g868 ( .A(n_869), .B(n_872), .C(n_876), .D(n_880), .Y(n_868) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
AOI22xp5_ASAP7_75t_L g896 ( .A1(n_897), .A2(n_898), .B1(n_942), .B2(n_943), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
HB1xp67_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
XOR2xp5_ASAP7_75t_L g900 ( .A(n_901), .B(n_941), .Y(n_900) );
NAND3xp33_ASAP7_75t_L g901 ( .A(n_902), .B(n_921), .C(n_931), .Y(n_901) );
AND4x1_ASAP7_75t_L g902 ( .A(n_903), .B(n_907), .C(n_911), .D(n_915), .Y(n_902) );
INVx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
OAI22xp33_ASAP7_75t_L g1020 ( .A1(n_941), .A2(n_1021), .B1(n_1022), .B2(n_1024), .Y(n_1020) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
XNOR2xp5_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .Y(n_944) );
NAND3x1_ASAP7_75t_SL g946 ( .A(n_947), .B(n_955), .C(n_981), .Y(n_946) );
OAI221xp5_ASAP7_75t_L g970 ( .A1(n_958), .A2(n_960), .B1(n_971), .B2(n_973), .C(n_975), .Y(n_970) );
INVxp67_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx3_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
OAI221xp5_ASAP7_75t_L g977 ( .A1(n_971), .A2(n_973), .B1(n_978), .B2(n_979), .C(n_980), .Y(n_977) );
INVx2_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
BUFx3_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
OAI21xp5_ASAP7_75t_L g988 ( .A1(n_989), .A2(n_997), .B(n_1190), .Y(n_988) );
CKINVDCx5p33_ASAP7_75t_R g989 ( .A(n_990), .Y(n_989) );
BUFx3_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx1_ASAP7_75t_L g1069 ( .A(n_991), .Y(n_1069) );
AND2x4_ASAP7_75t_L g991 ( .A(n_992), .B(n_995), .Y(n_991) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_992), .B(n_995), .Y(n_1062) );
HB1xp67_ASAP7_75t_L g1288 ( .A(n_992), .Y(n_1288) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
AND2x4_ASAP7_75t_L g1016 ( .A(n_993), .B(n_995), .Y(n_1016) );
INVx1_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_994), .B(n_1009), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_996), .Y(n_1009) );
NOR3xp33_ASAP7_75t_L g997 ( .A(n_998), .B(n_1130), .C(n_1168), .Y(n_997) );
AOI22xp5_ASAP7_75t_L g998 ( .A1(n_999), .A2(n_1066), .B1(n_1111), .B2(n_1119), .Y(n_998) );
NOR3xp33_ASAP7_75t_SL g999 ( .A(n_1000), .B(n_1076), .C(n_1079), .Y(n_999) );
A2O1A1Ixp33_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1029), .B(n_1037), .C(n_1051), .Y(n_1000) );
O2A1O1Ixp33_ASAP7_75t_L g1186 ( .A1(n_1001), .A2(n_1003), .B(n_1187), .C(n_1188), .Y(n_1186) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1002), .B(n_1033), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1017), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1003), .B(n_1056), .Y(n_1122) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1003), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1003), .B(n_1085), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1003), .B(n_1089), .Y(n_1147) );
NOR2xp33_ASAP7_75t_L g1183 ( .A(n_1003), .B(n_1043), .Y(n_1183) );
INVx4_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
OR2x2_ASAP7_75t_L g1054 ( .A(n_1004), .B(n_1040), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_1004), .B(n_1031), .Y(n_1078) );
INVx3_ASAP7_75t_L g1087 ( .A(n_1004), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1004), .B(n_1083), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_1004), .B(n_1017), .Y(n_1104) );
NOR2xp67_ASAP7_75t_SL g1106 ( .A(n_1004), .B(n_1065), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1004), .B(n_1033), .Y(n_1137) );
NAND3xp33_ASAP7_75t_L g1166 ( .A(n_1004), .B(n_1155), .C(n_1164), .Y(n_1166) );
AOI211xp5_ASAP7_75t_L g1170 ( .A1(n_1004), .A2(n_1098), .B(n_1171), .C(n_1172), .Y(n_1170) );
AND2x4_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1015), .Y(n_1004) );
AND2x4_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1010), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
OR2x2_ASAP7_75t_L g1023 ( .A(n_1008), .B(n_1011), .Y(n_1023) );
HB1xp67_ASAP7_75t_L g1287 ( .A(n_1009), .Y(n_1287) );
AND2x4_ASAP7_75t_L g1012 ( .A(n_1010), .B(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
OR2x2_ASAP7_75t_L g1024 ( .A(n_1011), .B(n_1014), .Y(n_1024) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
INVx2_ASAP7_75t_L g1046 ( .A(n_1016), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1017), .B(n_1034), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1017), .B(n_1122), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_1017), .B(n_1137), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1025), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1018), .B(n_1032), .Y(n_1083) );
INVx1_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_1019), .B(n_1032), .Y(n_1031) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1019), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1019), .B(n_1025), .Y(n_1110) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_1022), .A2(n_1024), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
OAI22xp33_ASAP7_75t_L g1047 ( .A1(n_1022), .A2(n_1048), .B1(n_1049), .B2(n_1050), .Y(n_1047) );
BUFx3_ASAP7_75t_L g1072 ( .A(n_1022), .Y(n_1072) );
BUFx6f_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
HB1xp67_ASAP7_75t_L g1050 ( .A(n_1024), .Y(n_1050) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1024), .Y(n_1075) );
INVx2_ASAP7_75t_L g1032 ( .A(n_1025), .Y(n_1032) );
NOR2xp33_ASAP7_75t_L g1189 ( .A(n_1029), .B(n_1096), .Y(n_1189) );
OR2x2_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1033), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1121 ( .A(n_1031), .B(n_1122), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1031), .B(n_1137), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_1032), .B(n_1056), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_1032), .B(n_1033), .Y(n_1065) );
INVx2_ASAP7_75t_L g1167 ( .A(n_1032), .Y(n_1167) );
OAI322xp33_ASAP7_75t_L g1181 ( .A1(n_1032), .A2(n_1058), .A3(n_1065), .B1(n_1089), .B2(n_1182), .C1(n_1184), .C2(n_1185), .Y(n_1181) );
OR2x2_ASAP7_75t_L g1077 ( .A(n_1033), .B(n_1078), .Y(n_1077) );
OR2x2_ASAP7_75t_L g1099 ( .A(n_1033), .B(n_1090), .Y(n_1099) );
BUFx3_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx2_ASAP7_75t_L g1056 ( .A(n_1034), .Y(n_1056) );
AOI222xp33_ASAP7_75t_L g1105 ( .A1(n_1034), .A2(n_1060), .B1(n_1085), .B2(n_1106), .C1(n_1107), .C2(n_1109), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1034), .B(n_1083), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1034), .B(n_1110), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1036), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1043), .Y(n_1037) );
AOI22xp5_ASAP7_75t_L g1080 ( .A1(n_1038), .A2(n_1081), .B1(n_1084), .B2(n_1086), .Y(n_1080) );
A2O1A1Ixp33_ASAP7_75t_L g1119 ( .A1(n_1038), .A2(n_1120), .B(n_1123), .C(n_1129), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1156 ( .A(n_1038), .B(n_1044), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1175 ( .A(n_1038), .B(n_1176), .Y(n_1175) );
INVx3_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
NOR2xp33_ASAP7_75t_L g1076 ( .A(n_1039), .B(n_1077), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1039), .B(n_1059), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_1039), .B(n_1097), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_1039), .B(n_1118), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g1039 ( .A(n_1040), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1040), .B(n_1060), .Y(n_1085) );
INVx1_ASAP7_75t_SL g1103 ( .A(n_1040), .Y(n_1103) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1040), .Y(n_1143) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1040), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1040), .B(n_1059), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1042), .Y(n_1040) );
OR2x2_ASAP7_75t_L g1058 ( .A(n_1043), .B(n_1059), .Y(n_1058) );
AND2x4_ASAP7_75t_SL g1097 ( .A(n_1043), .B(n_1059), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1043), .B(n_1060), .Y(n_1148) );
INVx2_ASAP7_75t_SL g1043 ( .A(n_1044), .Y(n_1043) );
INVx2_ASAP7_75t_L g1053 ( .A(n_1044), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1044), .B(n_1059), .Y(n_1129) );
INVx2_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
AOI221xp5_ASAP7_75t_L g1051 ( .A1(n_1052), .A2(n_1055), .B1(n_1057), .B2(n_1064), .C(n_1066), .Y(n_1051) );
NOR2xp33_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1054), .Y(n_1052) );
OAI211xp5_ASAP7_75t_SL g1079 ( .A1(n_1053), .A2(n_1080), .B(n_1091), .C(n_1105), .Y(n_1079) );
INVx2_ASAP7_75t_L g1108 ( .A(n_1053), .Y(n_1108) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1053), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1053), .B(n_1067), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1053), .B(n_1085), .Y(n_1172) );
O2A1O1Ixp33_ASAP7_75t_L g1173 ( .A1(n_1053), .A2(n_1174), .B(n_1177), .C(n_1178), .Y(n_1173) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1054), .Y(n_1152) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1055), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_1056), .B(n_1083), .Y(n_1082) );
NOR2x1_ASAP7_75t_L g1089 ( .A(n_1056), .B(n_1090), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1056), .B(n_1110), .Y(n_1109) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1059), .B(n_1124), .Y(n_1163) );
CKINVDCx6p67_ASAP7_75t_R g1059 ( .A(n_1060), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1060), .B(n_1103), .Y(n_1102) );
OR2x6_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1063), .Y(n_1060) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
BUFx3_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
OAI31xp33_ASAP7_75t_L g1131 ( .A1(n_1067), .A2(n_1132), .A3(n_1141), .B(n_1153), .Y(n_1131) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
OAI22xp33_ASAP7_75t_L g1070 ( .A1(n_1071), .A2(n_1072), .B1(n_1073), .B2(n_1074), .Y(n_1070) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1077), .Y(n_1177) );
OAI31xp33_ASAP7_75t_SL g1139 ( .A1(n_1081), .A2(n_1134), .A3(n_1136), .B(n_1140), .Y(n_1139) );
OAI21xp5_ASAP7_75t_L g1146 ( .A1(n_1081), .A2(n_1147), .B(n_1148), .Y(n_1146) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1083), .Y(n_1161) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_1084), .A2(n_1087), .B1(n_1113), .B2(n_1115), .Y(n_1112) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_1085), .B(n_1183), .Y(n_1182) );
NOR2xp33_ASAP7_75t_L g1086 ( .A(n_1087), .B(n_1088), .Y(n_1086) );
INVx2_ASAP7_75t_L g1114 ( .A(n_1087), .Y(n_1114) );
AOI22xp5_ASAP7_75t_L g1123 ( .A1(n_1087), .A2(n_1124), .B1(n_1125), .B2(n_1127), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1087), .B(n_1126), .Y(n_1157) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1090), .Y(n_1116) );
AOI221xp5_ASAP7_75t_L g1091 ( .A1(n_1092), .A2(n_1094), .B1(n_1095), .B2(n_1098), .C(n_1100), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_1094), .B(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1094), .Y(n_1138) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1097), .Y(n_1169) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
NOR2xp33_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1104), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1102), .B(n_1108), .Y(n_1107) );
OAI21xp5_ASAP7_75t_SL g1179 ( .A1(n_1102), .A2(n_1126), .B(n_1147), .Y(n_1179) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1106), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1107), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1109), .B(n_1114), .Y(n_1118) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1110), .Y(n_1162) );
AOI21xp33_ASAP7_75t_L g1111 ( .A1(n_1112), .A2(n_1116), .B(n_1117), .Y(n_1111) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
OAI21xp33_ASAP7_75t_L g1149 ( .A1(n_1128), .A2(n_1150), .B(n_1152), .Y(n_1149) );
NAND2xp5_ASAP7_75t_SL g1130 ( .A(n_1131), .B(n_1158), .Y(n_1130) );
A2O1A1Ixp33_ASAP7_75t_L g1132 ( .A1(n_1133), .A2(n_1135), .B(n_1138), .C(n_1139), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
A2O1A1Ixp33_ASAP7_75t_L g1178 ( .A1(n_1138), .A2(n_1144), .B(n_1176), .C(n_1179), .Y(n_1178) );
OAI211xp5_ASAP7_75t_SL g1141 ( .A1(n_1142), .A2(n_1144), .B(n_1146), .C(n_1149), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1148), .B(n_1151), .Y(n_1150) );
AOI21xp33_ASAP7_75t_L g1153 ( .A1(n_1154), .A2(n_1156), .B(n_1157), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
AOI32xp33_ASAP7_75t_L g1158 ( .A1(n_1159), .A2(n_1163), .A3(n_1164), .B1(n_1165), .B2(n_1167), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1162), .Y(n_1160) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
OAI211xp5_ASAP7_75t_SL g1168 ( .A1(n_1169), .A2(n_1170), .B(n_1173), .C(n_1180), .Y(n_1168) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1172), .Y(n_1188) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
NOR3xp33_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1186), .C(n_1189), .Y(n_1180) );
INVx2_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1223), .Y(n_1214) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1245), .Y(n_1280) );
HB1xp67_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1265), .Y(n_1258) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
CKINVDCx5p33_ASAP7_75t_R g1282 ( .A(n_1283), .Y(n_1282) );
A2O1A1Ixp33_ASAP7_75t_L g1285 ( .A1(n_1284), .A2(n_1286), .B(n_1288), .C(n_1289), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
endmodule