module fake_jpeg_12451_n_57 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_57);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_57;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_5),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_20),
.Y(n_24)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_0),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_14),
.B1(n_10),
.B2(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_22),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_21),
.A2(n_8),
.B1(n_14),
.B2(n_11),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_27),
.B(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_30),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_28),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_24),
.C(n_27),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_23),
.C(n_12),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_37),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

OAI21x1_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_42),
.B(n_43),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_19),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_35),
.B(n_32),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_47),
.B(n_48),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_12),
.B1(n_10),
.B2(n_32),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_49),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_52),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_7),
.C(n_2),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_2),
.B(n_4),
.Y(n_54)
);

MAJx2_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_52),
.C(n_4),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_55),
.B(n_53),
.Y(n_56)
);

BUFx24_ASAP7_75t_SL g57 ( 
.A(n_56),
.Y(n_57)
);


endmodule