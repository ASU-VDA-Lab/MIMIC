module real_jpeg_25556_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_1),
.B(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_17),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_13),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_5),
.B(n_13),
.Y(n_15)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_5),
.A2(n_18),
.B(n_19),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_5),
.B(n_18),
.Y(n_19)
);

AOI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_16),
.B(n_20),
.C(n_28),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_8),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_10),
.Y(n_8)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_9),
.B(n_35),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_9),
.B(n_35),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_10),
.A2(n_11),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g10 ( 
.A(n_11),
.Y(n_10)
);

OR2x2_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_14),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_17),
.B(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_17),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_31),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp33_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_32),
.B(n_33),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);


endmodule