module fake_jpeg_390_n_110 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_44),
.Y(n_46)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_0),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_34),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_61),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_41),
.B1(n_35),
.B2(n_32),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_30),
.B1(n_31),
.B2(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_63),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_54),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_64),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_30),
.B1(n_36),
.B2(n_29),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_36),
.B1(n_35),
.B2(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_31),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_19),
.B(n_10),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_75),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_56),
.B1(n_5),
.B2(n_6),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_28),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_74),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_1),
.B(n_3),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_4),
.B(n_5),
.C(n_7),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_3),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_4),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_17),
.C(n_25),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_83),
.C(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_7),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

AO22x1_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_13),
.B1(n_24),
.B2(n_22),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_8),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_26),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_18),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_8),
.B(n_9),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_11),
.C(n_12),
.Y(n_100)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_94),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_83),
.B1(n_70),
.B2(n_77),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_100),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_70),
.B1(n_11),
.B2(n_12),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_95),
.C(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_103),
.C(n_94),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_97),
.B(n_88),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_99),
.B(n_87),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_93),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_100),
.Y(n_110)
);


endmodule