module fake_aes_6991_n_1152 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1152);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1152;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_360;
wire n_345;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1016;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_1042;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_638;
wire n_563;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1025;
wire n_1011;
wire n_1132;
wire n_880;
wire n_1101;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_1138;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_950;
wire n_427;
wire n_910;
wire n_935;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_666;
wire n_621;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_1125;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_924;
wire n_912;
wire n_1043;
wire n_947;
wire n_378;
wire n_582;
wire n_1141;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1007;
wire n_859;
wire n_1117;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_1146;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_257;
wire n_992;
wire n_1127;
wire n_269;
INVx1_ASAP7_75t_L g252 ( .A(n_189), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_56), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_42), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_152), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_246), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_120), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_235), .Y(n_258) );
OR2x2_ASAP7_75t_L g259 ( .A(n_51), .B(n_114), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_118), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_2), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_4), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_150), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_86), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_28), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_225), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_166), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_222), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_91), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_87), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_161), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_18), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_132), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_100), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_220), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_5), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_117), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_247), .Y(n_278) );
INVxp33_ASAP7_75t_SL g279 ( .A(n_0), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_71), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_148), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_176), .Y(n_282) );
INVxp33_ASAP7_75t_L g283 ( .A(n_8), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_48), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_197), .Y(n_285) );
CKINVDCx16_ASAP7_75t_R g286 ( .A(n_58), .Y(n_286) );
BUFx10_ASAP7_75t_L g287 ( .A(n_19), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_52), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_165), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_66), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_45), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_137), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_214), .Y(n_293) );
CKINVDCx14_ASAP7_75t_R g294 ( .A(n_216), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_123), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_5), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_142), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_251), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_155), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_80), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_8), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_9), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_11), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_30), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_105), .Y(n_305) );
CKINVDCx16_ASAP7_75t_R g306 ( .A(n_179), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_92), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_218), .Y(n_308) );
INVx1_ASAP7_75t_SL g309 ( .A(n_49), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_199), .Y(n_310) );
BUFx10_ASAP7_75t_L g311 ( .A(n_210), .Y(n_311) );
BUFx5_ASAP7_75t_L g312 ( .A(n_208), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_81), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_133), .Y(n_314) );
INVxp33_ASAP7_75t_SL g315 ( .A(n_221), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_71), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_42), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_99), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_248), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_206), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_18), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_237), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_122), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_154), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_126), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_219), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_198), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_157), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_93), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_191), .Y(n_330) );
CKINVDCx16_ASAP7_75t_R g331 ( .A(n_115), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_46), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_51), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_141), .B(n_139), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_34), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_108), .Y(n_336) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_4), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_19), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_40), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_88), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_135), .Y(n_341) );
CKINVDCx16_ASAP7_75t_R g342 ( .A(n_232), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_9), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_104), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_20), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_187), .Y(n_346) );
INVxp67_ASAP7_75t_SL g347 ( .A(n_239), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_245), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_20), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_74), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_162), .Y(n_351) );
INVx1_ASAP7_75t_SL g352 ( .A(n_52), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_63), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_60), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_159), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_46), .B(n_175), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_146), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_125), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_134), .Y(n_359) );
INVx2_ASAP7_75t_SL g360 ( .A(n_119), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_138), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_173), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_85), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_47), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_164), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_243), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_169), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_209), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_156), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_94), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_63), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_95), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_59), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_145), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_200), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_229), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_70), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_116), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_36), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_33), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_136), .Y(n_381) );
BUFx10_ASAP7_75t_L g382 ( .A(n_3), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_180), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_312), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_376), .B(n_1), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_321), .Y(n_386) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_298), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_298), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_286), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_283), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_289), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_312), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_283), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_306), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_255), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_321), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_360), .B(n_6), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_276), .B(n_6), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_255), .B(n_7), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_312), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_294), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_252), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_294), .B(n_7), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_312), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_256), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_275), .B(n_10), .Y(n_406) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_298), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_331), .B(n_10), .Y(n_408) );
OAI22xp5_ASAP7_75t_SL g409 ( .A1(n_265), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_253), .B(n_12), .Y(n_410) );
OAI21x1_ASAP7_75t_L g411 ( .A1(n_275), .A2(n_78), .B(n_77), .Y(n_411) );
OAI22xp5_ASAP7_75t_SL g412 ( .A1(n_265), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_312), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_342), .B(n_14), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_260), .Y(n_415) );
NOR2x1_ASAP7_75t_L g416 ( .A(n_264), .B(n_15), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_387), .Y(n_417) );
INVx6_ASAP7_75t_L g418 ( .A(n_406), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_390), .B(n_311), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_384), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_395), .B(n_326), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_384), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_384), .Y(n_423) );
BUFx10_ASAP7_75t_L g424 ( .A(n_406), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_392), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_387), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_401), .B(n_323), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_395), .B(n_326), .Y(n_428) );
AND2x2_ASAP7_75t_SL g429 ( .A(n_406), .B(n_259), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_392), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_395), .B(n_363), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_390), .B(n_393), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_393), .B(n_311), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_401), .B(n_309), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_387), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_395), .B(n_363), .Y(n_436) );
INVx2_ASAP7_75t_SL g437 ( .A(n_391), .Y(n_437) );
INVx4_ASAP7_75t_L g438 ( .A(n_406), .Y(n_438) );
INVx3_ASAP7_75t_L g439 ( .A(n_406), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_402), .A2(n_261), .B1(n_272), .B2(n_262), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_391), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_387), .Y(n_442) );
INVx4_ASAP7_75t_L g443 ( .A(n_395), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_402), .A2(n_296), .B1(n_303), .B2(n_301), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_401), .B(n_266), .Y(n_445) );
INVx4_ASAP7_75t_L g446 ( .A(n_391), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_405), .B(n_312), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_405), .B(n_267), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_387), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_387), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_398), .B(n_287), .Y(n_451) );
AND3x2_ASAP7_75t_L g452 ( .A(n_408), .B(n_338), .C(n_356), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_415), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_398), .B(n_352), .Y(n_454) );
NOR2x1p5_ASAP7_75t_L g455 ( .A(n_394), .B(n_254), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_392), .Y(n_456) );
INVx4_ASAP7_75t_L g457 ( .A(n_403), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_400), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_415), .B(n_268), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_398), .B(n_287), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_386), .B(n_269), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_387), .Y(n_462) );
INVx8_ASAP7_75t_L g463 ( .A(n_403), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_400), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_429), .A2(n_403), .B1(n_414), .B2(n_408), .Y(n_465) );
OAI22xp5_ASAP7_75t_SL g466 ( .A1(n_454), .A2(n_412), .B1(n_409), .B2(n_280), .Y(n_466) );
NAND3xp33_ASAP7_75t_SL g467 ( .A(n_432), .B(n_394), .C(n_389), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_457), .B(n_445), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_457), .B(n_414), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_457), .B(n_414), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_457), .B(n_397), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_443), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_432), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_463), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_453), .B(n_400), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_443), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_432), .B(n_410), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_445), .B(n_397), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_463), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_453), .B(n_404), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_451), .B(n_460), .Y(n_481) );
O2A1O1Ixp5_ASAP7_75t_L g482 ( .A1(n_447), .A2(n_399), .B(n_385), .C(n_410), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_429), .A2(n_399), .B1(n_385), .B2(n_416), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_427), .B(n_416), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_453), .B(n_404), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_443), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_427), .B(n_386), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_434), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_451), .B(n_382), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_443), .Y(n_490) );
INVx3_ASAP7_75t_L g491 ( .A(n_443), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_463), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_419), .B(n_396), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_463), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_419), .B(n_396), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_451), .B(n_389), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_419), .B(n_258), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_433), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_424), .B(n_404), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_433), .B(n_263), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_463), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_433), .A2(n_310), .B1(n_319), .B2(n_257), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_424), .B(n_413), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_460), .B(n_277), .Y(n_504) );
INVx1_ASAP7_75t_SL g505 ( .A(n_434), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_460), .B(n_278), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_438), .B(n_315), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_418), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_424), .B(n_413), .Y(n_509) );
BUFx12f_ASAP7_75t_L g510 ( .A(n_455), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_438), .B(n_281), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_420), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_424), .B(n_413), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_454), .B(n_382), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_418), .Y(n_515) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_424), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_422), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_438), .B(n_270), .Y(n_518) );
INVx3_ASAP7_75t_L g519 ( .A(n_418), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_418), .Y(n_520) );
OR2x6_ASAP7_75t_L g521 ( .A(n_434), .B(n_412), .Y(n_521) );
INVx3_ASAP7_75t_L g522 ( .A(n_418), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_429), .B(n_285), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_422), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_454), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_439), .B(n_271), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_429), .A2(n_279), .B1(n_317), .B2(n_316), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_439), .B(n_305), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_439), .B(n_308), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_455), .A2(n_310), .B1(n_319), .B2(n_257), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_439), .A2(n_369), .B1(n_409), .B2(n_304), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_439), .B(n_313), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_459), .A2(n_339), .B1(n_343), .B2(n_332), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_421), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_421), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_428), .Y(n_536) );
NOR2xp33_ASAP7_75t_SL g537 ( .A(n_452), .B(n_369), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_448), .B(n_273), .Y(n_538) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_459), .A2(n_411), .B(n_349), .C(n_354), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_448), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_431), .B(n_336), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_452), .A2(n_333), .B1(n_335), .B2(n_291), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_440), .A2(n_380), .B1(n_364), .B2(n_371), .Y(n_543) );
INVx6_ASAP7_75t_L g544 ( .A(n_446), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_431), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_436), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_436), .B(n_344), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_461), .A2(n_411), .B(n_373), .C(n_377), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_437), .A2(n_411), .B(n_347), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_423), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_465), .A2(n_444), .B1(n_440), .B2(n_461), .Y(n_551) );
INVx3_ASAP7_75t_SL g552 ( .A(n_498), .Y(n_552) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_516), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_540), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_477), .B(n_444), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_519), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_519), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_516), .B(n_441), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_534), .B(n_441), .Y(n_559) );
AND2x6_ASAP7_75t_L g560 ( .A(n_474), .B(n_441), .Y(n_560) );
O2A1O1Ixp33_ASAP7_75t_L g561 ( .A1(n_525), .A2(n_425), .B(n_430), .C(n_423), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g562 ( .A1(n_526), .A2(n_430), .B(n_456), .C(n_425), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_535), .B(n_441), .Y(n_563) );
OAI21x1_ASAP7_75t_L g564 ( .A1(n_549), .A2(n_458), .B(n_456), .Y(n_564) );
AND3x2_ASAP7_75t_L g565 ( .A(n_537), .B(n_284), .C(n_280), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_499), .A2(n_437), .B(n_446), .Y(n_566) );
AOI21x1_ASAP7_75t_L g567 ( .A1(n_518), .A2(n_464), .B(n_458), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_536), .Y(n_568) );
OAI22x1_ASAP7_75t_L g569 ( .A1(n_531), .A2(n_288), .B1(n_290), .B2(n_284), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_505), .B(n_345), .Y(n_570) );
O2A1O1Ixp33_ASAP7_75t_SL g571 ( .A1(n_539), .A2(n_548), .B(n_480), .C(n_485), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_488), .B(n_288), .Y(n_572) );
OR2x6_ASAP7_75t_L g573 ( .A(n_474), .B(n_379), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_516), .B(n_446), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_473), .B(n_446), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_545), .B(n_446), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_546), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_478), .B(n_464), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_503), .A2(n_435), .B(n_426), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_481), .B(n_290), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_503), .A2(n_435), .B(n_426), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_481), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_516), .B(n_351), .Y(n_583) );
AO22x1_ASAP7_75t_L g584 ( .A1(n_496), .A2(n_337), .B1(n_353), .B2(n_302), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_509), .A2(n_435), .B(n_426), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_479), .A2(n_337), .B1(n_353), .B2(n_302), .Y(n_586) );
INVx2_ASAP7_75t_SL g587 ( .A(n_514), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_469), .A2(n_282), .B1(n_292), .B2(n_274), .Y(n_588) );
BUFx2_ASAP7_75t_L g589 ( .A(n_479), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_522), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_470), .B(n_356), .Y(n_591) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_491), .Y(n_592) );
AOI21xp33_ASAP7_75t_L g593 ( .A1(n_523), .A2(n_359), .B(n_357), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_509), .A2(n_450), .B(n_449), .Y(n_594) );
AO21x1_ASAP7_75t_L g595 ( .A1(n_526), .A2(n_295), .B(n_293), .Y(n_595) );
A2O1A1Ixp33_ASAP7_75t_L g596 ( .A1(n_538), .A2(n_297), .B(n_300), .C(n_299), .Y(n_596) );
NOR3xp33_ASAP7_75t_SL g597 ( .A(n_466), .B(n_365), .C(n_361), .Y(n_597) );
OAI22x1_ASAP7_75t_L g598 ( .A1(n_502), .A2(n_530), .B1(n_496), .B2(n_542), .Y(n_598) );
AO32x1_ASAP7_75t_L g599 ( .A1(n_539), .A2(n_348), .A3(n_307), .B1(n_314), .B2(n_330), .Y(n_599) );
A2O1A1Ixp33_ASAP7_75t_L g600 ( .A1(n_482), .A2(n_318), .B(n_322), .C(n_320), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_468), .B(n_366), .Y(n_601) );
BUFx2_ASAP7_75t_L g602 ( .A(n_489), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_522), .Y(n_603) );
NAND2x1p5_ASAP7_75t_L g604 ( .A(n_492), .B(n_350), .Y(n_604) );
NAND3xp33_ASAP7_75t_SL g605 ( .A(n_483), .B(n_375), .C(n_368), .Y(n_605) );
INVx1_ASAP7_75t_SL g606 ( .A(n_494), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_513), .A2(n_450), .B(n_449), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_471), .A2(n_325), .B1(n_340), .B2(n_328), .Y(n_608) );
AND2x4_ASAP7_75t_L g609 ( .A(n_493), .B(n_341), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_527), .A2(n_370), .B1(n_346), .B2(n_374), .Y(n_610) );
A2O1A1Ixp33_ASAP7_75t_L g611 ( .A1(n_507), .A2(n_367), .B(n_383), .C(n_355), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_496), .B(n_350), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_467), .B(n_16), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_513), .A2(n_450), .B(n_449), .Y(n_614) );
OAI21xp33_ASAP7_75t_SL g615 ( .A1(n_484), .A2(n_362), .B(n_358), .Y(n_615) );
NOR2x1p5_ASAP7_75t_SL g616 ( .A(n_512), .B(n_417), .Y(n_616) );
NOR2xp33_ASAP7_75t_SL g617 ( .A(n_501), .B(n_334), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_487), .A2(n_378), .B1(n_381), .B2(n_350), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_518), .A2(n_462), .B(n_442), .Y(n_619) );
BUFx3_ASAP7_75t_L g620 ( .A(n_510), .Y(n_620) );
AO32x2_ASAP7_75t_L g621 ( .A1(n_548), .A2(n_407), .A3(n_388), .B1(n_324), .B2(n_327), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_533), .A2(n_289), .B1(n_372), .B2(n_329), .C(n_298), .Y(n_622) );
NOR2x1_ASAP7_75t_R g623 ( .A(n_510), .B(n_324), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_475), .A2(n_462), .B(n_442), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_495), .A2(n_324), .B1(n_327), .B2(n_329), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_497), .B(n_16), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_475), .A2(n_462), .B(n_442), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_517), .A2(n_372), .B1(n_327), .B2(n_329), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_480), .A2(n_442), .B(n_417), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_500), .B(n_17), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_485), .A2(n_417), .B(n_327), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_504), .B(n_17), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_486), .A2(n_417), .B(n_372), .Y(n_633) );
O2A1O1Ixp33_ASAP7_75t_SL g634 ( .A1(n_528), .A2(n_131), .B(n_178), .C(n_250), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_517), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_524), .Y(n_636) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_524), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_521), .Y(n_638) );
NOR2xp33_ASAP7_75t_SL g639 ( .A(n_550), .B(n_388), .Y(n_639) );
A2O1A1Ixp33_ASAP7_75t_L g640 ( .A1(n_507), .A2(n_407), .B(n_388), .C(n_23), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_506), .B(n_21), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_521), .B(n_21), .Y(n_642) );
O2A1O1Ixp33_ASAP7_75t_L g643 ( .A1(n_521), .A2(n_22), .B(n_23), .C(n_24), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_508), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_490), .A2(n_407), .B(n_388), .C(n_25), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_472), .A2(n_407), .B1(n_388), .B2(n_25), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_472), .Y(n_647) );
AND2x2_ASAP7_75t_SL g648 ( .A(n_543), .B(n_22), .Y(n_648) );
NAND2x1p5_ASAP7_75t_L g649 ( .A(n_476), .B(n_388), .Y(n_649) );
NOR2xp67_ASAP7_75t_SL g650 ( .A(n_544), .B(n_388), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_541), .B(n_24), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_547), .B(n_26), .Y(n_652) );
AOI21x1_ASAP7_75t_L g653 ( .A1(n_529), .A2(n_407), .B(n_79), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_476), .B(n_26), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_532), .A2(n_407), .B(n_82), .Y(n_655) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_511), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_L g657 ( .A1(n_515), .A2(n_27), .B(n_28), .C(n_29), .Y(n_657) );
INVxp67_ASAP7_75t_SL g658 ( .A(n_520), .Y(n_658) );
NOR3xp33_ASAP7_75t_SL g659 ( .A(n_544), .B(n_29), .C(n_30), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_544), .B(n_31), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_465), .A2(n_32), .B1(n_34), .B2(n_35), .Y(n_661) );
BUFx12f_ASAP7_75t_L g662 ( .A(n_510), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_499), .A2(n_84), .B(n_83), .Y(n_663) );
O2A1O1Ixp33_ASAP7_75t_L g664 ( .A1(n_525), .A2(n_35), .B(n_36), .C(n_37), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_540), .B(n_37), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_510), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_505), .B(n_38), .Y(n_667) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_505), .Y(n_668) );
OAI21xp33_ASAP7_75t_L g669 ( .A1(n_465), .A2(n_38), .B(n_39), .Y(n_669) );
A2O1A1Ixp33_ASAP7_75t_L g670 ( .A1(n_632), .A2(n_39), .B(n_40), .C(n_41), .Y(n_670) );
OR2x2_ASAP7_75t_L g671 ( .A(n_586), .B(n_41), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_573), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_672) );
O2A1O1Ixp33_ASAP7_75t_L g673 ( .A1(n_611), .A2(n_43), .B(n_44), .C(n_47), .Y(n_673) );
OAI21xp5_ASAP7_75t_L g674 ( .A1(n_562), .A2(n_158), .B(n_244), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_648), .A2(n_598), .B1(n_668), .B2(n_580), .Y(n_675) );
INVxp67_ASAP7_75t_SL g676 ( .A(n_589), .Y(n_676) );
OAI221xp5_ASAP7_75t_SL g677 ( .A1(n_613), .A2(n_48), .B1(n_49), .B2(n_50), .C(n_53), .Y(n_677) );
AND2x4_ASAP7_75t_L g678 ( .A(n_554), .B(n_50), .Y(n_678) );
O2A1O1Ixp33_ASAP7_75t_SL g679 ( .A1(n_640), .A2(n_160), .B(n_242), .C(n_241), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_568), .Y(n_680) );
A2O1A1Ixp33_ASAP7_75t_L g681 ( .A1(n_630), .A2(n_53), .B(n_54), .C(n_55), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_578), .A2(n_153), .B(n_240), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_577), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_573), .A2(n_54), .B1(n_55), .B2(n_56), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_555), .B(n_57), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_573), .A2(n_57), .B1(n_58), .B2(n_59), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_602), .B(n_60), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_587), .B(n_61), .Y(n_688) );
BUFx3_ASAP7_75t_L g689 ( .A(n_662), .Y(n_689) );
OAI22xp33_ASAP7_75t_L g690 ( .A1(n_569), .A2(n_61), .B1(n_62), .B2(n_64), .Y(n_690) );
A2O1A1Ixp33_ASAP7_75t_L g691 ( .A1(n_651), .A2(n_62), .B(n_64), .C(n_65), .Y(n_691) );
CKINVDCx5p33_ASAP7_75t_R g692 ( .A(n_666), .Y(n_692) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_572), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_693) );
O2A1O1Ixp33_ASAP7_75t_SL g694 ( .A1(n_645), .A2(n_172), .B(n_238), .C(n_236), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_551), .A2(n_67), .B1(n_68), .B2(n_69), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g696 ( .A1(n_652), .A2(n_68), .B(n_69), .C(n_70), .Y(n_696) );
OR2x2_ASAP7_75t_L g697 ( .A(n_584), .B(n_72), .Y(n_697) );
AO31x2_ASAP7_75t_L g698 ( .A1(n_595), .A2(n_72), .A3(n_73), .B(n_74), .Y(n_698) );
BUFx5_ASAP7_75t_L g699 ( .A(n_560), .Y(n_699) );
O2A1O1Ixp33_ASAP7_75t_L g700 ( .A1(n_596), .A2(n_73), .B(n_75), .C(n_76), .Y(n_700) );
BUFx3_ASAP7_75t_L g701 ( .A(n_620), .Y(n_701) );
A2O1A1Ixp33_ASAP7_75t_L g702 ( .A1(n_561), .A2(n_75), .B(n_76), .C(n_89), .Y(n_702) );
AO31x2_ASAP7_75t_L g703 ( .A1(n_625), .A2(n_90), .A3(n_96), .B(n_97), .Y(n_703) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_553), .Y(n_704) );
OAI21xp5_ASAP7_75t_L g705 ( .A1(n_576), .A2(n_98), .B(n_101), .Y(n_705) );
AND2x4_ASAP7_75t_L g706 ( .A(n_582), .B(n_102), .Y(n_706) );
A2O1A1Ixp33_ASAP7_75t_L g707 ( .A1(n_669), .A2(n_103), .B(n_106), .C(n_107), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_635), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_L g709 ( .A1(n_615), .A2(n_109), .B(n_110), .C(n_111), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_552), .B(n_112), .Y(n_710) );
CKINVDCx5p33_ASAP7_75t_R g711 ( .A(n_638), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g712 ( .A1(n_641), .A2(n_113), .B(n_121), .C(n_124), .Y(n_712) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_553), .B(n_127), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_636), .Y(n_714) );
BUFx4_ASAP7_75t_R g715 ( .A(n_623), .Y(n_715) );
AND2x4_ASAP7_75t_L g716 ( .A(n_612), .B(n_128), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_665), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_644), .Y(n_718) );
AND2x4_ASAP7_75t_L g719 ( .A(n_656), .B(n_249), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_570), .B(n_129), .Y(n_720) );
A2O1A1Ixp33_ASAP7_75t_L g721 ( .A1(n_626), .A2(n_130), .B(n_140), .C(n_143), .Y(n_721) );
O2A1O1Ixp33_ASAP7_75t_L g722 ( .A1(n_551), .A2(n_144), .B(n_147), .C(n_149), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_610), .B(n_151), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g724 ( .A1(n_657), .A2(n_163), .B(n_167), .C(n_168), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_661), .Y(n_725) );
AOI221xp5_ASAP7_75t_L g726 ( .A1(n_610), .A2(n_170), .B1(n_171), .B2(n_174), .C(n_177), .Y(n_726) );
AO31x2_ASAP7_75t_L g727 ( .A1(n_625), .A2(n_181), .A3(n_182), .B(n_183), .Y(n_727) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_565), .A2(n_184), .B1(n_185), .B2(n_186), .Y(n_728) );
AO32x2_ASAP7_75t_L g729 ( .A1(n_618), .A2(n_188), .A3(n_190), .B1(n_192), .B2(n_193), .Y(n_729) );
AO31x2_ASAP7_75t_L g730 ( .A1(n_618), .A2(n_194), .A3(n_195), .B(n_196), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_566), .A2(n_201), .B(n_202), .Y(n_731) );
OAI22xp33_ASAP7_75t_L g732 ( .A1(n_606), .A2(n_203), .B1(n_204), .B2(n_205), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_559), .A2(n_207), .B(n_211), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_637), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_609), .B(n_212), .Y(n_735) );
OR2x2_ASAP7_75t_L g736 ( .A(n_609), .B(n_213), .Y(n_736) );
O2A1O1Ixp33_ASAP7_75t_L g737 ( .A1(n_591), .A2(n_215), .B(n_217), .C(n_223), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_593), .B(n_224), .Y(n_738) );
OA21x2_ASAP7_75t_L g739 ( .A1(n_655), .A2(n_226), .B(n_227), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_642), .A2(n_228), .B1(n_230), .B2(n_231), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_563), .A2(n_233), .B(n_234), .Y(n_741) );
O2A1O1Ixp33_ASAP7_75t_L g742 ( .A1(n_588), .A2(n_608), .B(n_664), .C(n_643), .Y(n_742) );
OR2x2_ASAP7_75t_L g743 ( .A(n_608), .B(n_588), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_667), .A2(n_605), .B1(n_575), .B2(n_601), .Y(n_744) );
O2A1O1Ixp33_ASAP7_75t_L g745 ( .A1(n_654), .A2(n_617), .B(n_659), .C(n_660), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_579), .A2(n_594), .B(n_581), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_597), .B(n_604), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_585), .A2(n_607), .B(n_614), .Y(n_748) );
OR2x2_ASAP7_75t_L g749 ( .A(n_590), .B(n_603), .Y(n_749) );
O2A1O1Ixp33_ASAP7_75t_L g750 ( .A1(n_617), .A2(n_622), .B(n_583), .C(n_556), .Y(n_750) );
INVx3_ASAP7_75t_SL g751 ( .A(n_560), .Y(n_751) );
A2O1A1Ixp33_ASAP7_75t_L g752 ( .A1(n_616), .A2(n_647), .B(n_633), .C(n_631), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g753 ( .A1(n_619), .A2(n_558), .B(n_574), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_567), .Y(n_754) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_560), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_629), .A2(n_627), .B(n_624), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_557), .Y(n_757) );
INVx4_ASAP7_75t_L g758 ( .A(n_560), .Y(n_758) );
INVx3_ASAP7_75t_L g759 ( .A(n_592), .Y(n_759) );
OR2x2_ASAP7_75t_L g760 ( .A(n_649), .B(n_658), .Y(n_760) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_628), .Y(n_761) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_621), .Y(n_762) );
AOI31xp67_ASAP7_75t_L g763 ( .A1(n_621), .A2(n_599), .A3(n_634), .B(n_639), .Y(n_763) );
CKINVDCx5p33_ASAP7_75t_R g764 ( .A(n_646), .Y(n_764) );
AOI21xp33_ASAP7_75t_L g765 ( .A1(n_650), .A2(n_663), .B(n_599), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_599), .A2(n_571), .B(n_549), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_621), .A2(n_465), .B1(n_457), .B2(n_540), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_568), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_568), .Y(n_769) );
BUFx3_ASAP7_75t_L g770 ( .A(n_662), .Y(n_770) );
BUFx6f_ASAP7_75t_L g771 ( .A(n_553), .Y(n_771) );
A2O1A1Ixp33_ASAP7_75t_L g772 ( .A1(n_632), .A2(n_630), .B(n_652), .C(n_651), .Y(n_772) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_668), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_571), .A2(n_549), .B(n_578), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_648), .A2(n_496), .B1(n_467), .B2(n_521), .Y(n_775) );
CKINVDCx5p33_ASAP7_75t_R g776 ( .A(n_662), .Y(n_776) );
OAI21x1_ASAP7_75t_L g777 ( .A1(n_564), .A2(n_653), .B(n_549), .Y(n_777) );
INVx3_ASAP7_75t_L g778 ( .A(n_553), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_602), .B(n_505), .Y(n_779) );
A2O1A1Ixp33_ASAP7_75t_L g780 ( .A1(n_632), .A2(n_630), .B(n_652), .C(n_651), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g781 ( .A1(n_571), .A2(n_549), .B(n_578), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_554), .B(n_540), .Y(n_782) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_662), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_568), .Y(n_784) );
BUFx10_ASAP7_75t_L g785 ( .A(n_668), .Y(n_785) );
OAI21xp5_ASAP7_75t_L g786 ( .A1(n_562), .A2(n_539), .B(n_548), .Y(n_786) );
INVx2_ASAP7_75t_SL g787 ( .A(n_668), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_568), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_668), .B(n_505), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_568), .Y(n_790) );
AO31x2_ASAP7_75t_L g791 ( .A1(n_595), .A2(n_539), .A3(n_548), .B(n_640), .Y(n_791) );
O2A1O1Ixp33_ASAP7_75t_SL g792 ( .A1(n_600), .A2(n_640), .B(n_562), .C(n_539), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_573), .A2(n_465), .B1(n_457), .B2(n_540), .Y(n_793) );
O2A1O1Ixp33_ASAP7_75t_SL g794 ( .A1(n_600), .A2(n_640), .B(n_562), .C(n_539), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_743), .B(n_680), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_675), .A2(n_775), .B1(n_793), .B2(n_764), .Y(n_796) );
INVx2_ASAP7_75t_SL g797 ( .A(n_689), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_782), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_725), .B(n_683), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_776), .Y(n_800) );
AOI21xp5_ASAP7_75t_L g801 ( .A1(n_746), .A2(n_748), .B(n_786), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_768), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_769), .B(n_784), .Y(n_803) );
INVx2_ASAP7_75t_SL g804 ( .A(n_770), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_788), .Y(n_805) );
INVx2_ASAP7_75t_SL g806 ( .A(n_785), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_790), .Y(n_807) );
OR2x6_ASAP7_75t_L g808 ( .A(n_758), .B(n_719), .Y(n_808) );
AOI22xp5_ASAP7_75t_SL g809 ( .A1(n_678), .A2(n_715), .B1(n_719), .B2(n_711), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_779), .B(n_789), .Y(n_810) );
INVx1_ASAP7_75t_SL g811 ( .A(n_760), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g812 ( .A1(n_756), .A2(n_780), .B(n_772), .Y(n_812) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_773), .Y(n_813) );
OR2x2_ASAP7_75t_L g814 ( .A(n_787), .B(n_671), .Y(n_814) );
OAI22xp33_ASAP7_75t_L g815 ( .A1(n_697), .A2(n_736), .B1(n_751), .B2(n_678), .Y(n_815) );
AO31x2_ASAP7_75t_L g816 ( .A1(n_754), .A2(n_752), .A3(n_707), .B(n_767), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_687), .A2(n_723), .B1(n_717), .B2(n_688), .Y(n_817) );
A2O1A1Ixp33_ASAP7_75t_L g818 ( .A1(n_742), .A2(n_745), .B(n_673), .C(n_700), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_708), .Y(n_819) );
A2O1A1Ixp33_ASAP7_75t_L g820 ( .A1(n_750), .A2(n_722), .B(n_738), .C(n_702), .Y(n_820) );
AOI21xp5_ASAP7_75t_L g821 ( .A1(n_794), .A2(n_792), .B(n_753), .Y(n_821) );
OR2x2_ASAP7_75t_L g822 ( .A(n_676), .B(n_701), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_718), .Y(n_823) );
NAND2xp5_ASAP7_75t_SL g824 ( .A(n_785), .B(n_706), .Y(n_824) );
BUFx12f_ASAP7_75t_L g825 ( .A(n_783), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_685), .B(n_714), .Y(n_826) );
A2O1A1Ixp33_ASAP7_75t_L g827 ( .A1(n_744), .A2(n_696), .B(n_691), .C(n_670), .Y(n_827) );
AND2x4_ASAP7_75t_L g828 ( .A(n_758), .B(n_747), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_698), .Y(n_829) );
CKINVDCx5p33_ASAP7_75t_R g830 ( .A(n_692), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_749), .Y(n_831) );
AO21x2_ASAP7_75t_L g832 ( .A1(n_765), .A2(n_674), .B(n_705), .Y(n_832) );
OAI21xp5_ASAP7_75t_L g833 ( .A1(n_724), .A2(n_735), .B(n_709), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_791), .B(n_757), .Y(n_834) );
OAI221xp5_ASAP7_75t_L g835 ( .A1(n_693), .A2(n_695), .B1(n_677), .B2(n_681), .C(n_672), .Y(n_835) );
OAI21x1_ASAP7_75t_L g836 ( .A1(n_778), .A2(n_713), .B(n_731), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_759), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_684), .Y(n_838) );
AO21x2_ASAP7_75t_L g839 ( .A1(n_679), .A2(n_694), .B(n_732), .Y(n_839) );
OAI21x1_ASAP7_75t_L g840 ( .A1(n_778), .A2(n_733), .B(n_741), .Y(n_840) );
BUFx4f_ASAP7_75t_SL g841 ( .A(n_759), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_706), .B(n_720), .Y(n_842) );
BUFx2_ASAP7_75t_L g843 ( .A(n_755), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_740), .A2(n_716), .B1(n_762), .B2(n_686), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_690), .Y(n_845) );
BUFx6f_ASAP7_75t_L g846 ( .A(n_704), .Y(n_846) );
AOI21x1_ASAP7_75t_L g847 ( .A1(n_761), .A2(n_739), .B(n_682), .Y(n_847) );
OA21x2_ASAP7_75t_L g848 ( .A1(n_712), .A2(n_721), .B(n_763), .Y(n_848) );
CKINVDCx14_ASAP7_75t_R g849 ( .A(n_728), .Y(n_849) );
AOI21xp5_ASAP7_75t_L g850 ( .A1(n_737), .A2(n_734), .B(n_716), .Y(n_850) );
AOI221xp5_ASAP7_75t_L g851 ( .A1(n_710), .A2(n_726), .B1(n_740), .B2(n_762), .C(n_704), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_704), .B(n_771), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_791), .B(n_699), .Y(n_853) );
OAI21x1_ASAP7_75t_L g854 ( .A1(n_771), .A2(n_699), .B(n_791), .Y(n_854) );
OAI211xp5_ASAP7_75t_L g855 ( .A1(n_762), .A2(n_729), .B(n_730), .C(n_727), .Y(n_855) );
BUFx2_ASAP7_75t_L g856 ( .A(n_771), .Y(n_856) );
BUFx3_ASAP7_75t_L g857 ( .A(n_699), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_730), .Y(n_858) );
AOI221xp5_ASAP7_75t_L g859 ( .A1(n_729), .A2(n_467), .B1(n_496), .B2(n_505), .C(n_775), .Y(n_859) );
OAI211xp5_ASAP7_75t_L g860 ( .A1(n_703), .A2(n_675), .B(n_775), .C(n_693), .Y(n_860) );
BUFx3_ASAP7_75t_L g861 ( .A(n_699), .Y(n_861) );
INVx2_ASAP7_75t_L g862 ( .A(n_727), .Y(n_862) );
BUFx2_ASAP7_75t_L g863 ( .A(n_789), .Y(n_863) );
INVx2_ASAP7_75t_L g864 ( .A(n_683), .Y(n_864) );
OAI21xp5_ASAP7_75t_L g865 ( .A1(n_786), .A2(n_781), .B(n_774), .Y(n_865) );
NOR2x1_ASAP7_75t_L g866 ( .A(n_689), .B(n_770), .Y(n_866) );
INVx1_ASAP7_75t_SL g867 ( .A(n_789), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_743), .B(n_568), .Y(n_868) );
A2O1A1Ixp33_ASAP7_75t_L g869 ( .A1(n_742), .A2(n_780), .B(n_772), .C(n_745), .Y(n_869) );
INVxp67_ASAP7_75t_L g870 ( .A(n_789), .Y(n_870) );
NAND2x1p5_ASAP7_75t_L g871 ( .A(n_758), .B(n_474), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_743), .B(n_568), .Y(n_872) );
INVxp67_ASAP7_75t_L g873 ( .A(n_789), .Y(n_873) );
BUFx4f_ASAP7_75t_SL g874 ( .A(n_689), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_782), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_782), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_743), .B(n_568), .Y(n_877) );
BUFx8_ASAP7_75t_L g878 ( .A(n_689), .Y(n_878) );
AO31x2_ASAP7_75t_L g879 ( .A1(n_766), .A2(n_754), .A3(n_539), .B(n_548), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_743), .B(n_568), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_743), .B(n_568), .Y(n_881) );
AO21x2_ASAP7_75t_L g882 ( .A1(n_766), .A2(n_786), .B(n_777), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_782), .Y(n_883) );
OR2x6_ASAP7_75t_L g884 ( .A(n_758), .B(n_573), .Y(n_884) );
OAI21xp5_ASAP7_75t_L g885 ( .A1(n_786), .A2(n_781), .B(n_774), .Y(n_885) );
AND2x2_ASAP7_75t_L g886 ( .A(n_789), .B(n_505), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_683), .Y(n_887) );
OR2x6_ASAP7_75t_L g888 ( .A(n_758), .B(n_573), .Y(n_888) );
A2O1A1Ixp33_ASAP7_75t_L g889 ( .A1(n_742), .A2(n_780), .B(n_772), .C(n_745), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_782), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_683), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_743), .B(n_568), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_743), .B(n_568), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_782), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_789), .B(n_505), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_743), .B(n_568), .Y(n_896) );
INVxp67_ASAP7_75t_SL g897 ( .A(n_789), .Y(n_897) );
OR2x2_ASAP7_75t_L g898 ( .A(n_811), .B(n_795), .Y(n_898) );
INVxp67_ASAP7_75t_SL g899 ( .A(n_897), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_811), .B(n_864), .Y(n_900) );
AOI22xp5_ASAP7_75t_L g901 ( .A1(n_808), .A2(n_859), .B1(n_838), .B2(n_849), .Y(n_901) );
OR2x6_ASAP7_75t_L g902 ( .A(n_808), .B(n_884), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_799), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_887), .B(n_891), .Y(n_904) );
HB1xp67_ASAP7_75t_L g905 ( .A(n_867), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_799), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_834), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_834), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_875), .B(n_876), .Y(n_909) );
NAND3xp33_ASAP7_75t_L g910 ( .A(n_812), .B(n_869), .C(n_889), .Y(n_910) );
BUFx2_ASAP7_75t_L g911 ( .A(n_808), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_883), .B(n_890), .Y(n_912) );
AOI33xp33_ASAP7_75t_L g913 ( .A1(n_867), .A2(n_894), .A3(n_796), .B1(n_817), .B2(n_895), .B3(n_886), .Y(n_913) );
OR2x6_ASAP7_75t_L g914 ( .A(n_884), .B(n_888), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_831), .B(n_819), .Y(n_915) );
OR2x6_ASAP7_75t_L g916 ( .A(n_884), .B(n_888), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_802), .B(n_805), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_810), .B(n_795), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_829), .Y(n_919) );
OA21x2_ASAP7_75t_L g920 ( .A1(n_801), .A2(n_865), .B(n_885), .Y(n_920) );
AND2x2_ASAP7_75t_L g921 ( .A(n_807), .B(n_803), .Y(n_921) );
INVx2_ASAP7_75t_SL g922 ( .A(n_822), .Y(n_922) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_835), .A2(n_870), .B1(n_873), .B2(n_845), .C(n_815), .Y(n_923) );
HB1xp67_ASAP7_75t_L g924 ( .A(n_863), .Y(n_924) );
OAI211xp5_ASAP7_75t_L g925 ( .A1(n_860), .A2(n_824), .B(n_835), .C(n_827), .Y(n_925) );
NAND3xp33_ASAP7_75t_L g926 ( .A(n_865), .B(n_885), .C(n_855), .Y(n_926) );
BUFx3_ASAP7_75t_L g927 ( .A(n_846), .Y(n_927) );
BUFx2_ASAP7_75t_L g928 ( .A(n_888), .Y(n_928) );
AOI221xp5_ASAP7_75t_L g929 ( .A1(n_868), .A2(n_896), .B1(n_893), .B2(n_872), .C(n_892), .Y(n_929) );
HB1xp67_ASAP7_75t_L g930 ( .A(n_803), .Y(n_930) );
AOI21xp5_ASAP7_75t_SL g931 ( .A1(n_844), .A2(n_851), .B(n_842), .Y(n_931) );
INVx2_ASAP7_75t_L g932 ( .A(n_882), .Y(n_932) );
INVx2_ASAP7_75t_L g933 ( .A(n_882), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_868), .Y(n_934) );
BUFx6f_ASAP7_75t_L g935 ( .A(n_854), .Y(n_935) );
BUFx3_ASAP7_75t_L g936 ( .A(n_841), .Y(n_936) );
AOI31xp33_ASAP7_75t_L g937 ( .A1(n_809), .A2(n_844), .A3(n_828), .B(n_871), .Y(n_937) );
INVx2_ASAP7_75t_SL g938 ( .A(n_806), .Y(n_938) );
HB1xp67_ASAP7_75t_L g939 ( .A(n_814), .Y(n_939) );
BUFx2_ASAP7_75t_L g940 ( .A(n_856), .Y(n_940) );
AO21x2_ASAP7_75t_L g941 ( .A1(n_862), .A2(n_858), .B(n_821), .Y(n_941) );
OAI221xp5_ASAP7_75t_L g942 ( .A1(n_818), .A2(n_893), .B1(n_892), .B2(n_881), .C(n_880), .Y(n_942) );
HB1xp67_ASAP7_75t_L g943 ( .A(n_823), .Y(n_943) );
AND2x2_ASAP7_75t_L g944 ( .A(n_872), .B(n_896), .Y(n_944) );
INVx2_ASAP7_75t_L g945 ( .A(n_879), .Y(n_945) );
AO21x2_ASAP7_75t_L g946 ( .A1(n_847), .A2(n_853), .B(n_832), .Y(n_946) );
INVxp33_ASAP7_75t_L g947 ( .A(n_866), .Y(n_947) );
INVx2_ASAP7_75t_L g948 ( .A(n_879), .Y(n_948) );
OAI21xp5_ASAP7_75t_SL g949 ( .A1(n_871), .A2(n_828), .B(n_880), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_881), .B(n_877), .Y(n_950) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_797), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_877), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_826), .Y(n_953) );
AO21x2_ASAP7_75t_L g954 ( .A1(n_832), .A2(n_820), .B(n_833), .Y(n_954) );
INVx2_ASAP7_75t_L g955 ( .A(n_879), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_826), .B(n_837), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_816), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_816), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_852), .B(n_833), .Y(n_959) );
AOI21xp5_ASAP7_75t_SL g960 ( .A1(n_857), .A2(n_861), .B(n_850), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_816), .Y(n_961) );
HB1xp67_ASAP7_75t_L g962 ( .A(n_804), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_848), .B(n_843), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_839), .A2(n_878), .B1(n_874), .B2(n_830), .Y(n_964) );
AOI221xp5_ASAP7_75t_L g965 ( .A1(n_800), .A2(n_878), .B1(n_825), .B2(n_836), .C(n_840), .Y(n_965) );
INVxp67_ASAP7_75t_L g966 ( .A(n_813), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_799), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_811), .B(n_864), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_811), .B(n_864), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_798), .B(n_505), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_799), .Y(n_971) );
AOI22xp5_ASAP7_75t_L g972 ( .A1(n_923), .A2(n_929), .B1(n_950), .B2(n_944), .Y(n_972) );
BUFx3_ASAP7_75t_L g973 ( .A(n_927), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_919), .Y(n_974) );
INVxp67_ASAP7_75t_L g975 ( .A(n_922), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_921), .B(n_959), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_919), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_921), .B(n_959), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_944), .B(n_950), .Y(n_979) );
AND2x2_ASAP7_75t_L g980 ( .A(n_907), .B(n_908), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_934), .B(n_952), .Y(n_981) );
BUFx2_ASAP7_75t_L g982 ( .A(n_902), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_907), .B(n_908), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_956), .B(n_900), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_956), .B(n_900), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_968), .B(n_969), .Y(n_986) );
OR2x2_ASAP7_75t_L g987 ( .A(n_898), .B(n_930), .Y(n_987) );
OR2x2_ASAP7_75t_L g988 ( .A(n_898), .B(n_899), .Y(n_988) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_922), .Y(n_989) );
AND2x4_ASAP7_75t_L g990 ( .A(n_963), .B(n_926), .Y(n_990) );
BUFx2_ASAP7_75t_L g991 ( .A(n_902), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_917), .B(n_963), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_903), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_903), .Y(n_994) );
BUFx3_ASAP7_75t_L g995 ( .A(n_927), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_906), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_967), .Y(n_997) );
OR2x2_ASAP7_75t_L g998 ( .A(n_905), .B(n_971), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_917), .B(n_971), .Y(n_999) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_904), .B(n_920), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_904), .B(n_920), .Y(n_1001) );
BUFx2_ASAP7_75t_SL g1002 ( .A(n_936), .Y(n_1002) );
INVx2_ASAP7_75t_L g1003 ( .A(n_920), .Y(n_1003) );
OR2x2_ASAP7_75t_L g1004 ( .A(n_918), .B(n_953), .Y(n_1004) );
INVx2_ASAP7_75t_L g1005 ( .A(n_932), .Y(n_1005) );
INVx3_ASAP7_75t_SL g1006 ( .A(n_902), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_953), .B(n_942), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_915), .B(n_954), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_910), .B(n_901), .Y(n_1009) );
AND2x4_ASAP7_75t_L g1010 ( .A(n_902), .B(n_945), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_954), .B(n_945), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_954), .B(n_948), .Y(n_1012) );
INVx1_ASAP7_75t_SL g1013 ( .A(n_940), .Y(n_1013) );
OR2x2_ASAP7_75t_L g1014 ( .A(n_943), .B(n_939), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_910), .B(n_901), .Y(n_1015) );
OR2x2_ASAP7_75t_L g1016 ( .A(n_924), .B(n_937), .Y(n_1016) );
INVx2_ASAP7_75t_L g1017 ( .A(n_1005), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_974), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_972), .A2(n_937), .B1(n_902), .B2(n_949), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_977), .Y(n_1020) );
AND2x4_ASAP7_75t_L g1021 ( .A(n_1000), .B(n_935), .Y(n_1021) );
NOR2x1_ASAP7_75t_L g1022 ( .A(n_1002), .B(n_949), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_980), .B(n_913), .Y(n_1023) );
OR2x2_ASAP7_75t_L g1024 ( .A(n_992), .B(n_955), .Y(n_1024) );
OR2x2_ASAP7_75t_L g1025 ( .A(n_992), .B(n_955), .Y(n_1025) );
AND2x4_ASAP7_75t_L g1026 ( .A(n_1000), .B(n_935), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_1001), .B(n_961), .Y(n_1027) );
INVx1_ASAP7_75t_SL g1028 ( .A(n_1013), .Y(n_1028) );
INVx1_ASAP7_75t_SL g1029 ( .A(n_1013), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_1001), .B(n_961), .Y(n_1030) );
OR2x2_ASAP7_75t_L g1031 ( .A(n_1008), .B(n_957), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_986), .B(n_958), .Y(n_1032) );
NAND2x1p5_ASAP7_75t_L g1033 ( .A(n_973), .B(n_911), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_986), .B(n_958), .Y(n_1034) );
NAND4xp25_ASAP7_75t_L g1035 ( .A(n_972), .B(n_925), .C(n_964), .D(n_931), .Y(n_1035) );
BUFx3_ASAP7_75t_L g1036 ( .A(n_973), .Y(n_1036) );
INVx2_ASAP7_75t_SL g1037 ( .A(n_973), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_983), .B(n_931), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_983), .B(n_909), .Y(n_1039) );
INVx2_ASAP7_75t_SL g1040 ( .A(n_995), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_976), .B(n_933), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_978), .B(n_933), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_978), .B(n_946), .Y(n_1043) );
OR2x2_ASAP7_75t_L g1044 ( .A(n_988), .B(n_966), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_984), .B(n_946), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_993), .B(n_912), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_984), .B(n_946), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_985), .B(n_946), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_985), .B(n_941), .Y(n_1049) );
BUFx4f_ASAP7_75t_L g1050 ( .A(n_1006), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_993), .B(n_965), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_979), .B(n_941), .Y(n_1052) );
INVx2_ASAP7_75t_SL g1053 ( .A(n_1036), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1043), .B(n_990), .Y(n_1054) );
BUFx2_ASAP7_75t_L g1055 ( .A(n_1022), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_1023), .B(n_979), .Y(n_1056) );
INVx2_ASAP7_75t_L g1057 ( .A(n_1017), .Y(n_1057) );
OR2x2_ASAP7_75t_L g1058 ( .A(n_1024), .B(n_988), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_1043), .B(n_990), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1018), .Y(n_1060) );
OR2x2_ASAP7_75t_L g1061 ( .A(n_1024), .B(n_987), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_1045), .B(n_990), .Y(n_1062) );
OR2x2_ASAP7_75t_L g1063 ( .A(n_1025), .B(n_1032), .Y(n_1063) );
OR2x2_ASAP7_75t_L g1064 ( .A(n_1025), .B(n_987), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_1045), .B(n_990), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_1047), .B(n_1011), .Y(n_1066) );
INVx1_ASAP7_75t_SL g1067 ( .A(n_1028), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1047), .B(n_1011), .Y(n_1068) );
HB1xp67_ASAP7_75t_L g1069 ( .A(n_1029), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_1048), .B(n_1012), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1020), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1020), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1048), .B(n_1012), .Y(n_1073) );
INVx2_ASAP7_75t_SL g1074 ( .A(n_1036), .Y(n_1074) );
AOI211xp5_ASAP7_75t_L g1075 ( .A1(n_1019), .A2(n_1016), .B(n_1015), .C(n_1009), .Y(n_1075) );
INVx2_ASAP7_75t_SL g1076 ( .A(n_1036), .Y(n_1076) );
NOR3xp33_ASAP7_75t_L g1077 ( .A(n_1035), .B(n_938), .C(n_1015), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_1052), .B(n_1003), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1052), .B(n_1003), .Y(n_1079) );
OR2x6_ASAP7_75t_L g1080 ( .A(n_1022), .B(n_982), .Y(n_1080) );
OR2x2_ASAP7_75t_L g1081 ( .A(n_1032), .B(n_1014), .Y(n_1081) );
OR2x2_ASAP7_75t_L g1082 ( .A(n_1031), .B(n_1014), .Y(n_1082) );
NAND2xp5_ASAP7_75t_SL g1083 ( .A(n_1019), .B(n_1016), .Y(n_1083) );
OR2x2_ASAP7_75t_L g1084 ( .A(n_1031), .B(n_998), .Y(n_1084) );
OR2x2_ASAP7_75t_L g1085 ( .A(n_1041), .B(n_998), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1039), .B(n_999), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_1049), .B(n_1010), .Y(n_1087) );
AND2x4_ASAP7_75t_L g1088 ( .A(n_1021), .B(n_1010), .Y(n_1088) );
AOI22xp5_ASAP7_75t_L g1089 ( .A1(n_1083), .A2(n_1035), .B1(n_1038), .B2(n_1009), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_1054), .B(n_1049), .Y(n_1090) );
INVxp67_ASAP7_75t_L g1091 ( .A(n_1069), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1060), .Y(n_1092) );
OA21x2_ASAP7_75t_L g1093 ( .A1(n_1055), .A2(n_1038), .B(n_1051), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_1056), .B(n_1034), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1054), .B(n_1041), .Y(n_1095) );
AND2x4_ASAP7_75t_L g1096 ( .A(n_1088), .B(n_1078), .Y(n_1096) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1057), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_1059), .B(n_1042), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_1066), .B(n_1027), .Y(n_1099) );
NAND2xp5_ASAP7_75t_SL g1100 ( .A(n_1055), .B(n_1050), .Y(n_1100) );
AND3x2_ASAP7_75t_L g1101 ( .A(n_1075), .B(n_951), .C(n_962), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1059), .B(n_1042), .Y(n_1102) );
OAI32xp33_ASAP7_75t_L g1103 ( .A1(n_1077), .A2(n_1044), .A3(n_989), .B1(n_975), .B2(n_1029), .Y(n_1103) );
NOR2x1_ASAP7_75t_L g1104 ( .A(n_1080), .B(n_1002), .Y(n_1104) );
AND2x4_ASAP7_75t_L g1105 ( .A(n_1088), .B(n_1021), .Y(n_1105) );
NAND2x1p5_ASAP7_75t_L g1106 ( .A(n_1053), .B(n_1050), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_1068), .B(n_1030), .Y(n_1107) );
INVx2_ASAP7_75t_L g1108 ( .A(n_1060), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1071), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1072), .Y(n_1110) );
INVx2_ASAP7_75t_L g1111 ( .A(n_1097), .Y(n_1111) );
INVx2_ASAP7_75t_L g1112 ( .A(n_1097), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_1089), .A2(n_1007), .B1(n_1051), .B2(n_1044), .Y(n_1113) );
OAI21xp33_ASAP7_75t_L g1114 ( .A1(n_1103), .A2(n_1065), .B(n_1062), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_1093), .B(n_1070), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1093), .B(n_1070), .Y(n_1116) );
OAI21xp5_ASAP7_75t_L g1117 ( .A1(n_1104), .A2(n_1067), .B(n_938), .Y(n_1117) );
OAI322xp33_ASAP7_75t_L g1118 ( .A1(n_1091), .A2(n_1082), .A3(n_1081), .B1(n_1063), .B2(n_1084), .C1(n_1086), .C2(n_1064), .Y(n_1118) );
NAND2x1_ASAP7_75t_L g1119 ( .A(n_1096), .B(n_1080), .Y(n_1119) );
AOI21xp33_ASAP7_75t_L g1120 ( .A1(n_1103), .A2(n_947), .B(n_1007), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g1121 ( .A1(n_1101), .A2(n_1079), .B1(n_1087), .B2(n_1073), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1092), .Y(n_1122) );
AOI211xp5_ASAP7_75t_L g1123 ( .A1(n_1120), .A2(n_1100), .B(n_1006), .C(n_1084), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_1114), .A2(n_982), .B1(n_991), .B2(n_1080), .Y(n_1124) );
AOI221x1_ASAP7_75t_L g1125 ( .A1(n_1117), .A2(n_1110), .B1(n_1109), .B2(n_1096), .C(n_1094), .Y(n_1125) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1122), .Y(n_1126) );
OR2x2_ASAP7_75t_L g1127 ( .A(n_1115), .B(n_1099), .Y(n_1127) );
OAI22xp33_ASAP7_75t_L g1128 ( .A1(n_1119), .A2(n_1106), .B1(n_1074), .B2(n_1076), .Y(n_1128) );
AOI221xp5_ASAP7_75t_L g1129 ( .A1(n_1118), .A2(n_1039), .B1(n_1107), .B2(n_1110), .C(n_1109), .Y(n_1129) );
AOI222xp33_ASAP7_75t_L g1130 ( .A1(n_1113), .A2(n_1090), .B1(n_1095), .B2(n_1102), .C1(n_1098), .C2(n_1096), .Y(n_1130) );
AOI21xp33_ASAP7_75t_L g1131 ( .A1(n_1121), .A2(n_1076), .B(n_1074), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1129), .B(n_1116), .Y(n_1132) );
OAI221xp5_ASAP7_75t_L g1133 ( .A1(n_1129), .A2(n_1124), .B1(n_1131), .B2(n_1123), .C(n_1130), .Y(n_1133) );
OAI322xp33_ASAP7_75t_L g1134 ( .A1(n_1128), .A2(n_1061), .A3(n_1058), .B1(n_1085), .B2(n_1111), .C1(n_1112), .C2(n_1004), .Y(n_1134) );
OAI211xp5_ASAP7_75t_L g1135 ( .A1(n_1125), .A2(n_936), .B(n_928), .C(n_911), .Y(n_1135) );
OAI211xp5_ASAP7_75t_SL g1136 ( .A1(n_1127), .A2(n_1111), .B(n_1046), .C(n_1037), .Y(n_1136) );
OAI221xp5_ASAP7_75t_L g1137 ( .A1(n_1126), .A2(n_1106), .B1(n_991), .B2(n_1006), .C(n_1108), .Y(n_1137) );
OAI221xp5_ASAP7_75t_L g1138 ( .A1(n_1133), .A2(n_1050), .B1(n_916), .B2(n_914), .C(n_1033), .Y(n_1138) );
NAND5xp2_ASAP7_75t_L g1139 ( .A(n_1135), .B(n_1033), .C(n_970), .D(n_996), .E(n_997), .Y(n_1139) );
AOI221xp5_ASAP7_75t_L g1140 ( .A1(n_1134), .A2(n_1090), .B1(n_1098), .B2(n_1095), .C(n_1102), .Y(n_1140) );
OAI211xp5_ASAP7_75t_L g1141 ( .A1(n_1132), .A2(n_960), .B(n_1040), .C(n_1037), .Y(n_1141) );
NOR3xp33_ASAP7_75t_L g1142 ( .A(n_1138), .B(n_1137), .C(n_1136), .Y(n_1142) );
NAND3xp33_ASAP7_75t_SL g1143 ( .A(n_1141), .B(n_1033), .C(n_940), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1142), .B(n_1140), .Y(n_1144) );
OR3x1_ASAP7_75t_L g1145 ( .A(n_1143), .B(n_1139), .C(n_994), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1144), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1145), .Y(n_1147) );
XNOR2xp5_ASAP7_75t_L g1148 ( .A(n_1147), .B(n_914), .Y(n_1148) );
OAI22xp5_ASAP7_75t_SL g1149 ( .A1(n_1148), .A2(n_1146), .B1(n_914), .B2(n_916), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1149), .Y(n_1150) );
OAI21xp5_ASAP7_75t_L g1151 ( .A1(n_1150), .A2(n_1105), .B(n_981), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_1151), .A2(n_1088), .B1(n_1021), .B2(n_1026), .Y(n_1152) );
endmodule