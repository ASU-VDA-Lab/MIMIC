module fake_jpeg_6521_n_308 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_308);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_30),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_34),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_25),
.B1(n_13),
.B2(n_27),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_40),
.B1(n_13),
.B2(n_25),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_27),
.B1(n_13),
.B2(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_57),
.Y(n_77)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_34),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_71),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_65),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_60),
.A2(n_74),
.B1(n_13),
.B2(n_29),
.Y(n_87)
);

CKINVDCx12_ASAP7_75t_R g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_35),
.Y(n_65)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_72),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_34),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_43),
.B(n_30),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_39),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_13),
.B1(n_27),
.B2(n_29),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_79),
.Y(n_99)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_80),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_75),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_48),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_91),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_16),
.B1(n_27),
.B2(n_69),
.Y(n_118)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_93),
.Y(n_117)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_67),
.Y(n_104)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_41),
.C(n_35),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_58),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_103),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_38),
.C(n_61),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_61),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_115),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_45),
.C(n_70),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_42),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_94),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_52),
.Y(n_116)
);

XNOR2x1_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_85),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_119),
.B1(n_77),
.B2(n_79),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_47),
.B1(n_44),
.B2(n_51),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_122),
.B(n_125),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_100),
.B(n_92),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_137),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_130),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVxp33_ASAP7_75t_SL g145 ( 
.A(n_129),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_133),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_132),
.A2(n_136),
.B(n_139),
.Y(n_147)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_134),
.A2(n_135),
.B1(n_142),
.B2(n_115),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_116),
.A2(n_92),
.B1(n_76),
.B2(n_16),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_23),
.B(n_26),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_100),
.B(n_30),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_140),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_31),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_103),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_102),
.B1(n_101),
.B2(n_98),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_143),
.B1(n_119),
.B2(n_109),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_16),
.B1(n_69),
.B2(n_89),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_112),
.A2(n_93),
.B(n_80),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_144),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_152),
.Y(n_188)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_135),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_156),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_170),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_130),
.B(n_108),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_159),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_131),
.B(n_105),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_132),
.A2(n_140),
.B1(n_128),
.B2(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_161),
.B(n_163),
.Y(n_185)
);

OAI32xp33_ASAP7_75t_L g162 ( 
.A1(n_126),
.A2(n_105),
.A3(n_22),
.B1(n_36),
.B2(n_31),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_168),
.Y(n_173)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_164),
.B(n_167),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_128),
.A2(n_78),
.B1(n_97),
.B2(n_31),
.Y(n_165)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_136),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_139),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_126),
.A2(n_90),
.B(n_37),
.Y(n_170)
);

NOR4xp25_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_90),
.C(n_52),
.D(n_45),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_143),
.C(n_139),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_167),
.B(n_122),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_172),
.B(n_190),
.Y(n_206)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_181),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_141),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_147),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_133),
.Y(n_180)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_120),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_182),
.A2(n_147),
.B1(n_150),
.B2(n_148),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_120),
.C(n_135),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_156),
.C(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_187),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_136),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_193),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_154),
.B(n_95),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_24),
.B(n_15),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_139),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_194),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_163),
.B(n_95),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_142),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_197),
.B(n_210),
.Y(n_237)
);

XNOR2x1_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_152),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_198),
.B(n_199),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_168),
.B1(n_165),
.B2(n_123),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_204),
.B1(n_207),
.B2(n_212),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_202),
.C(n_216),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_145),
.C(n_162),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_159),
.B1(n_157),
.B2(n_169),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_175),
.A2(n_161),
.B1(n_106),
.B2(n_18),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_106),
.Y(n_208)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_208),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_90),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_106),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_211),
.B(n_217),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_19),
.B1(n_23),
.B2(n_26),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_194),
.B1(n_187),
.B2(n_196),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_52),
.C(n_45),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_186),
.B(n_19),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_36),
.C(n_56),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_185),
.C(n_192),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_177),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_227),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_176),
.Y(n_221)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_178),
.Y(n_224)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_228),
.C(n_231),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_226),
.B(n_233),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_177),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_180),
.C(n_173),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_189),
.B1(n_173),
.B2(n_19),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_230),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_189),
.C(n_36),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_218),
.B(n_15),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_200),
.A2(n_26),
.B1(n_23),
.B2(n_15),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_219),
.B1(n_236),
.B2(n_14),
.Y(n_250)
);

INVx4_ASAP7_75t_SL g235 ( 
.A(n_214),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_235),
.A2(n_225),
.B(n_231),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_56),
.C(n_17),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_209),
.C(n_207),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_202),
.A2(n_14),
.B1(n_26),
.B2(n_22),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_238),
.B(n_12),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_SL g241 ( 
.A1(n_235),
.A2(n_205),
.B(n_214),
.C(n_215),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_251),
.B1(n_0),
.B2(n_1),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_245),
.B(n_248),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_228),
.B(n_214),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_246),
.B(n_2),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_213),
.Y(n_248)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_20),
.A3(n_14),
.B1(n_12),
.B2(n_17),
.C1(n_24),
.C2(n_56),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_17),
.C(n_21),
.Y(n_268)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_223),
.A2(n_24),
.B(n_22),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_255),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_17),
.C(n_20),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_17),
.C(n_21),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_229),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_255),
.B(n_229),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_257),
.C(n_262),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_237),
.Y(n_257)
);

FAx1_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_0),
.CI(n_1),
.CON(n_258),
.SN(n_258)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_258),
.A2(n_263),
.B(n_268),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_241),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_259)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_17),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_17),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_3),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_250),
.C(n_251),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_243),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_3),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_17),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_21),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_253),
.Y(n_273)
);

NOR2x1p5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_258),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_261),
.B(n_244),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_276),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_266),
.A2(n_241),
.B1(n_247),
.B2(n_239),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_275),
.B(n_279),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_254),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_265),
.C(n_257),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_256),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_282),
.B(n_277),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_288),
.B(n_291),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_280),
.C(n_273),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_287),
.B(n_289),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g298 ( 
.A1(n_290),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_276),
.B(n_267),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_281),
.B(n_270),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_296),
.A2(n_297),
.B(n_298),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_3),
.B(n_4),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_295),
.A2(n_283),
.B(n_284),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_21),
.C(n_9),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_299),
.A2(n_294),
.A3(n_21),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_7),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_302),
.A2(n_303),
.B(n_300),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_6),
.C(n_9),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_6),
.B(n_11),
.Y(n_306)
);

OAI211xp5_ASAP7_75t_SL g307 ( 
.A1(n_306),
.A2(n_6),
.B(n_11),
.C(n_21),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_11),
.C(n_21),
.Y(n_308)
);


endmodule