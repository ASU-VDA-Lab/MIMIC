module fake_jpeg_17855_n_162 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_162);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_11),
.B(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_37),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_33),
.A2(n_35),
.B1(n_38),
.B2(n_25),
.Y(n_68)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx2_ASAP7_75t_SL g64 ( 
.A(n_34),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_3),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_R g53 ( 
.A(n_36),
.B(n_30),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_31),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_5),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_6),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_42),
.A2(n_43),
.B(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_7),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_46),
.Y(n_51)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_50),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_62),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_54),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_32),
.Y(n_54)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_61),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_19),
.C(n_20),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_60),
.B(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_21),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_33),
.B1(n_44),
.B2(n_38),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_25),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_43),
.B(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_11),
.Y(n_73)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_19),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_34),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_26),
.B1(n_27),
.B2(n_20),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_67),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_86),
.B1(n_94),
.B2(n_98),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_39),
.B(n_19),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_85),
.C(n_91),
.Y(n_101)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_52),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_20),
.B(n_46),
.Y(n_85)
);

OA21x2_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_24),
.B(n_26),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_59),
.B(n_75),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_74),
.B(n_71),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_12),
.B1(n_57),
.B2(n_72),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_67),
.B(n_58),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_55),
.C(n_54),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_98),
.A2(n_77),
.B1(n_62),
.B2(n_71),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_69),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_105),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_69),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_84),
.A2(n_66),
.B(n_51),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_108),
.B1(n_80),
.B2(n_94),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_91),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_57),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_118),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_52),
.C(n_56),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_113),
.C(n_116),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_52),
.C(n_56),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_85),
.C(n_82),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_87),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_126),
.B1(n_97),
.B2(n_86),
.Y(n_136)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

BUFx24_ASAP7_75t_SL g127 ( 
.A(n_109),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_132),
.C(n_79),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_130),
.B(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_87),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_101),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_138),
.C(n_139),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_101),
.C(n_116),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_135),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_113),
.B(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_136),
.B(n_137),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_108),
.B1(n_86),
.B2(n_88),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_88),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g140 ( 
.A(n_124),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_83),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_97),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_131),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_148),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_147),
.C(n_123),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_119),
.Y(n_148)
);

AOI221xp5_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_125),
.B1(n_134),
.B2(n_138),
.C(n_120),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_150),
.B(n_151),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_133),
.C(n_139),
.Y(n_152)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

OAI21x1_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_146),
.B(n_128),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_100),
.Y(n_156)
);

OAI31xp33_ASAP7_75t_L g159 ( 
.A1(n_156),
.A2(n_100),
.A3(n_150),
.B(n_155),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_156),
.B(n_154),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_158),
.B(n_157),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_159),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_161),
.Y(n_162)
);


endmodule