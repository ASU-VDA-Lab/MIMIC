module fake_jpeg_26387_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_36),
.Y(n_52)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_38),
.Y(n_54)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_29),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_26),
.B1(n_20),
.B2(n_24),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_43),
.A2(n_50),
.B1(n_53),
.B2(n_16),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_32),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_45),
.C(n_55),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_26),
.B1(n_20),
.B2(n_28),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_48),
.B1(n_16),
.B2(n_28),
.Y(n_78)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_25),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_22),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_57),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_26),
.B1(n_20),
.B2(n_27),
.Y(n_50)
);

HAxp5_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_27),
.CON(n_51),
.SN(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_51),
.A2(n_56),
.B(n_49),
.C(n_21),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_33),
.B1(n_38),
.B2(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_69),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_61),
.Y(n_113)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_71),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_75),
.B(n_21),
.C(n_29),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_18),
.Y(n_65)
);

BUFx24_ASAP7_75t_SL g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_67),
.Y(n_92)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_22),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_22),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_22),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_34),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_38),
.B1(n_17),
.B2(n_22),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_81),
.B1(n_82),
.B2(n_48),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_23),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_39),
.Y(n_100)
);

OAI22x1_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_25),
.B1(n_30),
.B2(n_32),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_17),
.B1(n_22),
.B2(n_30),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_43),
.B1(n_50),
.B2(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_31),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_31),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_25),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_44),
.A2(n_18),
.B1(n_21),
.B2(n_28),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_64),
.B(n_70),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_42),
.B(n_39),
.C(n_55),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_55),
.Y(n_105)
);

NOR2x1_ASAP7_75t_R g122 ( 
.A(n_88),
.B(n_69),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_105),
.B(n_107),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_62),
.B(n_42),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_102),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_17),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_111),
.B(n_59),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_17),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_114),
.A2(n_113),
.B1(n_102),
.B2(n_99),
.Y(n_138)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_115),
.B(n_117),
.Y(n_153)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_118),
.B(n_124),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_121),
.A2(n_122),
.B(n_139),
.Y(n_152)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_131),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_58),
.C(n_72),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_129),
.C(n_112),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_114),
.A2(n_63),
.B1(n_59),
.B2(n_82),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_134),
.B1(n_138),
.B2(n_140),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_75),
.C(n_73),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_75),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_135),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_93),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_141),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_114),
.A2(n_68),
.B1(n_83),
.B2(n_74),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_55),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_101),
.B(n_61),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_96),
.A2(n_30),
.B1(n_0),
.B2(n_1),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_147),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_111),
.B1(n_96),
.B2(n_117),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_155),
.B(n_158),
.Y(n_173)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_156),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_89),
.B1(n_107),
.B2(n_109),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_157),
.B1(n_164),
.B2(n_166),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_138),
.A2(n_88),
.B(n_90),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_94),
.C(n_90),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_120),
.A2(n_92),
.B1(n_98),
.B2(n_108),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_116),
.A2(n_113),
.B(n_1),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_122),
.A2(n_92),
.B(n_113),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_170),
.B(n_125),
.Y(n_185)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_161),
.Y(n_188)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_110),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_162),
.B(n_169),
.Y(n_179)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_163),
.B(n_165),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_124),
.A2(n_110),
.B1(n_79),
.B2(n_3),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_123),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_116),
.A2(n_79),
.B1(n_2),
.B2(n_3),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_137),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_168),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_118),
.B(n_79),
.C(n_2),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_121),
.A2(n_0),
.B(n_3),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_172),
.B(n_175),
.Y(n_208)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

XNOR2x1_ASAP7_75t_SL g176 ( 
.A(n_152),
.B(n_132),
.Y(n_176)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_176),
.B(n_179),
.CI(n_151),
.CON(n_196),
.SN(n_196)
);

OAI322xp33_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_125),
.A3(n_136),
.B1(n_131),
.B2(n_126),
.C1(n_133),
.C2(n_130),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_159),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_160),
.B(n_130),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_178),
.B(n_189),
.Y(n_202)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_184),
.Y(n_209)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_185),
.A2(n_192),
.B1(n_170),
.B2(n_169),
.Y(n_211)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_163),
.B(n_11),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_142),
.Y(n_190)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_146),
.A2(n_15),
.B1(n_5),
.B2(n_6),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_193),
.A2(n_167),
.B1(n_161),
.B2(n_147),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_149),
.B(n_11),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_143),
.B1(n_9),
.B2(n_10),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_154),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_201),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_199),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_162),
.C(n_148),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_156),
.C(n_150),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_203),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_152),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_188),
.B1(n_195),
.B2(n_185),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_144),
.C(n_158),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_214),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_173),
.Y(n_210)
);

BUFx24_ASAP7_75t_SL g227 ( 
.A(n_210),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_211),
.A2(n_213),
.B1(n_193),
.B2(n_183),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_184),
.A2(n_155),
.B1(n_143),
.B2(n_0),
.Y(n_213)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_217),
.B(n_219),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_183),
.B1(n_175),
.B2(n_172),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

BUFx12_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_221),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_173),
.B(n_188),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_222),
.A2(n_225),
.B(n_229),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_202),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_224),
.Y(n_238)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_205),
.Y(n_231)
);

OAI22x1_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_180),
.B1(n_186),
.B2(n_182),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_199),
.C(n_200),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_236),
.C(n_240),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_235),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_206),
.C(n_203),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_210),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_240),
.Y(n_243)
);

XOR2x2_ASAP7_75t_SL g239 ( 
.A(n_229),
.B(n_201),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_196),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_196),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_244),
.C(n_251),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_227),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_238),
.A2(n_198),
.B1(n_180),
.B2(n_219),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_246),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_234),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_248),
.Y(n_255)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_233),
.A2(n_224),
.B1(n_218),
.B2(n_212),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_250),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_230),
.C(n_236),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_257),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_231),
.C(n_221),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_221),
.C(n_239),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_189),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_243),
.C(n_251),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_261),
.C(n_12),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_248),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_263),
.B(n_194),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_182),
.C(n_191),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_267),
.B(n_13),
.Y(n_269)
);

AOI322xp5_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_255),
.A3(n_9),
.B1(n_10),
.B2(n_12),
.C1(n_7),
.C2(n_14),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_SL g268 ( 
.A(n_265),
.B(n_266),
.Y(n_268)
);

AOI21x1_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_7),
.B(n_12),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_13),
.B(n_15),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_268),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_13),
.Y(n_272)
);


endmodule