module fake_netlist_6_4891_n_192 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_2, n_5, n_19, n_25, n_192);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;
input n_25;

output n_192;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_191;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_87;
wire n_189;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_29;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_108;
wire n_94;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_190;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_30;
wire n_79;
wire n_43;
wire n_171;
wire n_31;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVxp33_ASAP7_75t_SL g32 ( 
.A(n_16),
.Y(n_32)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVxp67_ASAP7_75t_SL g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_R g62 ( 
.A(n_42),
.B(n_21),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_29),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_29),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_39),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

AND2x4_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_45),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

NAND2x1p5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

NAND2x1_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_50),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_47),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_66),
.B1(n_70),
.B2(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_38),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_35),
.B(n_37),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_56),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_63),
.B1(n_57),
.B2(n_33),
.Y(n_91)
);

OAI321xp33_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_40),
.A3(n_41),
.B1(n_47),
.B2(n_67),
.C(n_69),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_56),
.B1(n_69),
.B2(n_68),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

OAI21x1_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_68),
.B(n_67),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_72),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_71),
.B(n_41),
.C(n_40),
.Y(n_99)
);

AO21x1_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_56),
.B(n_1),
.Y(n_100)
);

OAI21x1_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_77),
.B(n_76),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

OAI21x1_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_80),
.B(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NAND2x1p5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_79),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_78),
.B1(n_60),
.B2(n_88),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_90),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_SL g112 ( 
.A(n_107),
.B(n_90),
.C(n_62),
.Y(n_112)
);

OR2x6_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_96),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_107),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_96),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_110),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_102),
.B(n_105),
.Y(n_120)
);

NOR2x1_ASAP7_75t_SL g121 ( 
.A(n_116),
.B(n_113),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

AND2x4_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_113),
.Y(n_124)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_120),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_111),
.Y(n_128)
);

NAND4xp25_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_99),
.C(n_108),
.D(n_89),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_122),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_100),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_128),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_115),
.Y(n_136)
);

AND2x4_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_101),
.B(n_110),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_101),
.B(n_108),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

AOI211xp5_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_129),
.B(n_92),
.C(n_127),
.Y(n_143)
);

AOI322xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_130),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_6),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_130),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_138),
.A2(n_131),
.B1(n_113),
.B2(n_106),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_78),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_139),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

OAI211xp5_ASAP7_75t_SL g157 ( 
.A1(n_152),
.A2(n_144),
.B(n_141),
.C(n_132),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_154),
.B1(n_153),
.B2(n_155),
.Y(n_158)
);

AOI211xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_92),
.B(n_137),
.C(n_136),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_137),
.Y(n_160)
);

AOI221xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_133),
.B1(n_74),
.B2(n_75),
.C(n_87),
.Y(n_161)
);

AOI21x1_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_77),
.B(n_103),
.Y(n_162)
);

AOI221xp5_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_133),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_163)
);

OAI321xp33_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_0),
.A3(n_8),
.B1(n_9),
.B2(n_105),
.C(n_94),
.Y(n_164)
);

OAI211xp5_ASAP7_75t_SL g165 ( 
.A1(n_152),
.A2(n_98),
.B(n_94),
.C(n_102),
.Y(n_165)
);

AOI222xp33_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_81),
.B1(n_73),
.B2(n_96),
.C1(n_94),
.C2(n_23),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_73),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_160),
.Y(n_168)
);

XOR2x2_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_11),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_102),
.B1(n_81),
.B2(n_73),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_73),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_168),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_171),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_161),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_R g178 ( 
.A(n_166),
.B(n_18),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_20),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

AOI22x1_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_179),
.B1(n_178),
.B2(n_173),
.Y(n_185)
);

OAI22x1_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_179),
.B1(n_102),
.B2(n_103),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_181),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_185),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_182),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_189),
.A2(n_180),
.B1(n_182),
.B2(n_186),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_190),
.B(n_188),
.Y(n_192)
);


endmodule