module fake_netlist_5_961_n_196 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_30, n_20, n_5, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_196);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;

output n_196;

wire n_137;
wire n_168;
wire n_164;
wire n_191;
wire n_91;
wire n_82;
wire n_122;
wire n_194;
wire n_142;
wire n_176;
wire n_140;
wire n_124;
wire n_146;
wire n_136;
wire n_86;
wire n_182;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_180;
wire n_184;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_189;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_69;
wire n_58;
wire n_116;
wire n_195;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_179;
wire n_125;
wire n_35;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_193;
wire n_131;
wire n_151;
wire n_47;
wire n_173;
wire n_192;
wire n_53;
wire n_160;
wire n_188;
wire n_190;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_154;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_185;
wire n_183;
wire n_175;
wire n_169;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_181;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_178;
wire n_67;
wire n_121;
wire n_76;
wire n_36;
wire n_87;
wire n_150;
wire n_162;
wire n_170;
wire n_77;
wire n_64;
wire n_106;
wire n_102;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_174;
wire n_186;
wire n_134;
wire n_187;
wire n_104;
wire n_41;
wire n_32;
wire n_172;
wire n_103;
wire n_56;
wire n_51;
wire n_97;
wire n_141;
wire n_63;
wire n_166;
wire n_171;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVxp67_ASAP7_75t_SL g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVxp33_ASAP7_75t_SL g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVxp33_ASAP7_75t_SL g54 ( 
.A(n_7),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_1),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_2),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_3),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_7),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_39),
.B1(n_51),
.B2(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

AO22x2_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_51),
.B1(n_53),
.B2(n_38),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

NAND2x1p5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_50),
.Y(n_84)
);

OR2x6_ASAP7_75t_SL g85 ( 
.A(n_76),
.B(n_36),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

AO22x2_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_46),
.B1(n_52),
.B2(n_54),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_66),
.B(n_72),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

OR2x6_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_42),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

CKINVDCx11_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_74),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_69),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_65),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_90),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_72),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_69),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_69),
.Y(n_105)
);

O2A1O1Ixp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_60),
.B(n_73),
.C(n_74),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_101),
.A2(n_92),
.B1(n_32),
.B2(n_70),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_79),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_82),
.Y(n_110)
);

NOR2x2_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_92),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_98),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_64),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_82),
.Y(n_114)
);

NOR2x1_ASAP7_75t_SL g115 ( 
.A(n_112),
.B(n_100),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_98),
.Y(n_116)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_113),
.B(n_109),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_98),
.B(n_97),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

OA21x2_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_97),
.B(n_103),
.Y(n_121)
);

CKINVDCx8_ASAP7_75t_R g122 ( 
.A(n_119),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_109),
.B(n_113),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

OAI21x1_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_117),
.B(n_116),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_99),
.C(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

OA21x2_ASAP7_75t_L g132 ( 
.A1(n_123),
.A2(n_117),
.B(n_74),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_124),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_119),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

AO21x2_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_115),
.B(n_102),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_115),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_87),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_87),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_138),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_128),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_107),
.B1(n_87),
.B2(n_84),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_126),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_129),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_129),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

NAND2x1_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_135),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_130),
.Y(n_157)
);

XOR2x2_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_107),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_130),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_84),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_148),
.C(n_145),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_149),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_136),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_157),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_68),
.B(n_70),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_154),
.Y(n_173)
);

OAI31xp33_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_158),
.A3(n_68),
.B(n_63),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_169),
.A2(n_158),
.B1(n_111),
.B2(n_122),
.Y(n_175)
);

AND4x1_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_63),
.C(n_64),
.D(n_61),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

NAND3x1_ASAP7_75t_SL g178 ( 
.A(n_167),
.B(n_8),
.C(n_9),
.Y(n_178)
);

AND4x1_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_61),
.C(n_58),
.D(n_11),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_58),
.C(n_71),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_60),
.A3(n_8),
.B1(n_10),
.B2(n_12),
.C1(n_55),
.C2(n_71),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_170),
.B1(n_167),
.B2(n_172),
.Y(n_183)
);

AOI22x1_ASAP7_75t_L g184 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_174),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

NAND4xp25_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_60),
.C(n_10),
.D(n_102),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g187 ( 
.A1(n_176),
.A2(n_60),
.A3(n_71),
.B1(n_135),
.B2(n_119),
.C1(n_93),
.C2(n_89),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

AO22x1_ASAP7_75t_SL g189 ( 
.A1(n_184),
.A2(n_176),
.B1(n_135),
.B2(n_83),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_186),
.A2(n_185),
.B1(n_188),
.B2(n_183),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_130),
.B1(n_132),
.B2(n_71),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_71),
.A3(n_119),
.B1(n_86),
.B2(n_81),
.C1(n_132),
.C2(n_29),
.Y(n_192)
);

OAI322xp33_ASAP7_75t_L g193 ( 
.A1(n_190),
.A2(n_119),
.A3(n_103),
.B1(n_132),
.B2(n_25),
.C1(n_28),
.C2(n_19),
.Y(n_193)
);

AOI321xp33_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_191),
.A3(n_192),
.B1(n_103),
.B2(n_14),
.C(n_15),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

AOI221xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_132),
.B1(n_136),
.B2(n_193),
.C(n_190),
.Y(n_196)
);


endmodule