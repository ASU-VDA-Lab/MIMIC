module real_aes_8148_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_500;
wire n_307;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_1), .A2(n_5), .B1(n_465), .B2(n_470), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_2), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_3), .A2(n_35), .B1(n_102), .B2(n_160), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_4), .A2(n_69), .B1(n_482), .B2(n_486), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_6), .B(n_137), .Y(n_145) );
AND2x6_ASAP7_75t_L g117 ( .A(n_7), .B(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g507 ( .A(n_7), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_7), .B(n_514), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_8), .A2(n_391), .B1(n_392), .B2(n_405), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_8), .Y(n_391) );
AO22x2_ASAP7_75t_L g418 ( .A1(n_9), .A2(n_30), .B1(n_415), .B2(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g93 ( .A(n_10), .Y(n_93) );
INVx1_ASAP7_75t_L g96 ( .A(n_11), .Y(n_96) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_12), .B(n_98), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_13), .B(n_89), .Y(n_147) );
AO32x2_ASAP7_75t_L g198 ( .A1(n_14), .A2(n_88), .A3(n_131), .B1(n_137), .B2(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_15), .B(n_102), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_16), .B(n_89), .Y(n_119) );
AO22x2_ASAP7_75t_L g422 ( .A1(n_17), .A2(n_33), .B1(n_415), .B2(n_416), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_18), .A2(n_42), .B1(n_102), .B2(n_160), .Y(n_201) );
AOI22xp33_ASAP7_75t_SL g162 ( .A1(n_19), .A2(n_62), .B1(n_98), .B2(n_102), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_20), .B(n_102), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_21), .A2(n_407), .B1(n_408), .B2(n_495), .Y(n_406) );
INVx1_ASAP7_75t_L g495 ( .A(n_21), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_22), .A2(n_399), .B1(n_402), .B2(n_403), .Y(n_398) );
INVxp67_ASAP7_75t_L g402 ( .A(n_22), .Y(n_402) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_23), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_24), .B(n_133), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_25), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_26), .A2(n_65), .B1(n_490), .B2(n_492), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_27), .B(n_133), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_28), .Y(n_451) );
INVx2_ASAP7_75t_L g100 ( .A(n_29), .Y(n_100) );
NAND2xp5_ASAP7_75t_SL g124 ( .A(n_31), .B(n_102), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_32), .B(n_133), .Y(n_186) );
OAI221xp5_ASAP7_75t_L g499 ( .A1(n_33), .A2(n_47), .B1(n_57), .B2(n_500), .C(n_501), .Y(n_499) );
INVxp67_ASAP7_75t_L g502 ( .A(n_33), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_34), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_36), .A2(n_63), .B1(n_441), .B2(n_445), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_37), .B(n_102), .Y(n_140) );
INVx1_ASAP7_75t_L g520 ( .A(n_37), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_38), .A2(n_71), .B1(n_160), .B2(n_161), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_39), .B(n_102), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_40), .B(n_102), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_41), .B(n_110), .Y(n_144) );
AOI22xp5_ASAP7_75t_SL g509 ( .A1(n_41), .A2(n_407), .B1(n_408), .B2(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_41), .Y(n_510) );
AOI22xp33_ASAP7_75t_SL g151 ( .A1(n_43), .A2(n_49), .B1(n_98), .B2(n_102), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_44), .B(n_102), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_45), .B(n_102), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_46), .A2(n_61), .B1(n_400), .B2(n_401), .Y(n_399) );
CKINVDCx16_ASAP7_75t_R g401 ( .A(n_46), .Y(n_401) );
AO22x2_ASAP7_75t_L g414 ( .A1(n_47), .A2(n_67), .B1(n_415), .B2(n_416), .Y(n_414) );
INVxp67_ASAP7_75t_L g503 ( .A(n_47), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_48), .A2(n_60), .B1(n_475), .B2(n_478), .Y(n_474) );
INVx1_ASAP7_75t_L g118 ( .A(n_50), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_51), .B(n_102), .Y(n_113) );
INVx1_ASAP7_75t_L g92 ( .A(n_52), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_53), .Y(n_500) );
AO32x2_ASAP7_75t_L g157 ( .A1(n_54), .A2(n_131), .A3(n_137), .B1(n_158), .B2(n_163), .Y(n_157) );
INVx1_ASAP7_75t_L g127 ( .A(n_55), .Y(n_127) );
INVx1_ASAP7_75t_L g170 ( .A(n_56), .Y(n_170) );
AO22x2_ASAP7_75t_L g432 ( .A1(n_57), .A2(n_73), .B1(n_415), .B2(n_419), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_58), .B(n_98), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_59), .Y(n_423) );
INVx1_ASAP7_75t_L g400 ( .A(n_61), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_62), .A2(n_395), .B1(n_396), .B2(n_397), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_62), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_64), .B(n_160), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_66), .B(n_98), .Y(n_174) );
INVx2_ASAP7_75t_L g90 ( .A(n_68), .Y(n_90) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_70), .B(n_98), .Y(n_141) );
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_72), .A2(n_77), .B1(n_98), .B2(n_99), .Y(n_150) );
INVx1_ASAP7_75t_L g415 ( .A(n_74), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_74), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_75), .B(n_98), .Y(n_125) );
XOR2xp5_ASAP7_75t_L g521 ( .A(n_76), .B(n_522), .Y(n_521) );
AOI221xp5_ASAP7_75t_SL g78 ( .A1(n_79), .A2(n_384), .B1(n_389), .B2(n_496), .C(n_508), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
OR5x1_ASAP7_75t_L g81 ( .A(n_82), .B(n_275), .C(n_333), .D(n_369), .E(n_376), .Y(n_81) );
NAND3xp33_ASAP7_75t_SL g82 ( .A(n_83), .B(n_221), .C(n_245), .Y(n_82) );
AOI221xp5_ASAP7_75t_L g83 ( .A1(n_84), .A2(n_153), .B1(n_187), .B2(n_192), .C(n_202), .Y(n_83) );
OAI21xp5_ASAP7_75t_SL g355 ( .A1(n_84), .A2(n_356), .B(n_358), .Y(n_355) );
AND2x2_ASAP7_75t_L g84 ( .A(n_85), .B(n_134), .Y(n_84) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_85), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_120), .Y(n_85) );
INVx2_ASAP7_75t_L g191 ( .A(n_86), .Y(n_191) );
AND2x2_ASAP7_75t_L g204 ( .A(n_86), .B(n_136), .Y(n_204) );
AND2x2_ASAP7_75t_L g258 ( .A(n_86), .B(n_135), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_86), .B(n_121), .Y(n_273) );
OA21x2_ASAP7_75t_L g86 ( .A1(n_87), .A2(n_94), .B(n_119), .Y(n_86) );
OA21x2_ASAP7_75t_L g121 ( .A1(n_87), .A2(n_122), .B(n_132), .Y(n_121) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_89), .Y(n_137) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_91), .Y(n_89) );
AND2x2_ASAP7_75t_SL g133 ( .A(n_90), .B(n_91), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g91 ( .A(n_92), .B(n_93), .Y(n_91) );
OAI21xp5_ASAP7_75t_L g94 ( .A1(n_95), .A2(n_108), .B(n_117), .Y(n_94) );
O2A1O1Ixp33_ASAP7_75t_L g95 ( .A1(n_96), .A2(n_97), .B(n_101), .C(n_104), .Y(n_95) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
INVx3_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx2_ASAP7_75t_L g103 ( .A(n_100), .Y(n_103) );
INVx1_ASAP7_75t_L g111 ( .A(n_100), .Y(n_111) );
INVx3_ASAP7_75t_L g169 ( .A(n_102), .Y(n_169) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g160 ( .A(n_103), .Y(n_160) );
BUFx3_ASAP7_75t_L g161 ( .A(n_103), .Y(n_161) );
AND2x6_ASAP7_75t_L g387 ( .A(n_103), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_105), .A2(n_173), .B(n_174), .Y(n_172) );
INVx4_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx3_ASAP7_75t_L g116 ( .A(n_107), .Y(n_116) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_107), .Y(n_130) );
INVx1_ASAP7_75t_L g182 ( .A(n_107), .Y(n_182) );
INVx1_ASAP7_75t_L g388 ( .A(n_107), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_112), .B(n_113), .C(n_114), .Y(n_108) );
O2A1O1Ixp5_ASAP7_75t_L g126 ( .A1(n_109), .A2(n_127), .B(n_128), .C(n_129), .Y(n_126) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_114), .A2(n_143), .B(n_144), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g149 ( .A1(n_114), .A2(n_130), .B1(n_150), .B2(n_151), .Y(n_149) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_114), .A2(n_130), .B1(n_200), .B2(n_201), .Y(n_199) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g123 ( .A1(n_115), .A2(n_124), .B(n_125), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_115), .A2(n_140), .B(n_141), .Y(n_139) );
O2A1O1Ixp5_ASAP7_75t_SL g168 ( .A1(n_115), .A2(n_169), .B(n_170), .C(n_171), .Y(n_168) );
INVx5_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OAI22xp5_ASAP7_75t_SL g158 ( .A1(n_116), .A2(n_130), .B1(n_159), .B2(n_162), .Y(n_158) );
BUFx3_ASAP7_75t_L g131 ( .A(n_117), .Y(n_131) );
OAI21xp5_ASAP7_75t_L g138 ( .A1(n_117), .A2(n_139), .B(n_142), .Y(n_138) );
OAI21xp5_ASAP7_75t_L g167 ( .A1(n_117), .A2(n_168), .B(n_172), .Y(n_167) );
OAI21xp5_ASAP7_75t_L g177 ( .A1(n_117), .A2(n_178), .B(n_183), .Y(n_177) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_118), .Y(n_505) );
AND2x2_ASAP7_75t_L g291 ( .A(n_120), .B(n_232), .Y(n_291) );
AND2x2_ASAP7_75t_L g324 ( .A(n_120), .B(n_136), .Y(n_324) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g231 ( .A(n_121), .B(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g244 ( .A(n_121), .B(n_136), .Y(n_244) );
AND2x2_ASAP7_75t_L g251 ( .A(n_121), .B(n_232), .Y(n_251) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_121), .Y(n_260) );
AND2x2_ASAP7_75t_L g267 ( .A(n_121), .B(n_135), .Y(n_267) );
INVx1_ASAP7_75t_L g298 ( .A(n_121), .Y(n_298) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_126), .B(n_131), .Y(n_122) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_127), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_129), .A2(n_184), .B(n_185), .Y(n_183) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NAND3xp33_ASAP7_75t_L g148 ( .A(n_131), .B(n_149), .C(n_152), .Y(n_148) );
AND2x2_ASAP7_75t_L g386 ( .A(n_131), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g163 ( .A(n_133), .Y(n_163) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_133), .A2(n_167), .B(n_175), .Y(n_166) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_133), .A2(n_177), .B(n_186), .Y(n_176) );
INVx1_ASAP7_75t_L g274 ( .A(n_134), .Y(n_274) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_146), .Y(n_134) );
INVx2_ASAP7_75t_L g230 ( .A(n_135), .Y(n_230) );
AND2x2_ASAP7_75t_L g252 ( .A(n_135), .B(n_191), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_135), .B(n_298), .Y(n_303) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_136), .B(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g375 ( .A(n_136), .B(n_339), .Y(n_375) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B(n_145), .Y(n_136) );
INVx4_ASAP7_75t_L g152 ( .A(n_137), .Y(n_152) );
INVx2_ASAP7_75t_L g189 ( .A(n_146), .Y(n_189) );
INVx3_ASAP7_75t_L g290 ( .A(n_146), .Y(n_290) );
OR2x2_ASAP7_75t_L g320 ( .A(n_146), .B(n_321), .Y(n_320) );
NOR2x1_ASAP7_75t_L g346 ( .A(n_146), .B(n_230), .Y(n_346) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
INVx1_ASAP7_75t_L g233 ( .A(n_147), .Y(n_233) );
AO21x1_ASAP7_75t_L g232 ( .A1(n_149), .A2(n_152), .B(n_233), .Y(n_232) );
AOI33xp33_ASAP7_75t_L g366 ( .A1(n_153), .A2(n_204), .A3(n_218), .B1(n_290), .B2(n_367), .B3(n_368), .Y(n_366) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
OR2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_164), .Y(n_154) );
OR2x2_ASAP7_75t_L g219 ( .A(n_155), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_155), .B(n_216), .Y(n_278) );
OR2x2_ASAP7_75t_L g331 ( .A(n_155), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g257 ( .A(n_156), .B(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g282 ( .A(n_156), .B(n_164), .Y(n_282) );
AND2x2_ASAP7_75t_L g349 ( .A(n_156), .B(n_194), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_156), .A2(n_249), .B(n_375), .Y(n_374) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g196 ( .A(n_157), .Y(n_196) );
INVx1_ASAP7_75t_L g209 ( .A(n_157), .Y(n_209) );
AND2x2_ASAP7_75t_L g228 ( .A(n_157), .B(n_198), .Y(n_228) );
AND2x2_ASAP7_75t_L g277 ( .A(n_157), .B(n_197), .Y(n_277) );
INVx2_ASAP7_75t_SL g319 ( .A(n_164), .Y(n_319) );
OR2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_176), .Y(n_164) );
INVx2_ASAP7_75t_L g239 ( .A(n_165), .Y(n_239) );
INVx1_ASAP7_75t_L g370 ( .A(n_165), .Y(n_370) );
AND2x2_ASAP7_75t_L g383 ( .A(n_165), .B(n_264), .Y(n_383) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g210 ( .A(n_166), .Y(n_210) );
OR2x2_ASAP7_75t_L g216 ( .A(n_166), .B(n_217), .Y(n_216) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_166), .Y(n_227) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_176), .Y(n_194) );
AND2x2_ASAP7_75t_L g211 ( .A(n_176), .B(n_197), .Y(n_211) );
INVx1_ASAP7_75t_L g217 ( .A(n_176), .Y(n_217) );
INVx1_ASAP7_75t_L g224 ( .A(n_176), .Y(n_224) );
AND2x2_ASAP7_75t_L g249 ( .A(n_176), .B(n_198), .Y(n_249) );
INVx2_ASAP7_75t_L g265 ( .A(n_176), .Y(n_265) );
AND2x2_ASAP7_75t_L g358 ( .A(n_176), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_176), .B(n_239), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_181), .Y(n_178) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_SL g187 ( .A(n_188), .Y(n_187) );
OR2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
INVx2_ASAP7_75t_L g213 ( .A(n_189), .Y(n_213) );
INVx1_ASAP7_75t_L g242 ( .A(n_189), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_189), .B(n_273), .Y(n_339) );
INVx1_ASAP7_75t_SL g299 ( .A(n_190), .Y(n_299) );
INVx2_ASAP7_75t_L g220 ( .A(n_191), .Y(n_220) );
AND2x2_ASAP7_75t_L g289 ( .A(n_191), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g305 ( .A(n_191), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_195), .Y(n_192) );
INVx1_ASAP7_75t_L g367 ( .A(n_193), .Y(n_367) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g222 ( .A(n_195), .B(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g325 ( .A(n_195), .B(n_315), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_195), .A2(n_336), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
AND2x2_ASAP7_75t_L g238 ( .A(n_196), .B(n_239), .Y(n_238) );
BUFx2_ASAP7_75t_L g263 ( .A(n_196), .Y(n_263) );
INVx1_ASAP7_75t_L g287 ( .A(n_196), .Y(n_287) );
OR2x2_ASAP7_75t_L g351 ( .A(n_197), .B(n_210), .Y(n_351) );
NOR2xp67_ASAP7_75t_L g359 ( .A(n_197), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g264 ( .A(n_198), .B(n_265), .Y(n_264) );
BUFx2_ASAP7_75t_L g271 ( .A(n_198), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_205), .B1(n_212), .B2(n_214), .Y(n_202) );
OR2x2_ASAP7_75t_L g281 ( .A(n_203), .B(n_231), .Y(n_281) );
INVx1_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
AOI222xp33_ASAP7_75t_L g322 ( .A1(n_204), .A2(n_323), .B1(n_325), .B2(n_326), .C1(n_327), .C2(n_330), .Y(n_322) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_211), .Y(n_206) );
INVx1_ASAP7_75t_SL g207 ( .A(n_208), .Y(n_207) );
OR2x2_ASAP7_75t_L g269 ( .A(n_208), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
AND2x2_ASAP7_75t_SL g223 ( .A(n_210), .B(n_224), .Y(n_223) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_210), .Y(n_294) );
AND2x2_ASAP7_75t_L g342 ( .A(n_210), .B(n_211), .Y(n_342) );
INVx1_ASAP7_75t_L g360 ( .A(n_210), .Y(n_360) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g326 ( .A(n_213), .B(n_252), .Y(n_326) );
AND2x2_ASAP7_75t_L g368 ( .A(n_213), .B(n_244), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_218), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_215), .B(n_263), .Y(n_350) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_216), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g243 ( .A(n_220), .B(n_244), .Y(n_243) );
INVx3_ASAP7_75t_L g311 ( .A(n_220), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_225), .B(n_229), .C(n_234), .Y(n_221) );
INVxp67_ASAP7_75t_L g235 ( .A(n_222), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_223), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_223), .B(n_270), .Y(n_365) );
BUFx3_ASAP7_75t_L g329 ( .A(n_224), .Y(n_329) );
INVx1_ASAP7_75t_L g236 ( .A(n_225), .Y(n_236) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_228), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g255 ( .A(n_227), .B(n_249), .Y(n_255) );
INVx1_ASAP7_75t_SL g295 ( .A(n_228), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
INVx1_ASAP7_75t_L g285 ( .A(n_230), .Y(n_285) );
AND2x2_ASAP7_75t_L g308 ( .A(n_230), .B(n_291), .Y(n_308) );
INVx1_ASAP7_75t_SL g279 ( .A(n_231), .Y(n_279) );
INVx1_ASAP7_75t_L g306 ( .A(n_232), .Y(n_306) );
AOI31xp33_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .A3(n_237), .B(n_240), .Y(n_234) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g327 ( .A(n_238), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g301 ( .A(n_239), .Y(n_301) );
BUFx2_ASAP7_75t_L g315 ( .A(n_239), .Y(n_315) );
AND2x2_ASAP7_75t_L g343 ( .A(n_239), .B(n_264), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_243), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx1_ASAP7_75t_SL g316 ( .A(n_243), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_244), .B(n_311), .Y(n_357) );
AND2x2_ASAP7_75t_L g364 ( .A(n_244), .B(n_290), .Y(n_364) );
AOI211xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_250), .B(n_253), .C(n_268), .Y(n_245) );
INVxp67_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AOI221xp5_ASAP7_75t_L g276 ( .A1(n_250), .A2(n_277), .B1(n_278), .B2(n_279), .C(n_280), .Y(n_276) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AND2x2_ASAP7_75t_L g284 ( .A(n_251), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g321 ( .A(n_252), .Y(n_321) );
OAI32xp33_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_256), .A3(n_259), .B1(n_261), .B2(n_266), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_255), .A2(n_308), .B(n_309), .C(n_312), .Y(n_307) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
OAI21xp5_ASAP7_75t_SL g371 ( .A1(n_263), .A2(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_L g332 ( .A(n_264), .Y(n_332) );
INVxp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_270), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g318 ( .A(n_270), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g335 ( .A(n_272), .Y(n_335) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
NAND4xp25_ASAP7_75t_SL g275 ( .A(n_276), .B(n_288), .C(n_307), .D(n_322), .Y(n_275) );
AND2x2_ASAP7_75t_L g314 ( .A(n_277), .B(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g336 ( .A(n_277), .B(n_329), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_279), .B(n_311), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B1(n_283), .B2(n_286), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_281), .A2(n_332), .B1(n_363), .B2(n_365), .Y(n_362) );
O2A1O1Ixp33_ASAP7_75t_L g369 ( .A1(n_281), .A2(n_370), .B(n_371), .C(n_374), .Y(n_369) );
INVx2_ASAP7_75t_L g340 ( .A(n_282), .Y(n_340) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AOI222xp33_ASAP7_75t_L g334 ( .A1(n_284), .A2(n_318), .B1(n_335), .B2(n_336), .C1(n_337), .C2(n_340), .Y(n_334) );
O2A1O1Ixp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_291), .B(n_292), .C(n_296), .Y(n_288) );
INVx1_ASAP7_75t_L g354 ( .A(n_289), .Y(n_354) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OAI22xp33_ASAP7_75t_L g296 ( .A1(n_293), .A2(n_297), .B1(n_300), .B2(n_302), .Y(n_296) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g323 ( .A(n_305), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g381 ( .A(n_308), .Y(n_381) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OAI22xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_316), .B1(n_317), .B2(n_320), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_315), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g372 ( .A(n_320), .Y(n_372) );
INVx1_ASAP7_75t_L g353 ( .A(n_324), .Y(n_353) );
CKINVDCx16_ASAP7_75t_R g380 ( .A(n_326), .Y(n_380) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND5xp2_ASAP7_75t_L g333 ( .A(n_334), .B(n_341), .C(n_355), .D(n_361), .E(n_366), .Y(n_333) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B(n_344), .C(n_347), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI31xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_350), .A3(n_351), .B(n_352), .Y(n_347) );
INVx1_ASAP7_75t_L g373 ( .A(n_349), .Y(n_373) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI222xp33_ASAP7_75t_L g376 ( .A1(n_363), .A2(n_365), .B1(n_377), .B2(n_380), .C1(n_381), .C2(n_382), .Y(n_376) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_385), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_386), .Y(n_385) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_387), .A2(n_504), .B(n_519), .Y(n_518) );
XOR2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_406), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_392), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B1(n_398), .B2(n_404), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_398), .Y(n_404) );
INVx1_ASAP7_75t_L g403 ( .A(n_399), .Y(n_403) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g522 ( .A(n_408), .Y(n_522) );
NAND2x1_ASAP7_75t_L g408 ( .A(n_409), .B(n_463), .Y(n_408) );
NOR3xp33_ASAP7_75t_SL g409 ( .A(n_410), .B(n_433), .C(n_450), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B1(n_423), .B2(n_424), .Y(n_410) );
NAND2x1p5_ASAP7_75t_L g412 ( .A(n_413), .B(n_420), .Y(n_412) );
AND2x4_ASAP7_75t_L g442 ( .A(n_413), .B(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_L g448 ( .A(n_413), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_418), .Y(n_413) );
INVx2_ASAP7_75t_L g438 ( .A(n_414), .Y(n_438) );
AND2x2_ASAP7_75t_L g469 ( .A(n_414), .B(n_431), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_414), .B(n_432), .Y(n_473) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_417), .Y(n_419) );
AND2x2_ASAP7_75t_L g428 ( .A(n_418), .B(n_422), .Y(n_428) );
INVx2_ASAP7_75t_L g455 ( .A(n_418), .Y(n_455) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g443 ( .A(n_421), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g480 ( .A(n_421), .B(n_455), .Y(n_480) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g454 ( .A(n_422), .B(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g462 ( .A(n_422), .B(n_455), .Y(n_462) );
INVx1_ASAP7_75t_L g472 ( .A(n_422), .Y(n_472) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
CKINVDCx16_ASAP7_75t_R g425 ( .A(n_426), .Y(n_425) );
OR2x6_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x6_ASAP7_75t_L g436 ( .A(n_428), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g439 ( .A(n_432), .Y(n_439) );
INVx1_ASAP7_75t_L g444 ( .A(n_432), .Y(n_444) );
AND2x2_ASAP7_75t_L g457 ( .A(n_432), .B(n_438), .Y(n_457) );
OAI21xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B(n_440), .Y(n_433) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g477 ( .A(n_437), .B(n_462), .Y(n_477) );
AND2x6_ASAP7_75t_L g484 ( .A(n_437), .B(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g491 ( .A(n_437), .B(n_480), .Y(n_491) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g449 ( .A(n_444), .Y(n_449) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B1(n_458), .B2(n_459), .Y(n_450) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_456), .Y(n_453) );
INVx2_ASAP7_75t_L g485 ( .A(n_454), .Y(n_485) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2x1p5_ASAP7_75t_L g461 ( .A(n_457), .B(n_462), .Y(n_461) );
AND2x4_ASAP7_75t_L g494 ( .A(n_457), .B(n_480), .Y(n_494) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g468 ( .A(n_462), .B(n_469), .Y(n_468) );
AND4x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_474), .C(n_481), .D(n_489), .Y(n_463) );
BUFx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx5_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx8_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g479 ( .A(n_469), .B(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OR2x6_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVx1_ASAP7_75t_L g488 ( .A(n_473), .Y(n_488) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx6_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x4_ASAP7_75t_L g487 ( .A(n_480), .B(n_488), .Y(n_487) );
INVx4_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx11_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx2_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_498), .Y(n_497) );
AND3x1_ASAP7_75t_SL g498 ( .A(n_499), .B(n_504), .C(n_506), .Y(n_498) );
INVxp67_ASAP7_75t_L g514 ( .A(n_499), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
INVx1_ASAP7_75t_SL g516 ( .A(n_504), .Y(n_516) );
INVx1_ASAP7_75t_L g526 ( .A(n_504), .Y(n_526) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_505), .B(n_507), .Y(n_519) );
OR2x2_ASAP7_75t_SL g525 ( .A(n_506), .B(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
OAI322xp33_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_511), .A3(n_515), .B1(n_517), .B2(n_520), .C1(n_521), .C2(n_523), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
endmodule