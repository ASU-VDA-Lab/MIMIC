module fake_ariane_749_n_1746 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1746);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1746;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1733;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_159),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_107),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_17),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_16),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_58),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_53),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_38),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

BUFx8_ASAP7_75t_SL g171 ( 
.A(n_14),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_69),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_67),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_33),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_24),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_51),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_52),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_82),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_140),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_79),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_5),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_100),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_132),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_30),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_47),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_75),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_24),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_126),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_46),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_0),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_38),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_15),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_102),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_15),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_96),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_40),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_138),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_74),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_110),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_12),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_122),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_125),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_39),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_142),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_129),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_66),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_137),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_89),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_54),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_134),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_33),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_114),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_98),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_141),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_20),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_97),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_157),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_99),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_65),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_21),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_22),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_133),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_14),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_62),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_71),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_119),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_93),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_55),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_50),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_46),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_148),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_34),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_83),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_103),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_21),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_49),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_146),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_4),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_144),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_155),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_111),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_43),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_0),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_61),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_117),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_37),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_10),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_57),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_39),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_149),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_70),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_59),
.Y(n_260)
);

BUFx8_ASAP7_75t_SL g261 ( 
.A(n_90),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_84),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_22),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_25),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_3),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_11),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_101),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_26),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_76),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_153),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_19),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_108),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_12),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_17),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_68),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_34),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_32),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_13),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_20),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_56),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_44),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_81),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_124),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_91),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_19),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_23),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_31),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_127),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_72),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_60),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_25),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_85),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_18),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_104),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_41),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_95),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_27),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_105),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_135),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_31),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_7),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_121),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_113),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_41),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_40),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_35),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_27),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_42),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_88),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_26),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_147),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_2),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_29),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_6),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_1),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_130),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_9),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_274),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_274),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_171),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_261),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_179),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_274),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_191),
.B(n_1),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_274),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_233),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_234),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_274),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_265),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_190),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_235),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_265),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_236),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_221),
.B(n_2),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_251),
.B(n_3),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_247),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_273),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_273),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_286),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_286),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_284),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_172),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_183),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_172),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_176),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_288),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_176),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_183),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_188),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_188),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_239),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_163),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_239),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_164),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_187),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_201),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_203),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_219),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_238),
.B(n_4),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_256),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_305),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_208),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_241),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_163),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_228),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_312),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_241),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_199),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_315),
.Y(n_369)
);

NAND2xp33_ASAP7_75t_R g370 ( 
.A(n_160),
.B(n_92),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_232),
.Y(n_371)
);

BUFx2_ASAP7_75t_SL g372 ( 
.A(n_232),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_229),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_244),
.Y(n_374)
);

INVxp33_ASAP7_75t_SL g375 ( 
.A(n_168),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_244),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_238),
.B(n_5),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_232),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_199),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_260),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_174),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_243),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_250),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_260),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_197),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_178),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_279),
.B(n_6),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_198),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_254),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_246),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_255),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_277),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_279),
.B(n_7),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_319),
.Y(n_394)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_318),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_322),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_319),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_355),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_323),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_323),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_358),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_325),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_332),
.B(n_282),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_343),
.B(n_162),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_326),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_R g407 ( 
.A(n_321),
.B(n_205),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_325),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_328),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_328),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_342),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_343),
.B(n_165),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_336),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_342),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_331),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_348),
.B(n_258),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_361),
.A2(n_196),
.B1(n_195),
.B2(n_313),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_344),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_344),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_345),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_R g421 ( 
.A(n_356),
.B(n_206),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_341),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_348),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_345),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_327),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_346),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_347),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_366),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_347),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_357),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_349),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_349),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_368),
.B(n_216),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_350),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_324),
.B(n_216),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_350),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_368),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_320),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_362),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_351),
.B(n_218),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_353),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_363),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_365),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_363),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_367),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_367),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_340),
.B(n_282),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_364),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_374),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_373),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_374),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_376),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_364),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_376),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_380),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_382),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_380),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_384),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_385),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_384),
.B(n_169),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_329),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_329),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_381),
.B(n_218),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_415),
.B(n_371),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_401),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_423),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_460),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_464),
.A2(n_359),
.B1(n_387),
.B2(n_334),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_423),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_460),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_437),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_411),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_423),
.B(n_377),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_435),
.B(n_372),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_398),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_415),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_437),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_437),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_421),
.B(n_333),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_445),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_398),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_464),
.A2(n_352),
.B1(n_375),
.B2(n_335),
.Y(n_483)
);

NAND2xp33_ASAP7_75t_L g484 ( 
.A(n_421),
.B(n_383),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_441),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_464),
.B(n_360),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_449),
.Y(n_487)
);

AO22x1_ASAP7_75t_L g488 ( 
.A1(n_464),
.A2(n_291),
.B1(n_168),
.B2(n_193),
.Y(n_488)
);

BUFx6f_ASAP7_75t_SL g489 ( 
.A(n_464),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_445),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_404),
.B(n_372),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_445),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_404),
.B(n_389),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_401),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_430),
.B(n_391),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_450),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_449),
.B(n_330),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_402),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_SL g499 ( 
.A(n_430),
.B(n_370),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_420),
.A2(n_393),
.B1(n_354),
.B2(n_306),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_402),
.Y(n_501)
);

NAND3xp33_ASAP7_75t_L g502 ( 
.A(n_416),
.B(n_195),
.C(n_193),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_449),
.B(n_386),
.Y(n_503)
);

INVx5_ASAP7_75t_L g504 ( 
.A(n_411),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_408),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_420),
.A2(n_310),
.B1(n_300),
.B2(n_301),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_432),
.A2(n_285),
.B1(n_308),
.B2(n_314),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_454),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_450),
.Y(n_509)
);

INVx4_ASAP7_75t_SL g510 ( 
.A(n_411),
.Y(n_510)
);

INVx4_ASAP7_75t_SL g511 ( 
.A(n_411),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_432),
.A2(n_392),
.B1(n_390),
.B2(n_388),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_408),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_450),
.Y(n_514)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_441),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_439),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_440),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_434),
.A2(n_392),
.B1(n_390),
.B2(n_388),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_434),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_444),
.B(n_175),
.Y(n_520)
);

INVx4_ASAP7_75t_SL g521 ( 
.A(n_411),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_443),
.Y(n_522)
);

INVx4_ASAP7_75t_SL g523 ( 
.A(n_411),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_411),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_408),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_396),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_404),
.B(n_379),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_443),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_410),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_454),
.B(n_378),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_454),
.B(n_386),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_451),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_448),
.B(n_337),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_448),
.B(n_166),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_452),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_414),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_452),
.Y(n_537)
);

NAND3xp33_ASAP7_75t_L g538 ( 
.A(n_416),
.B(n_293),
.C(n_295),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_414),
.Y(n_539)
);

AND2x2_ASAP7_75t_SL g540 ( 
.A(n_441),
.B(n_177),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_414),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_441),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_459),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_435),
.A2(n_211),
.B1(n_231),
.B2(n_223),
.Y(n_544)
);

OR2x6_ASAP7_75t_L g545 ( 
.A(n_417),
.B(n_337),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_410),
.Y(n_546)
);

BUFx8_ASAP7_75t_SL g547 ( 
.A(n_428),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_457),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_448),
.B(n_338),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_406),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_459),
.A2(n_339),
.B1(n_338),
.B2(n_263),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_L g552 ( 
.A(n_407),
.B(n_289),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_463),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_463),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_433),
.B(n_405),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_419),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_419),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_441),
.B(n_181),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_414),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_433),
.B(n_209),
.Y(n_560)
);

AND2x6_ASAP7_75t_L g561 ( 
.A(n_419),
.B(n_289),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_428),
.Y(n_562)
);

OAI22xp33_ASAP7_75t_L g563 ( 
.A1(n_413),
.A2(n_196),
.B1(n_278),
.B2(n_281),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_419),
.B(n_339),
.Y(n_564)
);

BUFx6f_ASAP7_75t_SL g565 ( 
.A(n_422),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_414),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_414),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_419),
.B(n_210),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_410),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_414),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_405),
.B(n_182),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_436),
.B(n_220),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_436),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_425),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_417),
.B(n_240),
.Y(n_575)
);

BUFx6f_ASAP7_75t_SL g576 ( 
.A(n_418),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_407),
.B(n_240),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_418),
.Y(n_578)
);

INVx5_ASAP7_75t_L g579 ( 
.A(n_418),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_436),
.B(n_412),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_418),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_436),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_412),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_418),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_426),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_436),
.B(n_222),
.Y(n_586)
);

INVx6_ASAP7_75t_L g587 ( 
.A(n_418),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_418),
.B(n_184),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_427),
.Y(n_589)
);

INVx6_ASAP7_75t_L g590 ( 
.A(n_427),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_462),
.B(n_240),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_427),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_394),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_394),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_397),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_427),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_427),
.Y(n_597)
);

NAND2x1p5_ASAP7_75t_L g598 ( 
.A(n_427),
.B(n_200),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_397),
.Y(n_599)
);

AND2x6_ASAP7_75t_L g600 ( 
.A(n_427),
.B(n_289),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_424),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_462),
.B(n_263),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_461),
.B(n_202),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_424),
.B(n_160),
.Y(n_604)
);

AND2x6_ASAP7_75t_L g605 ( 
.A(n_424),
.B(n_289),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_395),
.Y(n_606)
);

AND3x2_ASAP7_75t_L g607 ( 
.A(n_429),
.B(n_275),
.C(n_214),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_461),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_399),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_429),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_429),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_L g612 ( 
.A1(n_575),
.A2(n_291),
.B1(n_268),
.B2(n_271),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_611),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_608),
.B(n_431),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_499),
.B(n_161),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_493),
.B(n_431),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_611),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_593),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_555),
.B(n_431),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_601),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_601),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_555),
.B(n_438),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_540),
.A2(n_170),
.B1(n_167),
.B2(n_161),
.Y(n_623)
);

OAI221xp5_ASAP7_75t_L g624 ( 
.A1(n_469),
.A2(n_304),
.B1(n_268),
.B2(n_271),
.C(n_276),
.Y(n_624)
);

NAND3xp33_ASAP7_75t_L g625 ( 
.A(n_469),
.B(n_276),
.C(n_278),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_540),
.B(n_499),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_601),
.Y(n_627)
);

A2O1A1Ixp33_ASAP7_75t_L g628 ( 
.A1(n_571),
.A2(n_403),
.B(n_409),
.C(n_456),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_583),
.B(n_438),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_591),
.B(n_438),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_533),
.A2(n_447),
.B1(n_458),
.B2(n_456),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_471),
.B(n_369),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_594),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_602),
.B(n_442),
.Y(n_634)
);

AOI22x1_ASAP7_75t_L g635 ( 
.A1(n_556),
.A2(n_453),
.B1(n_458),
.B2(n_456),
.Y(n_635)
);

A2O1A1Ixp33_ASAP7_75t_L g636 ( 
.A1(n_571),
.A2(n_403),
.B(n_409),
.C(n_455),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_485),
.B(n_167),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_533),
.A2(n_458),
.B1(n_455),
.B2(n_453),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_491),
.B(n_442),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_485),
.B(n_515),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_610),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_610),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_580),
.B(n_442),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_468),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_531),
.B(n_263),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_485),
.B(n_170),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_534),
.B(n_446),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_515),
.A2(n_287),
.B1(n_281),
.B2(n_304),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_486),
.B(n_446),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_560),
.B(n_446),
.Y(n_650)
);

NAND2x1p5_ASAP7_75t_L g651 ( 
.A(n_515),
.B(n_447),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_533),
.B(n_447),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_549),
.B(n_453),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_595),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_577),
.B(n_173),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_573),
.A2(n_455),
.B(n_462),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_574),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_610),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_549),
.B(n_400),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_466),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_548),
.B(n_287),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_532),
.B(n_173),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_486),
.B(n_257),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_549),
.B(n_400),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_489),
.A2(n_294),
.B1(n_180),
.B2(n_185),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_489),
.A2(n_294),
.B1(n_180),
.B2(n_185),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_475),
.A2(n_269),
.B1(n_270),
.B2(n_272),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_542),
.B(n_400),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_475),
.B(n_520),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_509),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_599),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_503),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_520),
.B(n_264),
.Y(n_673)
);

INVx8_ASAP7_75t_L g674 ( 
.A(n_565),
.Y(n_674)
);

OAI22xp33_ASAP7_75t_L g675 ( 
.A1(n_545),
.A2(n_293),
.B1(n_313),
.B2(n_295),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_542),
.B(n_400),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_542),
.B(n_186),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_609),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_524),
.B(n_186),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_494),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_477),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_524),
.B(n_189),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_SL g683 ( 
.A1(n_465),
.A2(n_297),
.B1(n_307),
.B2(n_317),
.Y(n_683)
);

AND2x4_ASAP7_75t_SL g684 ( 
.A(n_574),
.B(n_400),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_524),
.B(n_189),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_506),
.A2(n_297),
.B1(n_307),
.B2(n_311),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_492),
.B(n_192),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_519),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_492),
.B(n_192),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_506),
.A2(n_204),
.B1(n_316),
.B2(n_296),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_494),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_527),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_522),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_524),
.B(n_194),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_564),
.B(n_194),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_507),
.A2(n_280),
.B1(n_237),
.B2(n_226),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_564),
.B(n_269),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_483),
.B(n_266),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_502),
.B(n_270),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_497),
.B(n_272),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_548),
.B(n_298),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_550),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_474),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_487),
.A2(n_298),
.B1(n_303),
.B2(n_302),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_564),
.B(n_299),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_541),
.B(n_567),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_488),
.B(n_299),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_476),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_538),
.B(n_302),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_508),
.B(n_303),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_528),
.B(n_309),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_557),
.B(n_309),
.Y(n_712)
);

INVxp33_ASAP7_75t_L g713 ( 
.A(n_547),
.Y(n_713)
);

AND2x6_ASAP7_75t_SL g714 ( 
.A(n_545),
.B(n_290),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_535),
.B(n_267),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_482),
.B(n_8),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_537),
.B(n_212),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_505),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_543),
.B(n_207),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_484),
.A2(n_213),
.B1(n_292),
.B2(n_225),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_474),
.B(n_248),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_553),
.B(n_215),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_474),
.B(n_249),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_484),
.A2(n_245),
.B1(n_283),
.B2(n_217),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_554),
.B(n_558),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_558),
.B(n_224),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_582),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_481),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_541),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_490),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_517),
.B(n_253),
.Y(n_731)
);

O2A1O1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_604),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_557),
.B(n_11),
.Y(n_733)
);

O2A1O1Ixp5_ASAP7_75t_L g734 ( 
.A1(n_584),
.A2(n_227),
.B(n_230),
.C(n_242),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_541),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_513),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_496),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_568),
.B(n_252),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_525),
.Y(n_739)
);

NOR3xp33_ASAP7_75t_L g740 ( 
.A(n_495),
.B(n_259),
.C(n_262),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_541),
.B(n_289),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_514),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_572),
.B(n_13),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_467),
.B(n_470),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_586),
.B(n_16),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_472),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_509),
.B(n_18),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_467),
.B(n_23),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_478),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_525),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_529),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_529),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_516),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_546),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_546),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_495),
.B(n_395),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_498),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_567),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_507),
.A2(n_395),
.B1(n_29),
.B2(n_30),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_603),
.B(n_28),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_567),
.B(n_395),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_569),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_470),
.B(n_395),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_603),
.B(n_28),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_569),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_479),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_552),
.A2(n_395),
.B1(n_35),
.B2(n_36),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_479),
.B(n_32),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_479),
.B(n_36),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_530),
.B(n_526),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_480),
.B(n_37),
.Y(n_771)
);

AOI221xp5_ASAP7_75t_SL g772 ( 
.A1(n_512),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.C(n_45),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_480),
.B(n_45),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_584),
.B(n_536),
.Y(n_774)
);

NOR3xp33_ASAP7_75t_L g775 ( 
.A(n_563),
.B(n_526),
.C(n_516),
.Y(n_775)
);

INVx8_ASAP7_75t_L g776 ( 
.A(n_565),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_729),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_619),
.A2(n_584),
.B(n_473),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_622),
.A2(n_536),
.B(n_559),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_774),
.A2(n_536),
.B(n_559),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_672),
.B(n_562),
.Y(n_781)
);

BUFx5_ASAP7_75t_L g782 ( 
.A(n_752),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_729),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_774),
.A2(n_559),
.B(n_566),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_660),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_669),
.A2(n_552),
.B1(n_585),
.B2(n_545),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_692),
.B(n_544),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_706),
.A2(n_473),
.B(n_570),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_669),
.A2(n_576),
.B1(n_500),
.B2(n_590),
.Y(n_789)
);

NAND2xp33_ASAP7_75t_SL g790 ( 
.A(n_731),
.B(n_518),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_626),
.B(n_539),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_618),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_706),
.A2(n_473),
.B(n_570),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_614),
.B(n_500),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_643),
.A2(n_570),
.B(n_566),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_616),
.B(n_551),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_640),
.A2(n_539),
.B(n_566),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_626),
.B(n_539),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_644),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_632),
.B(n_501),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_625),
.A2(n_587),
.B1(n_590),
.B2(n_592),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_640),
.A2(n_596),
.B(n_589),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_629),
.A2(n_676),
.B(n_668),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_651),
.A2(n_623),
.B1(n_654),
.B2(n_633),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_628),
.A2(n_597),
.B(n_596),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_650),
.A2(n_597),
.B(n_589),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_700),
.B(n_512),
.Y(n_807)
);

OR2x6_ASAP7_75t_SL g808 ( 
.A(n_704),
.B(n_547),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_645),
.B(n_518),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_647),
.B(n_630),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_634),
.B(n_578),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_673),
.B(n_592),
.Y(n_812)
);

AOI21x1_ASAP7_75t_L g813 ( 
.A1(n_656),
.A2(n_578),
.B(n_581),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_673),
.B(n_590),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_698),
.A2(n_576),
.B1(n_587),
.B2(n_588),
.Y(n_815)
);

AOI21x1_ASAP7_75t_L g816 ( 
.A1(n_761),
.A2(n_581),
.B(n_588),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_744),
.B(n_567),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_671),
.Y(n_818)
);

O2A1O1Ixp5_ASAP7_75t_L g819 ( 
.A1(n_743),
.A2(n_606),
.B(n_598),
.C(n_587),
.Y(n_819)
);

NOR2x1_ASAP7_75t_R g820 ( 
.A(n_753),
.B(n_501),
.Y(n_820)
);

BUFx8_ASAP7_75t_SL g821 ( 
.A(n_657),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_698),
.A2(n_504),
.B(n_579),
.C(n_598),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_636),
.A2(n_579),
.B(n_504),
.Y(n_823)
);

O2A1O1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_624),
.A2(n_607),
.B(n_523),
.C(n_521),
.Y(n_824)
);

O2A1O1Ixp5_ASAP7_75t_L g825 ( 
.A1(n_745),
.A2(n_606),
.B(n_523),
.C(n_521),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_639),
.A2(n_579),
.B(n_504),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_744),
.B(n_504),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_729),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_738),
.A2(n_579),
.B(n_606),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_703),
.B(n_523),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_678),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_702),
.B(n_521),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_SL g833 ( 
.A(n_674),
.B(n_561),
.Y(n_833)
);

INVx11_ASAP7_75t_L g834 ( 
.A(n_674),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_688),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_649),
.B(n_511),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_649),
.B(n_639),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_620),
.A2(n_511),
.B(n_510),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_680),
.Y(n_839)
);

O2A1O1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_612),
.A2(n_511),
.B(n_510),
.C(n_561),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_651),
.A2(n_395),
.B1(n_510),
.B2(n_561),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_612),
.B(n_561),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_693),
.B(n_561),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_621),
.A2(n_641),
.B(n_627),
.Y(n_844)
);

NOR3xp33_ASAP7_75t_L g845 ( 
.A(n_675),
.B(n_605),
.C(n_600),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_691),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_652),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_771),
.B(n_395),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_653),
.A2(n_725),
.B1(n_759),
.B2(n_712),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_690),
.A2(n_605),
.B1(n_600),
.B2(n_64),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_642),
.A2(n_600),
.B(n_605),
.Y(n_851)
);

INVx1_ASAP7_75t_SL g852 ( 
.A(n_757),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_712),
.B(n_631),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_659),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_631),
.B(n_600),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_664),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_638),
.B(n_600),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_638),
.B(n_605),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_658),
.A2(n_605),
.B(n_63),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_675),
.A2(n_48),
.B(n_73),
.C(n_77),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_728),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_770),
.B(n_78),
.Y(n_862)
);

OAI21xp33_ASAP7_75t_L g863 ( 
.A1(n_667),
.A2(n_80),
.B(n_86),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_663),
.B(n_87),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_663),
.B(n_106),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_637),
.A2(n_677),
.B(n_646),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_730),
.A2(n_112),
.B(n_115),
.C(n_118),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_637),
.A2(n_677),
.B(n_646),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_674),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_687),
.A2(n_123),
.B(n_131),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_727),
.A2(n_143),
.B(n_150),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_689),
.A2(n_151),
.B(n_766),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_715),
.A2(n_717),
.B(n_719),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_734),
.A2(n_635),
.B(n_737),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_699),
.B(n_709),
.Y(n_875)
);

NOR2x1p5_ASAP7_75t_SL g876 ( 
.A(n_746),
.B(n_749),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_722),
.A2(n_694),
.B(n_685),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_710),
.B(n_661),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_699),
.B(n_709),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_708),
.Y(n_880)
);

AOI221xp5_ASAP7_75t_L g881 ( 
.A1(n_686),
.A2(n_648),
.B1(n_683),
.B2(n_775),
.C(n_696),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_679),
.A2(n_685),
.B(n_682),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_679),
.A2(n_682),
.B(n_694),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_655),
.B(n_615),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_742),
.A2(n_711),
.B(n_754),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_771),
.B(n_773),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_661),
.B(n_684),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_755),
.A2(n_765),
.B(n_750),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_681),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_763),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_670),
.A2(n_695),
.B(n_697),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_718),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_670),
.A2(n_705),
.B(n_762),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_759),
.A2(n_769),
.B1(n_768),
.B2(n_733),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_716),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_613),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_736),
.A2(n_751),
.B(n_739),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_729),
.B(n_758),
.Y(n_898)
);

NOR2xp67_ASAP7_75t_L g899 ( 
.A(n_665),
.B(n_666),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_768),
.A2(n_769),
.B1(n_733),
.B2(n_686),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_735),
.A2(n_758),
.B(n_756),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_617),
.A2(n_760),
.B(n_764),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_763),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_690),
.B(n_696),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_707),
.B(n_773),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_720),
.B(n_724),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_747),
.B(n_748),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_747),
.B(n_748),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_761),
.A2(n_726),
.B(n_741),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_776),
.B(n_713),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_741),
.A2(n_740),
.B(n_767),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_735),
.A2(n_758),
.B1(n_723),
.B2(n_721),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_732),
.A2(n_772),
.B(n_701),
.C(n_662),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_735),
.B(n_758),
.Y(n_914)
);

O2A1O1Ixp5_ASAP7_75t_L g915 ( 
.A1(n_735),
.A2(n_743),
.B(n_745),
.C(n_616),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_714),
.B(n_776),
.Y(n_916)
);

OAI21xp33_ASAP7_75t_L g917 ( 
.A1(n_776),
.A2(n_469),
.B(n_698),
.Y(n_917)
);

AOI22x1_ASAP7_75t_L g918 ( 
.A1(n_656),
.A2(n_727),
.B1(n_573),
.B2(n_582),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_669),
.B(n_608),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_618),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_700),
.B(n_468),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_660),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_763),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_644),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_674),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_700),
.B(n_468),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_692),
.B(n_669),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_703),
.B(n_548),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_619),
.A2(n_622),
.B(n_774),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_619),
.A2(n_622),
.B1(n_469),
.B2(n_669),
.Y(n_930)
);

CKINVDCx14_ASAP7_75t_R g931 ( 
.A(n_657),
.Y(n_931)
);

NAND2x1_ASAP7_75t_L g932 ( 
.A(n_729),
.B(n_587),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_619),
.A2(n_622),
.B(n_628),
.Y(n_933)
);

BUFx4f_ASAP7_75t_L g934 ( 
.A(n_674),
.Y(n_934)
);

BUFx8_ASAP7_75t_SL g935 ( 
.A(n_657),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_660),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_619),
.A2(n_622),
.B(n_774),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_692),
.B(n_669),
.Y(n_938)
);

OAI21x1_ASAP7_75t_L g939 ( 
.A1(n_635),
.A2(n_656),
.B(n_706),
.Y(n_939)
);

AOI21xp33_ASAP7_75t_L g940 ( 
.A1(n_698),
.A2(n_673),
.B(n_669),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_619),
.A2(n_622),
.B(n_774),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_619),
.A2(n_622),
.B(n_774),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_660),
.Y(n_943)
);

AOI21x1_ASAP7_75t_L g944 ( 
.A1(n_706),
.A2(n_656),
.B(n_622),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_669),
.B(n_548),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_618),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_692),
.B(n_669),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_669),
.B(n_608),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_644),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_669),
.A2(n_499),
.B1(n_626),
.B2(n_673),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_618),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_669),
.B(n_548),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_669),
.B(n_608),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_669),
.B(n_608),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_669),
.B(n_548),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_619),
.A2(n_622),
.B(n_774),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_669),
.A2(n_499),
.B1(n_626),
.B2(n_673),
.Y(n_957)
);

NOR2x1p5_ASAP7_75t_SL g958 ( 
.A(n_620),
.B(n_621),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_753),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_669),
.B(n_608),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_940),
.B(n_919),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_948),
.B(n_953),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_777),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_921),
.B(n_926),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_939),
.A2(n_813),
.B(n_944),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_934),
.Y(n_966)
);

AO31x2_ASAP7_75t_L g967 ( 
.A1(n_894),
.A2(n_900),
.A3(n_930),
.B(n_877),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_954),
.B(n_960),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_927),
.B(n_938),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_785),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_834),
.Y(n_971)
);

AOI21x1_ASAP7_75t_SL g972 ( 
.A1(n_907),
.A2(n_908),
.B(n_879),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_929),
.A2(n_941),
.B(n_937),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_942),
.A2(n_956),
.B(n_837),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_786),
.B(n_927),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_959),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_938),
.B(n_947),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_805),
.A2(n_918),
.B(n_816),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_809),
.B(n_878),
.Y(n_979)
);

OA21x2_ASAP7_75t_L g980 ( 
.A1(n_915),
.A2(n_819),
.B(n_933),
.Y(n_980)
);

OAI21xp33_ASAP7_75t_L g981 ( 
.A1(n_875),
.A2(n_886),
.B(n_881),
.Y(n_981)
);

OA22x2_ASAP7_75t_L g982 ( 
.A1(n_917),
.A2(n_957),
.B1(n_950),
.B2(n_895),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_777),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_803),
.A2(n_873),
.B(n_810),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_947),
.B(n_847),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_825),
.A2(n_806),
.B(n_819),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_869),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_864),
.A2(n_865),
.B(n_905),
.C(n_790),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_854),
.B(n_856),
.Y(n_989)
);

OAI21x1_ASAP7_75t_SL g990 ( 
.A1(n_866),
.A2(n_868),
.B(n_891),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_792),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_864),
.A2(n_865),
.B(n_905),
.C(n_906),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_924),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_791),
.A2(n_798),
.B(n_915),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_799),
.B(n_949),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_807),
.B(n_787),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_818),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_826),
.A2(n_778),
.B(n_779),
.Y(n_998)
);

AO31x2_ASAP7_75t_L g999 ( 
.A1(n_882),
.A2(n_883),
.A3(n_822),
.B(n_798),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_853),
.B(n_904),
.Y(n_1000)
);

AO31x2_ASAP7_75t_L g1001 ( 
.A1(n_791),
.A2(n_849),
.A3(n_885),
.B(n_913),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_890),
.B(n_923),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_825),
.A2(n_901),
.B(n_802),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_SL g1004 ( 
.A1(n_902),
.A2(n_911),
.B(n_804),
.Y(n_1004)
);

NAND2x1p5_ASAP7_75t_L g1005 ( 
.A(n_890),
.B(n_923),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_780),
.A2(n_784),
.B(n_829),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_795),
.A2(n_955),
.B(n_952),
.Y(n_1007)
);

OAI22x1_ASAP7_75t_L g1008 ( 
.A1(n_945),
.A2(n_787),
.B1(n_800),
.B2(n_895),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_794),
.B(n_796),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_874),
.A2(n_788),
.B(n_793),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_880),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_781),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_924),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_799),
.B(n_949),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_812),
.B(n_831),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_823),
.A2(n_872),
.B(n_893),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_897),
.A2(n_888),
.B(n_838),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_777),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_925),
.B(n_903),
.Y(n_1019)
);

AND2x6_ASAP7_75t_L g1020 ( 
.A(n_842),
.B(n_777),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_783),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_887),
.B(n_928),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_844),
.A2(n_909),
.B(n_898),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_797),
.A2(n_811),
.B(n_814),
.Y(n_1024)
);

AOI21x1_ASAP7_75t_SL g1025 ( 
.A1(n_862),
.A2(n_914),
.B(n_843),
.Y(n_1025)
);

INVx4_ASAP7_75t_L g1026 ( 
.A(n_934),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_814),
.A2(n_842),
.B(n_812),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_835),
.B(n_920),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_898),
.A2(n_871),
.B(n_836),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_946),
.B(n_951),
.Y(n_1030)
);

AO22x1_ASAP7_75t_L g1031 ( 
.A1(n_916),
.A2(n_852),
.B1(n_910),
.B2(n_889),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_932),
.A2(n_848),
.B(n_870),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_851),
.A2(n_840),
.B(n_912),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_899),
.A2(n_884),
.B(n_863),
.C(n_876),
.Y(n_1034)
);

O2A1O1Ixp5_ASAP7_75t_L g1035 ( 
.A1(n_832),
.A2(n_884),
.B(n_801),
.C(n_827),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_931),
.B(n_820),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_783),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_861),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_896),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_783),
.B(n_828),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_783),
.Y(n_1041)
);

NAND2xp33_ASAP7_75t_SL g1042 ( 
.A(n_828),
.B(n_817),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_839),
.B(n_922),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_828),
.A2(n_857),
.B(n_855),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_821),
.B(n_935),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_846),
.B(n_943),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_789),
.B(n_815),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_828),
.B(n_833),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_859),
.A2(n_841),
.B(n_824),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_892),
.B(n_936),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_808),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_SL g1052 ( 
.A1(n_858),
.A2(n_830),
.B(n_860),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_782),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_867),
.A2(n_830),
.B(n_958),
.Y(n_1054)
);

NOR2x1_ASAP7_75t_SL g1055 ( 
.A(n_782),
.B(n_845),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_850),
.A2(n_782),
.B(n_845),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_782),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_782),
.B(n_850),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_782),
.A2(n_937),
.B(n_929),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_916),
.A2(n_939),
.B(n_813),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_939),
.A2(n_813),
.B(n_944),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_890),
.B(n_923),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_959),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_792),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_894),
.A2(n_900),
.B1(n_908),
.B2(n_907),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_939),
.A2(n_813),
.B(n_944),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_939),
.A2(n_813),
.B(n_944),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_SL g1068 ( 
.A1(n_894),
.A2(n_957),
.B(n_950),
.Y(n_1068)
);

O2A1O1Ixp5_ASAP7_75t_L g1069 ( 
.A1(n_900),
.A2(n_894),
.B(n_908),
.C(n_907),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_939),
.A2(n_813),
.B(n_944),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_777),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_919),
.B(n_948),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_929),
.A2(n_941),
.B(n_937),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_939),
.A2(n_813),
.B(n_944),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_939),
.A2(n_813),
.B(n_944),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_939),
.A2(n_813),
.B(n_944),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_777),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_919),
.B(n_948),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_919),
.B(n_948),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_834),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_894),
.A2(n_900),
.B1(n_908),
.B2(n_907),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_939),
.A2(n_813),
.B(n_944),
.Y(n_1082)
);

AOI221xp5_ASAP7_75t_L g1083 ( 
.A1(n_940),
.A2(n_675),
.B1(n_698),
.B2(n_612),
.C(n_881),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_940),
.A2(n_879),
.B(n_875),
.C(n_864),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_939),
.A2(n_813),
.B(n_944),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_919),
.B(n_948),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_919),
.B(n_948),
.Y(n_1087)
);

AOI21x1_ASAP7_75t_L g1088 ( 
.A1(n_813),
.A2(n_883),
.B(n_882),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_919),
.B(n_948),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_777),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_921),
.B(n_926),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_777),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_940),
.A2(n_879),
.B(n_875),
.C(n_864),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_939),
.A2(n_813),
.B(n_944),
.Y(n_1094)
);

O2A1O1Ixp5_ASAP7_75t_L g1095 ( 
.A1(n_900),
.A2(n_894),
.B(n_908),
.C(n_907),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_940),
.A2(n_879),
.B(n_875),
.C(n_864),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_929),
.A2(n_941),
.B(n_937),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_939),
.A2(n_813),
.B(n_944),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_792),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_929),
.A2(n_941),
.B(n_937),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_SL g1101 ( 
.A(n_894),
.B(n_940),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_929),
.A2(n_941),
.B(n_937),
.Y(n_1102)
);

AOI21x1_ASAP7_75t_L g1103 ( 
.A1(n_813),
.A2(n_883),
.B(n_882),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_880),
.Y(n_1104)
);

INVx5_ASAP7_75t_L g1105 ( 
.A(n_777),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_929),
.A2(n_941),
.B(n_937),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1028),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_992),
.A2(n_988),
.B(n_1083),
.C(n_981),
.Y(n_1108)
);

AND2x6_ASAP7_75t_L g1109 ( 
.A(n_1040),
.B(n_1053),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1065),
.A2(n_1081),
.B(n_1059),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1065),
.A2(n_1081),
.B(n_984),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_969),
.B(n_977),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_964),
.B(n_1091),
.Y(n_1113)
);

AND2x6_ASAP7_75t_L g1114 ( 
.A(n_1040),
.B(n_1057),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_969),
.A2(n_977),
.B1(n_1084),
.B2(n_1093),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1069),
.A2(n_1095),
.B(n_1096),
.Y(n_1116)
);

AOI21xp33_ASAP7_75t_SL g1117 ( 
.A1(n_961),
.A2(n_1045),
.B(n_975),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1101),
.A2(n_982),
.B1(n_979),
.B2(n_996),
.Y(n_1118)
);

BUFx12f_ASAP7_75t_L g1119 ( 
.A(n_971),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_962),
.B(n_968),
.Y(n_1120)
);

INVxp67_ASAP7_75t_SL g1121 ( 
.A(n_1013),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_974),
.A2(n_1097),
.B(n_973),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1028),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1030),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1030),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_970),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_976),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_962),
.B(n_968),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1104),
.B(n_1022),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1072),
.B(n_1078),
.Y(n_1130)
);

HAxp5_ASAP7_75t_L g1131 ( 
.A(n_1101),
.B(n_1014),
.CON(n_1131),
.SN(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_991),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_SL g1133 ( 
.A(n_1027),
.B(n_1068),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_1026),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1102),
.A2(n_1106),
.B(n_1073),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1073),
.A2(n_1100),
.B(n_1027),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1104),
.B(n_1022),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1072),
.B(n_1078),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1079),
.B(n_1086),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_1079),
.B(n_1086),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1087),
.B(n_1089),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1011),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_987),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_1105),
.Y(n_1144)
);

CKINVDCx6p67_ASAP7_75t_R g1145 ( 
.A(n_1051),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_1026),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_1105),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_997),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1087),
.B(n_1089),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_1012),
.B(n_993),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_985),
.B(n_1063),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1038),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1100),
.A2(n_998),
.B(n_1029),
.Y(n_1153)
);

AND2x2_ASAP7_75t_SL g1154 ( 
.A(n_1047),
.B(n_1015),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1006),
.A2(n_1024),
.B(n_1058),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1064),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1015),
.A2(n_985),
.B1(n_1058),
.B2(n_1034),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_SL g1158 ( 
.A1(n_1007),
.A2(n_994),
.B(n_1032),
.C(n_1024),
.Y(n_1158)
);

AOI21xp33_ASAP7_75t_L g1159 ( 
.A1(n_1004),
.A2(n_1008),
.B(n_1009),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1039),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_995),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1019),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_1080),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1002),
.B(n_1062),
.Y(n_1164)
);

BUFx12f_ASAP7_75t_L g1165 ( 
.A(n_966),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_1105),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1099),
.B(n_1002),
.Y(n_1167)
);

AO21x2_ASAP7_75t_L g1168 ( 
.A1(n_990),
.A2(n_994),
.B(n_965),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_983),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_983),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_989),
.B(n_1031),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_989),
.B(n_1005),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1036),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1000),
.B(n_1020),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_1041),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1005),
.B(n_1000),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1020),
.B(n_967),
.Y(n_1177)
);

OAI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_1041),
.A2(n_963),
.B1(n_1021),
.B2(n_1071),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_983),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_SL g1180 ( 
.A1(n_1048),
.A2(n_1055),
.B(n_1044),
.Y(n_1180)
);

INVx5_ASAP7_75t_L g1181 ( 
.A(n_1020),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_963),
.B(n_1021),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_967),
.A2(n_980),
.B1(n_1052),
.B2(n_1071),
.Y(n_1183)
);

INVx4_ASAP7_75t_SL g1184 ( 
.A(n_1020),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_1018),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1016),
.A2(n_980),
.B(n_986),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_1018),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1077),
.B(n_1037),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1043),
.B(n_1046),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1046),
.B(n_967),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1050),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_1018),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1037),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1077),
.B(n_1092),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_1037),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1090),
.Y(n_1196)
);

BUFx12f_ASAP7_75t_L g1197 ( 
.A(n_1090),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1001),
.B(n_1090),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1056),
.A2(n_1085),
.B(n_1061),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1092),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1066),
.A2(n_1082),
.B(n_1070),
.Y(n_1201)
);

OR2x6_ASAP7_75t_L g1202 ( 
.A(n_1092),
.B(n_1054),
.Y(n_1202)
);

BUFx4_ASAP7_75t_SL g1203 ( 
.A(n_972),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1060),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1067),
.A2(n_1074),
.B(n_1098),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1042),
.A2(n_1017),
.B1(n_1023),
.B2(n_1033),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1075),
.A2(n_1094),
.B(n_1076),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_1003),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_999),
.B(n_1049),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1010),
.A2(n_978),
.B(n_1035),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1025),
.A2(n_1088),
.B(n_1103),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1028),
.Y(n_1212)
);

NAND2x1p5_ASAP7_75t_L g1213 ( 
.A(n_976),
.B(n_987),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_992),
.A2(n_988),
.B(n_1065),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_964),
.B(n_1091),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1028),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_969),
.B(n_977),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_976),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_976),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_992),
.A2(n_940),
.B(n_988),
.C(n_1083),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_969),
.B(n_977),
.Y(n_1221)
);

INVx5_ASAP7_75t_L g1222 ( 
.A(n_1026),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1104),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1028),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1028),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_992),
.A2(n_988),
.B(n_1065),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_976),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1083),
.A2(n_940),
.B1(n_346),
.B2(n_327),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_969),
.B(n_977),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_992),
.A2(n_988),
.B(n_1065),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_961),
.B(n_526),
.Y(n_1231)
);

CKINVDCx11_ASAP7_75t_R g1232 ( 
.A(n_1104),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_1026),
.Y(n_1233)
);

O2A1O1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_992),
.A2(n_988),
.B(n_940),
.C(n_1065),
.Y(n_1234)
);

OR2x2_ASAP7_75t_L g1235 ( 
.A(n_979),
.B(n_964),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_SL g1236 ( 
.A1(n_961),
.A2(n_900),
.B1(n_1081),
.B2(n_1065),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_992),
.A2(n_1081),
.B1(n_1065),
.B2(n_988),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1104),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1105),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_964),
.Y(n_1240)
);

INVx4_ASAP7_75t_L g1241 ( 
.A(n_1144),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1236),
.A2(n_1231),
.B1(n_1133),
.B2(n_1154),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1110),
.A2(n_1111),
.B(n_1214),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1236),
.A2(n_1220),
.B1(n_1108),
.B2(n_1237),
.Y(n_1244)
);

AOI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1135),
.A2(n_1153),
.B(n_1122),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1160),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1223),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1132),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1148),
.Y(n_1249)
);

BUFx4f_ASAP7_75t_SL g1250 ( 
.A(n_1163),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1152),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1228),
.A2(n_1171),
.B1(n_1118),
.B2(n_1120),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1184),
.B(n_1181),
.Y(n_1253)
);

BUFx8_ASAP7_75t_L g1254 ( 
.A(n_1119),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1143),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1198),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1144),
.Y(n_1257)
);

OA21x2_ASAP7_75t_L g1258 ( 
.A1(n_1186),
.A2(n_1210),
.B(n_1155),
.Y(n_1258)
);

OAI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1133),
.A2(n_1235),
.B1(n_1118),
.B2(n_1240),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1131),
.B(n_1176),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1140),
.A2(n_1215),
.B1(n_1113),
.B2(n_1237),
.Y(n_1261)
);

AOI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1211),
.A2(n_1201),
.B(n_1205),
.Y(n_1262)
);

AOI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1207),
.A2(n_1199),
.B(n_1230),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1209),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1156),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1217),
.A2(n_1221),
.B1(n_1229),
.B2(n_1112),
.Y(n_1266)
);

BUFx2_ASAP7_75t_SL g1267 ( 
.A(n_1181),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1117),
.B(n_1217),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1126),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1183),
.A2(n_1136),
.B(n_1206),
.Y(n_1270)
);

NOR2x1_ASAP7_75t_SL g1271 ( 
.A(n_1172),
.B(n_1174),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1183),
.A2(n_1116),
.B(n_1226),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1128),
.B(n_1130),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1191),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1107),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1177),
.B(n_1174),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1123),
.Y(n_1277)
);

BUFx2_ASAP7_75t_SL g1278 ( 
.A(n_1222),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1138),
.B(n_1139),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1124),
.B(n_1125),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1147),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_1232),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1212),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1216),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1224),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1225),
.Y(n_1286)
);

INVx6_ASAP7_75t_L g1287 ( 
.A(n_1222),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1202),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1167),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1189),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_SL g1291 ( 
.A1(n_1157),
.A2(n_1115),
.B1(n_1149),
.B2(n_1141),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1234),
.A2(n_1117),
.B(n_1115),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1151),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1121),
.Y(n_1294)
);

CKINVDCx11_ASAP7_75t_R g1295 ( 
.A(n_1165),
.Y(n_1295)
);

AO21x1_ASAP7_75t_L g1296 ( 
.A1(n_1157),
.A2(n_1116),
.B(n_1159),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1204),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1159),
.A2(n_1158),
.B(n_1168),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1162),
.A2(n_1238),
.B1(n_1137),
.B2(n_1129),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1221),
.B(n_1229),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1180),
.A2(n_1175),
.B(n_1208),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1161),
.Y(n_1302)
);

OA21x2_ASAP7_75t_L g1303 ( 
.A1(n_1208),
.A2(n_1209),
.B(n_1168),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1238),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1175),
.A2(n_1134),
.B(n_1146),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1134),
.A2(n_1146),
.B(n_1196),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1150),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1142),
.A2(n_1219),
.B1(n_1218),
.B2(n_1233),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1164),
.B(n_1187),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1233),
.A2(n_1222),
.B1(n_1127),
.B2(n_1227),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1182),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1109),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1203),
.A2(n_1213),
.B(n_1178),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1200),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_1169),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1114),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1114),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1114),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1182),
.Y(n_1319)
);

BUFx2_ASAP7_75t_R g1320 ( 
.A(n_1173),
.Y(n_1320)
);

AOI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1188),
.A2(n_1194),
.B(n_1185),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1194),
.B(n_1179),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1169),
.Y(n_1323)
);

CKINVDCx6p67_ASAP7_75t_R g1324 ( 
.A(n_1145),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_SL g1325 ( 
.A1(n_1166),
.A2(n_1239),
.B1(n_1197),
.B2(n_1192),
.Y(n_1325)
);

INVx5_ASAP7_75t_L g1326 ( 
.A(n_1166),
.Y(n_1326)
);

OAI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1166),
.A2(n_1239),
.B1(n_1195),
.B2(n_1193),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_1170),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1170),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1195),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1177),
.B(n_1190),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1160),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1198),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1228),
.A2(n_1083),
.B1(n_940),
.B2(n_402),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1160),
.Y(n_1335)
);

AO21x1_ASAP7_75t_L g1336 ( 
.A1(n_1237),
.A2(n_1101),
.B(n_1081),
.Y(n_1336)
);

INVx11_ASAP7_75t_L g1337 ( 
.A(n_1119),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1228),
.A2(n_1083),
.B1(n_940),
.B2(n_402),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1160),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1231),
.A2(n_1083),
.B1(n_1101),
.B2(n_786),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1232),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1228),
.A2(n_1083),
.B1(n_940),
.B2(n_402),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_SL g1343 ( 
.A1(n_1236),
.A2(n_1101),
.B1(n_346),
.B2(n_327),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1220),
.A2(n_992),
.B(n_988),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1144),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1228),
.A2(n_1083),
.B1(n_940),
.B2(n_402),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1122),
.A2(n_1135),
.B(n_1153),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1297),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1243),
.A2(n_1244),
.B(n_1344),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1264),
.B(n_1260),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1247),
.Y(n_1351)
);

INVxp67_ASAP7_75t_SL g1352 ( 
.A(n_1256),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1331),
.B(n_1276),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1283),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1286),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1286),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1288),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1331),
.B(n_1276),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1268),
.B(n_1266),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1317),
.Y(n_1360)
);

OA21x2_ASAP7_75t_L g1361 ( 
.A1(n_1272),
.A2(n_1270),
.B(n_1245),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1303),
.Y(n_1362)
);

AOI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1262),
.A2(n_1263),
.B(n_1296),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1268),
.B(n_1300),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_1317),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1304),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1264),
.B(n_1260),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1280),
.B(n_1248),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1253),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1294),
.Y(n_1370)
);

AO21x2_ASAP7_75t_L g1371 ( 
.A1(n_1259),
.A2(n_1296),
.B(n_1298),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1318),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1302),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1250),
.Y(n_1374)
);

INVx1_ASAP7_75t_SL g1375 ( 
.A(n_1255),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1273),
.B(n_1279),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1280),
.B(n_1249),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_SL g1378 ( 
.A1(n_1336),
.A2(n_1292),
.B(n_1271),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1301),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1255),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1291),
.B(n_1290),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1288),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1318),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1293),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1251),
.B(n_1265),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1307),
.B(n_1275),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1277),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1284),
.B(n_1285),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1272),
.A2(n_1270),
.B(n_1336),
.Y(n_1389)
);

AOI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1347),
.A2(n_1258),
.B(n_1301),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1289),
.B(n_1242),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1256),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1333),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1333),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1274),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1337),
.Y(n_1396)
);

NOR2xp67_ASAP7_75t_SL g1397 ( 
.A(n_1278),
.B(n_1267),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1313),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1246),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1261),
.B(n_1298),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1254),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1332),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1335),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1298),
.B(n_1347),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1339),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1347),
.B(n_1329),
.Y(n_1406)
);

AO21x2_ASAP7_75t_L g1407 ( 
.A1(n_1340),
.A2(n_1321),
.B(n_1269),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1258),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1258),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1305),
.A2(n_1306),
.B(n_1312),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1316),
.Y(n_1411)
);

AO21x1_ASAP7_75t_SL g1412 ( 
.A1(n_1252),
.A2(n_1323),
.B(n_1319),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1329),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1320),
.B(n_1282),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1406),
.B(n_1315),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1364),
.B(n_1308),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1406),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1348),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1398),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1375),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1362),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1389),
.B(n_1315),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1351),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1387),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1389),
.B(n_1314),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1389),
.B(n_1311),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1359),
.B(n_1281),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1404),
.B(n_1350),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1404),
.B(n_1330),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1353),
.B(n_1299),
.Y(n_1430)
);

INVxp67_ASAP7_75t_SL g1431 ( 
.A(n_1352),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1353),
.B(n_1257),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1361),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1380),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1349),
.B(n_1281),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1367),
.B(n_1400),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_SL g1437 ( 
.A1(n_1378),
.A2(n_1343),
.B1(n_1346),
.B2(n_1342),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1370),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1358),
.B(n_1309),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1358),
.B(n_1392),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1392),
.Y(n_1441)
);

NOR2x1_ASAP7_75t_R g1442 ( 
.A(n_1396),
.B(n_1295),
.Y(n_1442)
);

AO21x2_ASAP7_75t_L g1443 ( 
.A1(n_1390),
.A2(n_1371),
.B(n_1363),
.Y(n_1443)
);

NOR4xp25_ASAP7_75t_SL g1444 ( 
.A(n_1397),
.B(n_1278),
.C(n_1287),
.D(n_1324),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1368),
.B(n_1241),
.Y(n_1445)
);

AO21x2_ASAP7_75t_L g1446 ( 
.A1(n_1371),
.A2(n_1322),
.B(n_1327),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1393),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1360),
.B(n_1326),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1377),
.B(n_1345),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1393),
.B(n_1394),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1361),
.B(n_1241),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1361),
.B(n_1241),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1394),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1408),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1438),
.B(n_1373),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1438),
.B(n_1416),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1416),
.B(n_1384),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1423),
.B(n_1366),
.Y(n_1458)
);

AOI221xp5_ASAP7_75t_L g1459 ( 
.A1(n_1437),
.A2(n_1381),
.B1(n_1338),
.B2(n_1334),
.C(n_1391),
.Y(n_1459)
);

OAI221xp5_ASAP7_75t_SL g1460 ( 
.A1(n_1437),
.A2(n_1425),
.B1(n_1439),
.B2(n_1434),
.C(n_1420),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1423),
.B(n_1385),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1428),
.B(n_1360),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1420),
.B(n_1414),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1428),
.B(n_1365),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_SL g1465 ( 
.A(n_1442),
.B(n_1401),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1428),
.B(n_1365),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1430),
.A2(n_1412),
.B1(n_1407),
.B2(n_1371),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1418),
.Y(n_1468)
);

AOI22x1_ASAP7_75t_SL g1469 ( 
.A1(n_1442),
.A2(n_1374),
.B1(n_1341),
.B2(n_1254),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1436),
.B(n_1372),
.Y(n_1470)
);

OAI211xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1450),
.A2(n_1376),
.B(n_1386),
.C(n_1409),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1427),
.B(n_1395),
.Y(n_1472)
);

NAND3xp33_ASAP7_75t_L g1473 ( 
.A(n_1425),
.B(n_1395),
.C(n_1388),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_L g1474 ( 
.A(n_1425),
.B(n_1408),
.C(n_1409),
.Y(n_1474)
);

AND2x2_ASAP7_75t_SL g1475 ( 
.A(n_1448),
.B(n_1369),
.Y(n_1475)
);

AOI221xp5_ASAP7_75t_L g1476 ( 
.A1(n_1426),
.A2(n_1378),
.B1(n_1403),
.B2(n_1399),
.C(n_1354),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1434),
.B(n_1372),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1440),
.B(n_1383),
.Y(n_1478)
);

AOI21xp33_ASAP7_75t_L g1479 ( 
.A1(n_1446),
.A2(n_1411),
.B(n_1379),
.Y(n_1479)
);

NOR3xp33_ASAP7_75t_L g1480 ( 
.A(n_1435),
.B(n_1310),
.C(n_1363),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1417),
.B(n_1383),
.Y(n_1481)
);

OAI21xp33_ASAP7_75t_L g1482 ( 
.A1(n_1431),
.A2(n_1383),
.B(n_1397),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1440),
.B(n_1439),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1439),
.B(n_1324),
.Y(n_1484)
);

NAND3xp33_ASAP7_75t_L g1485 ( 
.A(n_1435),
.B(n_1399),
.C(n_1403),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1417),
.B(n_1410),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1440),
.B(n_1295),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1432),
.B(n_1413),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1432),
.B(n_1354),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1431),
.B(n_1355),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1441),
.B(n_1355),
.Y(n_1491)
);

NAND3xp33_ASAP7_75t_L g1492 ( 
.A(n_1433),
.B(n_1405),
.C(n_1402),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1441),
.B(n_1447),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1429),
.B(n_1410),
.Y(n_1494)
);

NAND3xp33_ASAP7_75t_L g1495 ( 
.A(n_1422),
.B(n_1382),
.C(n_1357),
.Y(n_1495)
);

NAND3xp33_ASAP7_75t_L g1496 ( 
.A(n_1433),
.B(n_1405),
.C(n_1402),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1447),
.B(n_1356),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1494),
.B(n_1415),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1493),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1494),
.B(n_1415),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1486),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1468),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1491),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1486),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1497),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1468),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1490),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1456),
.B(n_1453),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1492),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1470),
.B(n_1451),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1483),
.B(n_1450),
.Y(n_1511)
);

INVxp67_ASAP7_75t_SL g1512 ( 
.A(n_1474),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1472),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1473),
.B(n_1453),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1474),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1489),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1492),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1455),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1461),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1475),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1457),
.B(n_1424),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1496),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1485),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1462),
.B(n_1452),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1475),
.Y(n_1525)
);

NOR2x1_ASAP7_75t_L g1526 ( 
.A(n_1485),
.B(n_1421),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1475),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1458),
.B(n_1454),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1464),
.B(n_1419),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1464),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1496),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1466),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1476),
.B(n_1424),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1521),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1530),
.B(n_1466),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1527),
.B(n_1495),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1516),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1523),
.B(n_1481),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1516),
.Y(n_1539)
);

NAND3xp33_ASAP7_75t_SL g1540 ( 
.A(n_1515),
.B(n_1482),
.C(n_1459),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1530),
.B(n_1481),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1515),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1528),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1502),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1533),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1530),
.B(n_1487),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1533),
.B(n_1478),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1502),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1528),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1530),
.B(n_1484),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1528),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1530),
.B(n_1482),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1518),
.B(n_1469),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1523),
.B(n_1426),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1508),
.B(n_1488),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1521),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1502),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1508),
.B(n_1477),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1527),
.B(n_1480),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1513),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1501),
.B(n_1445),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1518),
.B(n_1426),
.Y(n_1562)
);

NAND2x1_ASAP7_75t_L g1563 ( 
.A(n_1515),
.B(n_1526),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1513),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1502),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1514),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1503),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1503),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1506),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1511),
.B(n_1449),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1505),
.Y(n_1571)
);

AOI32xp33_ASAP7_75t_L g1572 ( 
.A1(n_1512),
.A2(n_1526),
.A3(n_1501),
.B1(n_1531),
.B2(n_1517),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1537),
.Y(n_1573)
);

AOI21xp33_ASAP7_75t_SL g1574 ( 
.A1(n_1572),
.A2(n_1514),
.B(n_1463),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1542),
.A2(n_1512),
.B1(n_1460),
.B2(n_1527),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1547),
.B(n_1555),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1542),
.A2(n_1527),
.B1(n_1520),
.B2(n_1525),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1537),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1539),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1539),
.Y(n_1580)
);

NAND2x1_ASAP7_75t_SL g1581 ( 
.A(n_1552),
.B(n_1527),
.Y(n_1581)
);

NAND2x1p5_ASAP7_75t_L g1582 ( 
.A(n_1563),
.B(n_1520),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1546),
.Y(n_1583)
);

AND2x2_ASAP7_75t_SL g1584 ( 
.A(n_1553),
.B(n_1465),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1546),
.B(n_1498),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1544),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1566),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1545),
.B(n_1507),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1550),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1547),
.B(n_1511),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1560),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1560),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1550),
.B(n_1498),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1561),
.B(n_1498),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1540),
.B(n_1469),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1534),
.B(n_1556),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1564),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1561),
.B(n_1500),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1536),
.B(n_1520),
.Y(n_1599)
);

NOR2xp67_ASAP7_75t_L g1600 ( 
.A(n_1552),
.B(n_1525),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1563),
.A2(n_1525),
.B1(n_1514),
.B2(n_1501),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1554),
.A2(n_1532),
.B1(n_1529),
.B2(n_1511),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1559),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1559),
.A2(n_1467),
.B1(n_1517),
.B2(n_1509),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1559),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1555),
.B(n_1507),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1564),
.B(n_1499),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1567),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1567),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1536),
.B(n_1504),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1571),
.Y(n_1611)
);

OAI33xp33_ASAP7_75t_L g1612 ( 
.A1(n_1543),
.A2(n_1531),
.A3(n_1517),
.B1(n_1509),
.B2(n_1522),
.B3(n_1499),
.Y(n_1612)
);

INVxp67_ASAP7_75t_SL g1613 ( 
.A(n_1538),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1568),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1568),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1586),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1612),
.A2(n_1509),
.B1(n_1522),
.B2(n_1517),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1582),
.B(n_1536),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1582),
.B(n_1594),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1605),
.B(n_1543),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1586),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1573),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1584),
.B(n_1574),
.Y(n_1623)
);

NOR2x1_ASAP7_75t_L g1624 ( 
.A(n_1595),
.B(n_1571),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1598),
.B(n_1549),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1576),
.B(n_1549),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1612),
.A2(n_1522),
.B1(n_1412),
.B2(n_1419),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1578),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1595),
.B(n_1337),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1584),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1606),
.B(n_1551),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1606),
.B(n_1551),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1585),
.B(n_1593),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1590),
.B(n_1558),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1610),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1583),
.B(n_1535),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1587),
.Y(n_1637)
);

INVx4_ASAP7_75t_L g1638 ( 
.A(n_1605),
.Y(n_1638)
);

NOR2x1_ASAP7_75t_L g1639 ( 
.A(n_1575),
.B(n_1558),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1610),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1587),
.B(n_1505),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1610),
.B(n_1535),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1603),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1589),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1581),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1599),
.B(n_1541),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1613),
.B(n_1562),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1613),
.B(n_1519),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1579),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1580),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1588),
.B(n_1570),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1643),
.B(n_1604),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1643),
.B(n_1596),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1637),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1637),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1644),
.B(n_1591),
.Y(n_1656)
);

OAI322xp33_ASAP7_75t_L g1657 ( 
.A1(n_1623),
.A2(n_1601),
.A3(n_1577),
.B1(n_1611),
.B2(n_1609),
.C1(n_1608),
.C2(n_1597),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1634),
.B(n_1607),
.Y(n_1658)
);

NOR3xp33_ASAP7_75t_L g1659 ( 
.A(n_1624),
.B(n_1614),
.C(n_1592),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1638),
.B(n_1600),
.Y(n_1660)
);

INVx1_ASAP7_75t_SL g1661 ( 
.A(n_1630),
.Y(n_1661)
);

OAI22xp33_ASAP7_75t_SL g1662 ( 
.A1(n_1630),
.A2(n_1599),
.B1(n_1615),
.B2(n_1602),
.Y(n_1662)
);

NAND2xp33_ASAP7_75t_SL g1663 ( 
.A(n_1618),
.B(n_1599),
.Y(n_1663)
);

AOI221xp5_ASAP7_75t_L g1664 ( 
.A1(n_1617),
.A2(n_1504),
.B1(n_1471),
.B2(n_1479),
.C(n_1557),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1622),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1638),
.B(n_1254),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1633),
.B(n_1541),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1644),
.B(n_1519),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1633),
.B(n_1500),
.Y(n_1669)
);

NAND2x1_ASAP7_75t_L g1670 ( 
.A(n_1618),
.B(n_1645),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1624),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1642),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1645),
.B(n_1529),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1644),
.B(n_1570),
.Y(n_1674)
);

INVx1_ASAP7_75t_SL g1675 ( 
.A(n_1635),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1639),
.A2(n_1443),
.B1(n_1433),
.B2(n_1557),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1661),
.B(n_1633),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1675),
.B(n_1672),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1676),
.A2(n_1639),
.B1(n_1627),
.B2(n_1645),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1654),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1671),
.B(n_1638),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1663),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1664),
.A2(n_1616),
.B1(n_1621),
.B2(n_1647),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_1670),
.Y(n_1684)
);

OAI21xp33_ASAP7_75t_L g1685 ( 
.A1(n_1662),
.A2(n_1632),
.B(n_1631),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1666),
.B(n_1638),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1671),
.B(n_1620),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_1666),
.Y(n_1688)
);

NOR2xp67_ASAP7_75t_L g1689 ( 
.A(n_1660),
.B(n_1635),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1667),
.B(n_1620),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1669),
.B(n_1642),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1652),
.B(n_1620),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1676),
.A2(n_1621),
.B1(n_1616),
.B2(n_1647),
.Y(n_1693)
);

BUFx2_ASAP7_75t_L g1694 ( 
.A(n_1660),
.Y(n_1694)
);

NOR2x1_ASAP7_75t_L g1695 ( 
.A(n_1655),
.B(n_1629),
.Y(n_1695)
);

OAI221xp5_ASAP7_75t_L g1696 ( 
.A1(n_1679),
.A2(n_1659),
.B1(n_1653),
.B2(n_1632),
.C(n_1631),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_SL g1697 ( 
.A(n_1692),
.B(n_1618),
.Y(n_1697)
);

NOR3xp33_ASAP7_75t_L g1698 ( 
.A(n_1688),
.B(n_1659),
.C(n_1657),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1685),
.A2(n_1658),
.B(n_1656),
.C(n_1665),
.Y(n_1699)
);

NAND4xp75_ASAP7_75t_L g1700 ( 
.A(n_1695),
.B(n_1673),
.C(n_1640),
.D(n_1635),
.Y(n_1700)
);

AOI21xp33_ASAP7_75t_L g1701 ( 
.A1(n_1684),
.A2(n_1621),
.B(n_1616),
.Y(n_1701)
);

OAI322xp33_ASAP7_75t_L g1702 ( 
.A1(n_1680),
.A2(n_1640),
.A3(n_1674),
.B1(n_1668),
.B2(n_1648),
.C1(n_1641),
.C2(n_1649),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1682),
.B(n_1640),
.Y(n_1703)
);

AOI211xp5_ASAP7_75t_L g1704 ( 
.A1(n_1689),
.A2(n_1620),
.B(n_1619),
.C(n_1649),
.Y(n_1704)
);

AOI221xp5_ASAP7_75t_L g1705 ( 
.A1(n_1683),
.A2(n_1648),
.B1(n_1650),
.B2(n_1628),
.C(n_1622),
.Y(n_1705)
);

AOI221xp5_ASAP7_75t_L g1706 ( 
.A1(n_1693),
.A2(n_1678),
.B1(n_1680),
.B2(n_1677),
.C(n_1687),
.Y(n_1706)
);

AND5x1_ASAP7_75t_L g1707 ( 
.A(n_1706),
.B(n_1686),
.C(n_1694),
.D(n_1690),
.E(n_1681),
.Y(n_1707)
);

O2A1O1Ixp33_ASAP7_75t_L g1708 ( 
.A1(n_1698),
.A2(n_1699),
.B(n_1703),
.C(n_1696),
.Y(n_1708)
);

NOR2xp67_ASAP7_75t_L g1709 ( 
.A(n_1697),
.B(n_1691),
.Y(n_1709)
);

NOR3xp33_ASAP7_75t_L g1710 ( 
.A(n_1701),
.B(n_1700),
.C(n_1702),
.Y(n_1710)
);

NOR2x1_ASAP7_75t_L g1711 ( 
.A(n_1704),
.B(n_1628),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1705),
.B(n_1634),
.Y(n_1712)
);

INVxp67_ASAP7_75t_L g1713 ( 
.A(n_1703),
.Y(n_1713)
);

AND5x1_ASAP7_75t_L g1714 ( 
.A(n_1706),
.B(n_1642),
.C(n_1619),
.D(n_1646),
.E(n_1626),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1698),
.B(n_1636),
.Y(n_1715)
);

NOR3xp33_ASAP7_75t_L g1716 ( 
.A(n_1708),
.B(n_1710),
.C(n_1713),
.Y(n_1716)
);

AND3x1_ASAP7_75t_L g1717 ( 
.A(n_1715),
.B(n_1619),
.C(n_1646),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1711),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1712),
.B(n_1626),
.Y(n_1719)
);

INVxp67_ASAP7_75t_SL g1720 ( 
.A(n_1707),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1718),
.Y(n_1721)
);

NOR2x1_ASAP7_75t_L g1722 ( 
.A(n_1719),
.B(n_1709),
.Y(n_1722)
);

AOI31xp33_ASAP7_75t_L g1723 ( 
.A1(n_1720),
.A2(n_1714),
.A3(n_1646),
.B(n_1650),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1717),
.Y(n_1724)
);

INVxp67_ASAP7_75t_SL g1725 ( 
.A(n_1716),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1717),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1725),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1722),
.Y(n_1728)
);

NAND5xp2_ASAP7_75t_L g1729 ( 
.A(n_1724),
.B(n_1726),
.C(n_1723),
.D(n_1721),
.E(n_1636),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1723),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1726),
.A2(n_1641),
.B1(n_1651),
.B2(n_1625),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1728),
.Y(n_1732)
);

AOI22x1_ASAP7_75t_L g1733 ( 
.A1(n_1730),
.A2(n_1625),
.B1(n_1651),
.B2(n_1510),
.Y(n_1733)
);

INVx3_ASAP7_75t_SL g1734 ( 
.A(n_1727),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1732),
.Y(n_1735)
);

OAI221xp5_ASAP7_75t_L g1736 ( 
.A1(n_1735),
.A2(n_1734),
.B1(n_1731),
.B2(n_1733),
.C(n_1729),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1736),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1736),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1738),
.A2(n_1731),
.B1(n_1625),
.B2(n_1544),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1737),
.B(n_1548),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1740),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1739),
.A2(n_1565),
.B(n_1548),
.Y(n_1742)
);

AOI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1741),
.A2(n_1565),
.B(n_1569),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1743),
.A2(n_1742),
.B1(n_1569),
.B2(n_1443),
.Y(n_1744)
);

OAI221xp5_ASAP7_75t_R g1745 ( 
.A1(n_1744),
.A2(n_1444),
.B1(n_1328),
.B2(n_1325),
.C(n_1524),
.Y(n_1745)
);

AOI211xp5_ASAP7_75t_L g1746 ( 
.A1(n_1745),
.A2(n_1444),
.B(n_1345),
.C(n_1257),
.Y(n_1746)
);


endmodule