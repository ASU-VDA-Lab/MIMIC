module fake_jpeg_11097_n_107 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_10),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_32),
.Y(n_45)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_0),
.B(n_1),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_23),
.B1(n_19),
.B2(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_3),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_34),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_34),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_25),
.A2(n_22),
.B1(n_23),
.B2(n_19),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_26),
.B1(n_29),
.B2(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_18),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_14),
.B1(n_18),
.B2(n_11),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_45),
.B1(n_12),
.B2(n_13),
.Y(n_62)
);

OR2x2_ASAP7_75t_SL g46 ( 
.A(n_24),
.B(n_2),
.Y(n_46)
);

NOR2xp67_ASAP7_75t_R g54 ( 
.A(n_46),
.B(n_16),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_34),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_54),
.B(n_60),
.Y(n_67)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_52),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_61),
.B1(n_51),
.B2(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_58),
.Y(n_65)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_13),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_16),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_12),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_46),
.B1(n_17),
.B2(n_43),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_17),
.B(n_27),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_48),
.C(n_37),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_27),
.B1(n_43),
.B2(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_62),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_49),
.B1(n_63),
.B2(n_57),
.Y(n_78)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_78),
.B(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_50),
.C(n_56),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_67),
.C(n_65),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_83),
.C(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_65),
.B(n_54),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_81),
.C(n_80),
.Y(n_92)
);

AO221x1_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_88),
.B1(n_74),
.B2(n_79),
.C(n_76),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_67),
.B(n_73),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_71),
.B1(n_69),
.B2(n_75),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_95),
.Y(n_97)
);

BUFx24_ASAP7_75t_SL g93 ( 
.A(n_85),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_93),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_68),
.C(n_60),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_90),
.C(n_86),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_47),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_6),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_102),
.Y(n_104)
);

NAND5xp2_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_6),
.C(n_7),
.D(n_8),
.E(n_96),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_100),
.B(n_98),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_103),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_7),
.Y(n_107)
);


endmodule