module fake_ibex_2036_n_2939 (n_151, n_85, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_545, n_194, n_249, n_334, n_312, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_531, n_15, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_527, n_465, n_48, n_325, n_57, n_301, n_496, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_13, n_122, n_523, n_116, n_370, n_431, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_490, n_52, n_448, n_99, n_466, n_269, n_156, n_126, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_536, n_352, n_290, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_514, n_429, n_275, n_541, n_98, n_129, n_267, n_245, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_66, n_305, n_307, n_192, n_140, n_484, n_480, n_416, n_365, n_4, n_6, n_539, n_100, n_179, n_354, n_206, n_392, n_516, n_548, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_546, n_199, n_495, n_410, n_308, n_463, n_411, n_135, n_520, n_512, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_517, n_211, n_218, n_314, n_132, n_277, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_532, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_476, n_461, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_311, n_406, n_97, n_197, n_528, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_425, n_2939);

input n_151;
input n_85;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_194;
input n_249;
input n_334;
input n_312;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_531;
input n_15;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_523;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_490;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_126;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_536;
input n_352;
input n_290;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_514;
input n_429;
input n_275;
input n_541;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_480;
input n_416;
input n_365;
input n_4;
input n_6;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_516;
input n_548;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_546;
input n_199;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_520;
input n_512;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_476;
input n_461;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2939;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_2569;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_1079;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1954;
wire n_1859;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_1308;
wire n_556;
wire n_1138;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_884;
wire n_667;
wire n_2396;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2724;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_557;
wire n_641;
wire n_1937;
wire n_2311;
wire n_893;
wire n_1654;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_852;
wire n_1427;
wire n_1133;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2814;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2922;
wire n_2347;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1960;
wire n_1723;
wire n_2663;
wire n_793;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_2906;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_554;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_605;
wire n_2373;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_971;
wire n_1326;
wire n_702;
wire n_1350;
wire n_906;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_2541;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_2723;
wire n_1616;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_2256;
wire n_606;
wire n_737;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2879;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2718;
wire n_2377;
wire n_2577;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_2573;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_591;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_2838;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_594;
wire n_2361;
wire n_1566;
wire n_1464;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_660;
wire n_2590;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_576;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_607;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2823;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_2905;
wire n_803;
wire n_2570;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_2095;
wire n_555;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_2903;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_2463;
wire n_2654;
wire n_717;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_668;
wire n_871;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_588;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_916;
wire n_2298;
wire n_2771;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_2772;
wire n_2778;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1845;
wire n_1104;
wire n_1667;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_626;
wire n_1941;
wire n_1707;
wire n_2422;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_634;
wire n_961;
wire n_991;
wire n_1331;
wire n_1349;
wire n_1223;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_2862;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_598;
wire n_2141;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_2920;
wire n_604;
wire n_1598;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_1625;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2555;
wire n_2639;
wire n_2330;
wire n_636;
wire n_1259;
wire n_2108;
wire n_2535;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2709;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_2665;
wire n_1124;
wire n_611;
wire n_1690;
wire n_2688;
wire n_2881;
wire n_1673;
wire n_2018;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_2758;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_648;
wire n_571;
wire n_1169;
wire n_1946;
wire n_1726;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_2447;
wire n_2818;
wire n_1057;
wire n_1473;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_775;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_1167;
wire n_818;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_2608;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2861;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_1256;
wire n_2798;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_1961;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_688;
wire n_1547;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1542;
wire n_1097;
wire n_2518;
wire n_2784;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_1147;
wire n_747;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_1029;
wire n_2394;
wire n_770;
wire n_1635;
wire n_1572;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_2323;
wire n_740;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_1986;
wire n_2882;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_2734;
wire n_2870;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_580;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2928;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_999;
wire n_2634;
wire n_1092;
wire n_1808;
wire n_560;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_2931;
wire n_2492;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_1142;
wire n_783;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2357;
wire n_2303;
wire n_2653;
wire n_2855;
wire n_2618;
wire n_924;
wire n_2937;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_2092;
wire n_566;
wire n_581;
wire n_1365;
wire n_1472;
wire n_2443;
wire n_2802;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2704;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_1736;
wire n_2907;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_2754;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1947;
wire n_1675;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_908;
wire n_1346;
wire n_565;
wire n_2834;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_529),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_8),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_342),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_280),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_358),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_297),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_434),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_179),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_408),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_353),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_63),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_387),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_84),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_232),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_12),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_420),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_6),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_39),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_334),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_311),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_548),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_186),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_553),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_478),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_451),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_481),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_521),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_319),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_471),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_528),
.B(n_403),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_106),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_550),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_183),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_172),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_345),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_27),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_35),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_231),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_67),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_511),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_136),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_243),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_543),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_173),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_204),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_17),
.Y(n_599)
);

NOR2xp67_ASAP7_75t_L g600 ( 
.A(n_116),
.B(n_314),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_306),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_482),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_527),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_462),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_477),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_36),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_40),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_486),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_416),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_476),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_519),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_356),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_183),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_11),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_541),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_391),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_383),
.Y(n_617)
);

NOR2xp67_ASAP7_75t_L g618 ( 
.A(n_228),
.B(n_195),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_208),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_115),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_419),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_307),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_233),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_208),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_522),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_84),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_542),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_178),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_516),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_544),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_401),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_309),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_322),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_549),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_213),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_427),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_538),
.Y(n_637)
);

BUFx5_ASAP7_75t_L g638 ( 
.A(n_520),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_295),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_335),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_325),
.Y(n_641)
);

NOR2xp67_ASAP7_75t_L g642 ( 
.A(n_66),
.B(n_356),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_479),
.Y(n_643)
);

BUFx10_ASAP7_75t_L g644 ( 
.A(n_37),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_381),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_152),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_272),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_111),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_119),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_499),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_97),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_483),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_342),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_245),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_58),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_420),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_89),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_16),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_151),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_47),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_337),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_15),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_170),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_408),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_143),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_169),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_390),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_255),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_385),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_79),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_313),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_531),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_371),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_274),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_23),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_552),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_14),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_517),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_159),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_251),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_256),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_258),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_269),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_147),
.Y(n_684)
);

NOR2xp67_ASAP7_75t_L g685 ( 
.A(n_248),
.B(n_82),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_235),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_324),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_459),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_489),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_321),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_364),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_498),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_272),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_10),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_305),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_526),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_307),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_260),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_36),
.Y(n_699)
);

BUFx5_ASAP7_75t_L g700 ( 
.A(n_237),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_40),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_118),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_515),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_247),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_340),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_184),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_14),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_535),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_537),
.B(n_360),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_107),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_458),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_370),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_174),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_104),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_259),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_438),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_319),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_132),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_376),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_368),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_385),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_101),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_378),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_300),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_114),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_269),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_79),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_152),
.Y(n_728)
);

BUFx10_ASAP7_75t_L g729 ( 
.A(n_258),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_396),
.B(n_71),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_547),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_524),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_508),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_423),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_190),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_410),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_370),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_72),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_93),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_422),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_523),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_98),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_171),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_90),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_125),
.Y(n_745)
);

NOR2xp67_ASAP7_75t_L g746 ( 
.A(n_44),
.B(n_267),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_386),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_469),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_372),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_386),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_209),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_160),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_427),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_382),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_525),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_492),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_192),
.Y(n_757)
);

CKINVDCx14_ASAP7_75t_R g758 ( 
.A(n_493),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_322),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_197),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_205),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_391),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_233),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_435),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_488),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_70),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_257),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_291),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_480),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_0),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_354),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_394),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_214),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_184),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_6),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_96),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_445),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_545),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_514),
.Y(n_779)
);

CKINVDCx16_ASAP7_75t_R g780 ( 
.A(n_56),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_347),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_289),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_407),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_120),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_293),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_290),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_490),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_257),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_433),
.B(n_97),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_362),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_167),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_464),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_176),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_232),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_277),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_122),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_63),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_396),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_225),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_414),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_323),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_167),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_88),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_44),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_447),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_165),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_402),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_536),
.Y(n_808)
);

CKINVDCx16_ASAP7_75t_R g809 ( 
.A(n_207),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_372),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_203),
.Y(n_811)
);

NOR2xp67_ASAP7_75t_L g812 ( 
.A(n_9),
.B(n_155),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_238),
.Y(n_813)
);

CKINVDCx16_ASAP7_75t_R g814 ( 
.A(n_518),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_435),
.Y(n_815)
);

CKINVDCx16_ASAP7_75t_R g816 ( 
.A(n_211),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_491),
.B(n_77),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_42),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_80),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_69),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_509),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_290),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_76),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_271),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_357),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_237),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_7),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_546),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_229),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_266),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_175),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_127),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_90),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_28),
.Y(n_834)
);

BUFx2_ASAP7_75t_SL g835 ( 
.A(n_513),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_101),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_70),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_451),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_265),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_77),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_446),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_397),
.Y(n_842)
);

CKINVDCx16_ASAP7_75t_R g843 ( 
.A(n_105),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_50),
.Y(n_844)
);

NOR2xp67_ASAP7_75t_L g845 ( 
.A(n_359),
.B(n_401),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_414),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_475),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_128),
.Y(n_848)
);

BUFx10_ASAP7_75t_L g849 ( 
.A(n_423),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_410),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_146),
.Y(n_851)
);

BUFx8_ASAP7_75t_SL g852 ( 
.A(n_164),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_217),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_0),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_443),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_51),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_185),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_242),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_61),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_512),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_81),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_324),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_135),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_234),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_551),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_380),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_198),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_303),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_104),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_201),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_31),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_455),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_470),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_227),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_323),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_366),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_83),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_35),
.Y(n_878)
);

INVxp67_ASAP7_75t_L g879 ( 
.A(n_12),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_392),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_265),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_438),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_82),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_220),
.Y(n_884)
);

BUFx8_ASAP7_75t_SL g885 ( 
.A(n_421),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_106),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_436),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_507),
.Y(n_888)
);

BUFx5_ASAP7_75t_L g889 ( 
.A(n_116),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_534),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_102),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_68),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_298),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_400),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_343),
.Y(n_895)
);

NOR2xp67_ASAP7_75t_L g896 ( 
.A(n_219),
.B(n_140),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_510),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_150),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_504),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_487),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_456),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_263),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_127),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_813),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_644),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_700),
.Y(n_906)
);

OAI22x1_ASAP7_75t_R g907 ( 
.A1(n_562),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_700),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_694),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_813),
.B(n_2),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_700),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_696),
.B(n_3),
.Y(n_912)
);

BUFx8_ASAP7_75t_SL g913 ( 
.A(n_852),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_611),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_611),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_611),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_607),
.B(n_4),
.Y(n_917)
);

CKINVDCx16_ASAP7_75t_R g918 ( 
.A(n_780),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_611),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_607),
.B(n_4),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_876),
.Y(n_921)
);

INVx5_ASAP7_75t_L g922 ( 
.A(n_676),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_700),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_786),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_876),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_903),
.B(n_5),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_814),
.Y(n_927)
);

OA21x2_ASAP7_75t_L g928 ( 
.A1(n_604),
.A2(n_460),
.B(n_457),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_903),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_571),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_571),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_644),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_638),
.B(n_5),
.Y(n_933)
);

BUFx8_ASAP7_75t_L g934 ( 
.A(n_700),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_809),
.B(n_7),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_644),
.Y(n_936)
);

BUFx8_ASAP7_75t_L g937 ( 
.A(n_700),
.Y(n_937)
);

BUFx12f_ASAP7_75t_L g938 ( 
.A(n_729),
.Y(n_938)
);

AOI22x1_ASAP7_75t_SL g939 ( 
.A1(n_562),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_563),
.B(n_11),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_700),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_565),
.B(n_13),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_567),
.B(n_15),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_SL g944 ( 
.A1(n_566),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_944)
);

BUFx12f_ASAP7_75t_L g945 ( 
.A(n_729),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_634),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_683),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_889),
.Y(n_948)
);

BUFx8_ASAP7_75t_L g949 ( 
.A(n_889),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_590),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_889),
.Y(n_951)
);

INVx5_ASAP7_75t_L g952 ( 
.A(n_676),
.Y(n_952)
);

BUFx8_ASAP7_75t_SL g953 ( 
.A(n_852),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_590),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_816),
.A2(n_843),
.B1(n_556),
.B2(n_558),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_669),
.B(n_19),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_669),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_634),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_885),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_889),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_675),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_675),
.Y(n_962)
);

INVx5_ASAP7_75t_L g963 ( 
.A(n_676),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_634),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_729),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_638),
.B(n_20),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_889),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_570),
.B(n_20),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_573),
.B(n_21),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_575),
.B(n_21),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_634),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_603),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_698),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_643),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_643),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_735),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_643),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_889),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_581),
.B(n_22),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_735),
.Y(n_980)
);

NOR2x1_ASAP7_75t_L g981 ( 
.A(n_805),
.B(n_461),
.Y(n_981)
);

BUFx8_ASAP7_75t_SL g982 ( 
.A(n_885),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_849),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_643),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_566),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_805),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_860),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_588),
.B(n_22),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_592),
.B(n_24),
.Y(n_989)
);

INVx6_ASAP7_75t_L g990 ( 
.A(n_849),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_838),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_838),
.Y(n_992)
);

BUFx8_ASAP7_75t_SL g993 ( 
.A(n_589),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_599),
.B(n_601),
.Y(n_994)
);

AND2x6_ASAP7_75t_L g995 ( 
.A(n_732),
.B(n_463),
.Y(n_995)
);

OA21x2_ASAP7_75t_L g996 ( 
.A1(n_604),
.A2(n_466),
.B(n_465),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_869),
.B(n_24),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_860),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_849),
.B(n_25),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_869),
.B(n_25),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_574),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_638),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_785),
.B(n_26),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_758),
.B(n_26),
.Y(n_1004)
);

BUFx12f_ASAP7_75t_L g1005 ( 
.A(n_556),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_638),
.Y(n_1006)
);

AND2x6_ASAP7_75t_L g1007 ( 
.A(n_732),
.B(n_467),
.Y(n_1007)
);

AND2x2_ASAP7_75t_SL g1008 ( 
.A(n_817),
.B(n_468),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_879),
.B(n_27),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_890),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_947),
.B(n_557),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_914),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_922),
.B(n_952),
.Y(n_1013)
);

AO21x2_ASAP7_75t_L g1014 ( 
.A1(n_933),
.A2(n_580),
.B(n_577),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_934),
.B(n_625),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_934),
.B(n_625),
.Y(n_1016)
);

NAND2xp33_ASAP7_75t_L g1017 ( 
.A(n_995),
.B(n_638),
.Y(n_1017)
);

NAND3xp33_ASAP7_75t_L g1018 ( 
.A(n_937),
.B(n_902),
.C(n_558),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_910),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_922),
.B(n_596),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_906),
.Y(n_1021)
);

AND3x2_ASAP7_75t_L g1022 ( 
.A(n_909),
.B(n_657),
.C(n_730),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_922),
.B(n_578),
.Y(n_1023)
);

INVx8_ASAP7_75t_L g1024 ( 
.A(n_922),
.Y(n_1024)
);

CKINVDCx6p67_ASAP7_75t_R g1025 ( 
.A(n_918),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_910),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_952),
.B(n_689),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_911),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_952),
.B(n_578),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_952),
.B(n_963),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_917),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_937),
.B(n_637),
.Y(n_1032)
);

AOI21x1_ASAP7_75t_L g1033 ( 
.A1(n_908),
.A2(n_672),
.B(n_637),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_924),
.B(n_586),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_923),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_1005),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_941),
.Y(n_1037)
);

OR2x6_ASAP7_75t_L g1038 ( 
.A(n_938),
.B(n_600),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_926),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_913),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_963),
.B(n_586),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_956),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_949),
.B(n_672),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_956),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_990),
.B(n_932),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_990),
.B(n_598),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_948),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_951),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_997),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_990),
.B(n_598),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_1008),
.A2(n_955),
.B1(n_1000),
.B2(n_997),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_1000),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_963),
.B(n_587),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_963),
.B(n_587),
.Y(n_1054)
);

NAND3xp33_ASAP7_75t_L g1055 ( 
.A(n_949),
.B(n_902),
.C(n_594),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_932),
.B(n_591),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_960),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_967),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_SL g1059 ( 
.A(n_1008),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_SL g1060 ( 
.A1(n_985),
.A2(n_613),
.B1(n_632),
.B2(n_589),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_904),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_921),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_925),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_1002),
.B(n_678),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_927),
.A2(n_828),
.B1(n_610),
.B2(n_594),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_978),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_914),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1006),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_914),
.Y(n_1069)
);

AND3x2_ASAP7_75t_L g1070 ( 
.A(n_935),
.B(n_614),
.C(n_606),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_1001),
.B(n_678),
.Y(n_1071)
);

INVx8_ASAP7_75t_L g1072 ( 
.A(n_945),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_929),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1010),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_904),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_914),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_920),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_965),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_965),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_913),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_983),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_930),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_915),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_915),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_931),
.Y(n_1085)
);

INVx5_ASAP7_75t_L g1086 ( 
.A(n_995),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_983),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_905),
.B(n_591),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_1001),
.B(n_692),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_953),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_915),
.Y(n_1091)
);

NAND2xp33_ASAP7_75t_L g1092 ( 
.A(n_995),
.B(n_638),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_936),
.B(n_692),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_959),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_950),
.B(n_847),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_915),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_981),
.B(n_847),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_953),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_954),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_982),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_957),
.Y(n_1101)
);

INVxp33_ASAP7_75t_L g1102 ( 
.A(n_999),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_916),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_916),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1004),
.B(n_595),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_961),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_962),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_916),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_973),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_972),
.B(n_638),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_976),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_980),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_919),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_912),
.A2(n_874),
.B1(n_884),
.B2(n_597),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_986),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_994),
.B(n_884),
.Y(n_1116)
);

CKINVDCx11_ASAP7_75t_R g1117 ( 
.A(n_985),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_919),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_991),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_992),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_940),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_940),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_919),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_942),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_994),
.B(n_886),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_972),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_942),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_989),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_919),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_946),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_982),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_943),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_946),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_943),
.Y(n_1134)
);

NAND2xp33_ASAP7_75t_L g1135 ( 
.A(n_995),
.B(n_890),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1003),
.B(n_874),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_946),
.Y(n_1137)
);

INVxp33_ASAP7_75t_L g1138 ( 
.A(n_993),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_958),
.Y(n_1139)
);

AND2x6_ASAP7_75t_L g1140 ( 
.A(n_995),
.B(n_582),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_968),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1003),
.B(n_886),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1009),
.B(n_892),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_968),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_1007),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_SL g1146 ( 
.A(n_1007),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_958),
.Y(n_1147)
);

NAND3xp33_ASAP7_75t_L g1148 ( 
.A(n_1009),
.B(n_893),
.C(n_892),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_969),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_970),
.B(n_893),
.Y(n_1150)
);

AOI21x1_ASAP7_75t_L g1151 ( 
.A1(n_928),
.A2(n_602),
.B(n_593),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_970),
.B(n_605),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_979),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_979),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_964),
.Y(n_1155)
);

OR2x6_ASAP7_75t_L g1156 ( 
.A(n_944),
.B(n_618),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_993),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_988),
.B(n_615),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_988),
.B(n_630),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_966),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_971),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_971),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1007),
.B(n_895),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_939),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_996),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_971),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_996),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_974),
.Y(n_1168)
);

AO22x2_ASAP7_75t_L g1169 ( 
.A1(n_907),
.A2(n_789),
.B1(n_651),
.B2(n_656),
.Y(n_1169)
);

NAND2xp33_ASAP7_75t_L g1170 ( 
.A(n_974),
.B(n_890),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_974),
.B(n_650),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_974),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_975),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_975),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_998),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_998),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_975),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_977),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_977),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_977),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_984),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_998),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_984),
.Y(n_1183)
);

BUFx10_ASAP7_75t_L g1184 ( 
.A(n_984),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_984),
.B(n_652),
.Y(n_1185)
);

OAI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_987),
.A2(n_613),
.B1(n_682),
.B2(n_632),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1126),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1144),
.B(n_554),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1077),
.B(n_576),
.Y(n_1189)
);

INVxp67_ASAP7_75t_L g1190 ( 
.A(n_1154),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1121),
.B(n_576),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1154),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1061),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1122),
.B(n_579),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1124),
.B(n_579),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1061),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1086),
.B(n_585),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1062),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1126),
.Y(n_1199)
);

NAND2xp33_ASAP7_75t_L g1200 ( 
.A(n_1140),
.B(n_585),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1063),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1127),
.B(n_610),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1073),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1051),
.A2(n_828),
.B1(n_726),
.B2(n_734),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1132),
.B(n_873),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1086),
.B(n_873),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1134),
.B(n_1141),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_1072),
.Y(n_1208)
);

NAND2xp33_ASAP7_75t_L g1209 ( 
.A(n_1140),
.B(n_888),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1145),
.Y(n_1210)
);

NAND2xp33_ASAP7_75t_L g1211 ( 
.A(n_1140),
.B(n_897),
.Y(n_1211)
);

INVxp67_ASAP7_75t_L g1212 ( 
.A(n_1011),
.Y(n_1212)
);

NOR3xp33_ASAP7_75t_L g1213 ( 
.A(n_1186),
.B(n_569),
.C(n_561),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1149),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1116),
.B(n_895),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1153),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1150),
.B(n_897),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1026),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1081),
.B(n_899),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1026),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1056),
.B(n_642),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1081),
.B(n_899),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1087),
.B(n_733),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1125),
.B(n_608),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1087),
.B(n_787),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1158),
.B(n_627),
.Y(n_1226)
);

BUFx8_ASAP7_75t_L g1227 ( 
.A(n_1098),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1158),
.B(n_629),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1075),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_1034),
.B(n_898),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1120),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1128),
.B(n_898),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1033),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1031),
.A2(n_622),
.B(n_623),
.C(n_621),
.Y(n_1234)
);

AOI221xp5_ASAP7_75t_L g1235 ( 
.A1(n_1169),
.A2(n_635),
.B1(n_636),
.B2(n_633),
.C(n_628),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1052),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1082),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1039),
.B(n_688),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1018),
.B(n_703),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1078),
.B(n_900),
.Y(n_1240)
);

NOR2xp67_ASAP7_75t_L g1241 ( 
.A(n_1157),
.B(n_29),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1052),
.Y(n_1242)
);

INVxp67_ASAP7_75t_L g1243 ( 
.A(n_1065),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1042),
.A2(n_641),
.B1(n_645),
.B2(n_639),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1085),
.Y(n_1245)
);

OR2x2_ASAP7_75t_L g1246 ( 
.A(n_1072),
.B(n_1036),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_SL g1247 ( 
.A(n_1055),
.B(n_708),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1044),
.B(n_711),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1019),
.B(n_756),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1099),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1079),
.B(n_731),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1072),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1049),
.B(n_765),
.Y(n_1253)
);

INVxp67_ASAP7_75t_L g1254 ( 
.A(n_1046),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1050),
.Y(n_1255)
);

OR2x6_ASAP7_75t_L g1256 ( 
.A(n_1169),
.B(n_685),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1045),
.B(n_1136),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1142),
.B(n_1143),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1152),
.B(n_779),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1152),
.B(n_792),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1015),
.B(n_741),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1159),
.B(n_1160),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1101),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1015),
.B(n_748),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1088),
.B(n_755),
.Y(n_1265)
);

AO221x1_ASAP7_75t_L g1266 ( 
.A1(n_1186),
.A2(n_682),
.B1(n_738),
.B2(n_734),
.C(n_726),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1159),
.B(n_1105),
.Y(n_1267)
);

BUFx5_ASAP7_75t_L g1268 ( 
.A(n_1165),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1016),
.B(n_769),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1014),
.B(n_821),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1016),
.B(n_778),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1025),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1014),
.B(n_865),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1024),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1106),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1102),
.B(n_808),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1024),
.Y(n_1277)
);

INVx8_ASAP7_75t_L g1278 ( 
.A(n_1024),
.Y(n_1278)
);

AO221x1_ASAP7_75t_L g1279 ( 
.A1(n_1169),
.A2(n_738),
.B1(n_826),
.B2(n_763),
.C(n_751),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1059),
.A2(n_559),
.B1(n_568),
.B2(n_560),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1107),
.Y(n_1281)
);

OAI221xp5_ASAP7_75t_L g1282 ( 
.A1(n_1114),
.A2(n_699),
.B1(n_715),
.B2(n_680),
.C(n_667),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1059),
.A2(n_763),
.B1(n_826),
.B2(n_751),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1109),
.Y(n_1284)
);

AOI221xp5_ASAP7_75t_L g1285 ( 
.A1(n_1102),
.A2(n_1148),
.B1(n_1112),
.B2(n_1119),
.C(n_1115),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1071),
.B(n_572),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1111),
.Y(n_1287)
);

NAND3xp33_ASAP7_75t_L g1288 ( 
.A(n_1017),
.B(n_612),
.C(n_609),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1095),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1095),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1089),
.B(n_616),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1089),
.B(n_617),
.Y(n_1292)
);

O2A1O1Ixp5_ASAP7_75t_L g1293 ( 
.A1(n_1163),
.A2(n_709),
.B(n_583),
.C(n_651),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1171),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1032),
.B(n_746),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1093),
.B(n_619),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1093),
.B(n_835),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1094),
.B(n_620),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1068),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1171),
.Y(n_1300)
);

INVx1_ASAP7_75t_SL g1301 ( 
.A(n_1023),
.Y(n_1301)
);

NOR3xp33_ASAP7_75t_L g1302 ( 
.A(n_1117),
.B(n_795),
.C(n_727),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1185),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1029),
.B(n_624),
.Y(n_1304)
);

INVxp33_ASAP7_75t_L g1305 ( 
.A(n_1060),
.Y(n_1305)
);

NAND2x1_ASAP7_75t_L g1306 ( 
.A(n_1013),
.B(n_890),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1041),
.B(n_626),
.Y(n_1307)
);

INVx8_ASAP7_75t_L g1308 ( 
.A(n_1146),
.Y(n_1308)
);

AND3x4_ASAP7_75t_L g1309 ( 
.A(n_1117),
.B(n_845),
.C(n_812),
.Y(n_1309)
);

OR2x6_ASAP7_75t_L g1310 ( 
.A(n_1100),
.B(n_896),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1053),
.B(n_631),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1021),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1054),
.B(n_640),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1020),
.B(n_1027),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1020),
.B(n_647),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1027),
.B(n_648),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1032),
.B(n_654),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1043),
.B(n_555),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1184),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1043),
.B(n_658),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1185),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1030),
.B(n_555),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1131),
.B(n_855),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1028),
.B(n_584),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1028),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1035),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1064),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1064),
.Y(n_1328)
);

INVxp67_ASAP7_75t_L g1329 ( 
.A(n_1038),
.Y(n_1329)
);

NOR3xp33_ASAP7_75t_L g1330 ( 
.A(n_1164),
.B(n_663),
.C(n_659),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1017),
.B(n_656),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1038),
.B(n_664),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1070),
.B(n_665),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1097),
.B(n_668),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1037),
.Y(n_1335)
);

BUFx8_ASAP7_75t_L g1336 ( 
.A(n_1138),
.Y(n_1336)
);

A2O1A1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1092),
.A2(n_649),
.B(n_653),
.C(n_646),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1037),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1097),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1047),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_SL g1341 ( 
.A(n_1167),
.B(n_880),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1110),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1047),
.Y(n_1343)
);

INVx2_ASAP7_75t_SL g1344 ( 
.A(n_1022),
.Y(n_1344)
);

NAND3xp33_ASAP7_75t_L g1345 ( 
.A(n_1135),
.B(n_673),
.C(n_670),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1048),
.B(n_712),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1048),
.Y(n_1347)
);

INVxp67_ASAP7_75t_L g1348 ( 
.A(n_1040),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1040),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1135),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1057),
.B(n_719),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1058),
.B(n_555),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1058),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1066),
.Y(n_1354)
);

NOR2xp67_ASAP7_75t_L g1355 ( 
.A(n_1080),
.B(n_30),
.Y(n_1355)
);

O2A1O1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1156),
.A2(n_655),
.B(n_661),
.C(n_660),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1151),
.B(n_719),
.Y(n_1357)
);

OR2x6_ASAP7_75t_L g1358 ( 
.A(n_1156),
.B(n_740),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1184),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1138),
.B(n_686),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_SL g1361 ( 
.A(n_1184),
.B(n_564),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1164),
.B(n_690),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1180),
.B(n_564),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1172),
.Y(n_1364)
);

NAND2xp33_ASAP7_75t_L g1365 ( 
.A(n_1012),
.B(n_564),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1174),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1174),
.B(n_740),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1168),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1173),
.B(n_749),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1080),
.B(n_693),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1170),
.A2(n_666),
.B1(n_671),
.B2(n_662),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1177),
.B(n_749),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1178),
.B(n_777),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1090),
.B(n_695),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1181),
.B(n_777),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1012),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1069),
.Y(n_1377)
);

BUFx5_ASAP7_75t_L g1378 ( 
.A(n_1170),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1090),
.B(n_701),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1012),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1074),
.B(n_783),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1074),
.B(n_702),
.Y(n_1382)
);

INVx8_ASAP7_75t_L g1383 ( 
.A(n_1012),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1076),
.A2(n_677),
.B1(n_679),
.B2(n_674),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1067),
.B(n_753),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1183),
.B(n_704),
.Y(n_1386)
);

NAND2xp33_ASAP7_75t_L g1387 ( 
.A(n_1067),
.B(n_753),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1083),
.B(n_783),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1084),
.A2(n_880),
.B1(n_901),
.B2(n_836),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1067),
.B(n_753),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1084),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1067),
.B(n_705),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1091),
.B(n_793),
.Y(n_1393)
);

OR2x6_ASAP7_75t_L g1394 ( 
.A(n_1096),
.B(n_804),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1147),
.Y(n_1395)
);

INVx8_ASAP7_75t_L g1396 ( 
.A(n_1147),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1103),
.B(n_706),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1104),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1108),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1108),
.B(n_877),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1113),
.Y(n_1401)
);

AND2x4_ASAP7_75t_SL g1402 ( 
.A(n_1155),
.B(n_836),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1118),
.B(n_713),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1118),
.B(n_877),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1123),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1129),
.Y(n_1406)
);

NAND2xp33_ASAP7_75t_L g1407 ( 
.A(n_1130),
.B(n_754),
.Y(n_1407)
);

INVx8_ASAP7_75t_L g1408 ( 
.A(n_1133),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1137),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1137),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1139),
.B(n_718),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1207),
.B(n_720),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1190),
.B(n_901),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1214),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1216),
.B(n_1192),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1278),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1191),
.B(n_721),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1191),
.B(n_722),
.Y(n_1418)
);

AO21x1_ASAP7_75t_L g1419 ( 
.A1(n_1270),
.A2(n_684),
.B(n_681),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1289),
.A2(n_691),
.B1(n_697),
.B2(n_687),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1278),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1278),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1218),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1212),
.B(n_723),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1220),
.Y(n_1425)
);

AOI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1357),
.A2(n_1162),
.B(n_1161),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1205),
.B(n_724),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_R g1428 ( 
.A(n_1208),
.B(n_725),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1215),
.B(n_728),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1205),
.B(n_1258),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1233),
.A2(n_1314),
.B(n_1262),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1268),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1262),
.A2(n_1175),
.B(n_1166),
.Y(n_1433)
);

NOR2x1_ASAP7_75t_L g1434 ( 
.A(n_1246),
.B(n_707),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1301),
.B(n_739),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1257),
.B(n_742),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1268),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1217),
.B(n_745),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1227),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1301),
.B(n_752),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1198),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1188),
.B(n_757),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1217),
.B(n_759),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1270),
.A2(n_1175),
.B(n_1166),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1273),
.A2(n_1179),
.B(n_1176),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1273),
.A2(n_1179),
.B(n_1176),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1357),
.A2(n_714),
.B(n_710),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1227),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1293),
.A2(n_717),
.B(n_716),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1194),
.B(n_760),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1195),
.B(n_762),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1201),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1189),
.B(n_764),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1268),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_SL g1455 ( 
.A(n_1210),
.B(n_772),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1402),
.Y(n_1456)
);

BUFx12f_ASAP7_75t_L g1457 ( 
.A(n_1336),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1268),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1267),
.B(n_1203),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1268),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1389),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1236),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1319),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1210),
.B(n_766),
.Y(n_1464)
);

NOR3xp33_ASAP7_75t_L g1465 ( 
.A(n_1204),
.B(n_770),
.C(n_768),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1342),
.A2(n_1182),
.B(n_737),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1243),
.A2(n_781),
.B1(n_782),
.B2(n_773),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1285),
.B(n_784),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1252),
.B(n_736),
.Y(n_1469)
);

A2O1A1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1290),
.A2(n_744),
.B(n_747),
.C(n_743),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1232),
.B(n_788),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1226),
.B(n_791),
.Y(n_1472)
);

A2O1A1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1245),
.A2(n_761),
.B(n_767),
.C(n_750),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1350),
.A2(n_774),
.B(n_771),
.Y(n_1474)
);

AOI33xp33_ASAP7_75t_L g1475 ( 
.A1(n_1244),
.A2(n_796),
.A3(n_776),
.B1(n_797),
.B2(n_790),
.B3(n_775),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1230),
.B(n_1254),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1228),
.B(n_1263),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1329),
.B(n_798),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1337),
.A2(n_803),
.B(n_799),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1255),
.B(n_806),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1275),
.B(n_794),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1200),
.A2(n_810),
.B(n_807),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1256),
.A2(n_815),
.B1(n_822),
.B2(n_818),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1209),
.A2(n_829),
.B(n_823),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1202),
.B(n_801),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1281),
.B(n_802),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1237),
.B(n_811),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1242),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1211),
.A2(n_834),
.B(n_832),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1231),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1250),
.B(n_819),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1319),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1331),
.A2(n_846),
.B(n_839),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1284),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1280),
.B(n_820),
.Y(n_1495)
);

INVx4_ASAP7_75t_L g1496 ( 
.A(n_1308),
.Y(n_1496)
);

O2A1O1Ixp5_ASAP7_75t_L g1497 ( 
.A1(n_1318),
.A2(n_891),
.B(n_857),
.C(n_859),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1287),
.B(n_824),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1229),
.Y(n_1499)
);

O2A1O1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1234),
.A2(n_864),
.B(n_866),
.C(n_851),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1295),
.B(n_867),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1324),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1327),
.A2(n_870),
.B(n_868),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1331),
.A2(n_878),
.B(n_872),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1256),
.A2(n_882),
.B1(n_883),
.B2(n_881),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1224),
.B(n_825),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1328),
.A2(n_894),
.B(n_887),
.Y(n_1507)
);

CKINVDCx6p67_ASAP7_75t_R g1508 ( 
.A(n_1349),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1202),
.B(n_827),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1324),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_SL g1511 ( 
.A1(n_1266),
.A2(n_830),
.B1(n_833),
.B2(n_831),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1274),
.B(n_1277),
.Y(n_1512)
);

O2A1O1Ixp5_ASAP7_75t_L g1513 ( 
.A1(n_1297),
.A2(n_850),
.B(n_875),
.C(n_800),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1288),
.B(n_837),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1199),
.Y(n_1515)
);

O2A1O1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1282),
.A2(n_840),
.B(n_842),
.C(n_841),
.Y(n_1516)
);

NOR3xp33_ASAP7_75t_L g1517 ( 
.A(n_1204),
.B(n_1283),
.C(n_1389),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1346),
.Y(n_1518)
);

AND2x2_ASAP7_75t_SL g1519 ( 
.A(n_1341),
.B(n_800),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1219),
.B(n_844),
.Y(n_1520)
);

BUFx8_ASAP7_75t_L g1521 ( 
.A(n_1344),
.Y(n_1521)
);

O2A1O1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1213),
.A2(n_848),
.B(n_854),
.C(n_853),
.Y(n_1522)
);

INVxp67_ASAP7_75t_L g1523 ( 
.A(n_1341),
.Y(n_1523)
);

O2A1O1Ixp33_ASAP7_75t_L g1524 ( 
.A1(n_1356),
.A2(n_858),
.B(n_861),
.C(n_856),
.Y(n_1524)
);

INVxp67_ASAP7_75t_L g1525 ( 
.A(n_1298),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1222),
.B(n_862),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1265),
.B(n_863),
.Y(n_1527)
);

OAI21xp33_ASAP7_75t_L g1528 ( 
.A1(n_1286),
.A2(n_1292),
.B(n_1291),
.Y(n_1528)
);

CKINVDCx10_ASAP7_75t_R g1529 ( 
.A(n_1310),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1346),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1351),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1187),
.Y(n_1532)
);

OAI21xp33_ASAP7_75t_L g1533 ( 
.A1(n_1296),
.A2(n_871),
.B(n_850),
.Y(n_1533)
);

NOR2x1_ASAP7_75t_L g1534 ( 
.A(n_1323),
.B(n_800),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1382),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1304),
.A2(n_1311),
.B(n_1307),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1283),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1256),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1235),
.B(n_28),
.Y(n_1539)
);

O2A1O1Ixp33_ASAP7_75t_L g1540 ( 
.A1(n_1259),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_1540)
);

NAND2x1p5_ASAP7_75t_L g1541 ( 
.A(n_1199),
.B(n_32),
.Y(n_1541)
);

AO21x1_ASAP7_75t_L g1542 ( 
.A1(n_1295),
.A2(n_33),
.B(n_34),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1358),
.B(n_33),
.Y(n_1543)
);

OAI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1294),
.A2(n_1303),
.B(n_1300),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1260),
.B(n_34),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1260),
.B(n_37),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1386),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1397),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1308),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1308),
.B(n_38),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1367),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1358),
.B(n_38),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1359),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1317),
.B(n_39),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1367),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1320),
.B(n_41),
.Y(n_1556)
);

INVx2_ASAP7_75t_SL g1557 ( 
.A(n_1221),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1253),
.B(n_41),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1358),
.B(n_42),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1253),
.B(n_1249),
.Y(n_1560)
);

OR2x6_ASAP7_75t_L g1561 ( 
.A(n_1272),
.B(n_43),
.Y(n_1561)
);

AO21x1_ASAP7_75t_L g1562 ( 
.A1(n_1381),
.A2(n_43),
.B(n_45),
.Y(n_1562)
);

AOI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1276),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1563)
);

A2O1A1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1321),
.A2(n_49),
.B(n_46),
.C(n_48),
.Y(n_1564)
);

O2A1O1Ixp33_ASAP7_75t_L g1565 ( 
.A1(n_1261),
.A2(n_51),
.B(n_48),
.C(n_50),
.Y(n_1565)
);

AND2x6_ASAP7_75t_L g1566 ( 
.A(n_1339),
.B(n_472),
.Y(n_1566)
);

OAI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1343),
.A2(n_474),
.B(n_473),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1221),
.B(n_1223),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1334),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1384),
.A2(n_55),
.B1(n_52),
.B2(n_54),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1225),
.B(n_1313),
.Y(n_1571)
);

A2O1A1Ixp33_ASAP7_75t_L g1572 ( 
.A1(n_1347),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_1572)
);

O2A1O1Ixp33_ASAP7_75t_SL g1573 ( 
.A1(n_1306),
.A2(n_1363),
.B(n_1197),
.C(n_1206),
.Y(n_1573)
);

BUFx2_ASAP7_75t_SL g1574 ( 
.A(n_1241),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1360),
.B(n_57),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1264),
.B(n_58),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1269),
.B(n_1271),
.Y(n_1577)
);

CKINVDCx8_ASAP7_75t_R g1578 ( 
.A(n_1310),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1279),
.B(n_59),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1240),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1394),
.A2(n_65),
.B1(n_62),
.B2(n_64),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1193),
.Y(n_1582)
);

AOI33xp33_ASAP7_75t_L g1583 ( 
.A1(n_1332),
.A2(n_65),
.A3(n_68),
.B1(n_62),
.B2(n_64),
.B3(n_67),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1315),
.B(n_69),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1248),
.B(n_1238),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1316),
.B(n_1353),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1196),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1383),
.Y(n_1588)
);

NOR2x1_ASAP7_75t_L g1589 ( 
.A(n_1310),
.B(n_1309),
.Y(n_1589)
);

AND2x4_ASAP7_75t_SL g1590 ( 
.A(n_1302),
.B(n_71),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1394),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_1383),
.Y(n_1592)
);

A2O1A1Ixp33_ASAP7_75t_L g1593 ( 
.A1(n_1369),
.A2(n_76),
.B(n_74),
.C(n_75),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1333),
.B(n_75),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1362),
.B(n_78),
.Y(n_1595)
);

BUFx12f_ASAP7_75t_L g1596 ( 
.A(n_1336),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1305),
.B(n_78),
.Y(n_1597)
);

OAI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1312),
.A2(n_485),
.B(n_484),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1370),
.B(n_80),
.Y(n_1599)
);

INVx4_ASAP7_75t_L g1600 ( 
.A(n_1383),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1345),
.B(n_81),
.Y(n_1601)
);

A2O1A1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1369),
.A2(n_86),
.B(n_83),
.C(n_85),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1394),
.A2(n_88),
.B1(n_85),
.B2(n_87),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1251),
.B(n_87),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1374),
.B(n_1379),
.Y(n_1605)
);

A2O1A1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1372),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1299),
.B(n_91),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1326),
.B(n_92),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1372),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1373),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1325),
.A2(n_495),
.B(n_494),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1392),
.B(n_94),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1239),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_1613)
);

INVx2_ASAP7_75t_SL g1614 ( 
.A(n_1247),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1348),
.B(n_95),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1335),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1338),
.B(n_98),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1340),
.A2(n_497),
.B(n_496),
.Y(n_1618)
);

OAI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1354),
.A2(n_501),
.B(n_500),
.Y(n_1619)
);

OAI321xp33_ASAP7_75t_L g1620 ( 
.A1(n_1375),
.A2(n_102),
.A3(n_105),
.B1(n_99),
.B2(n_100),
.C(n_103),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_SL g1621 ( 
.A1(n_1330),
.A2(n_103),
.B1(n_99),
.B2(n_100),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1403),
.B(n_1411),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1371),
.B(n_107),
.Y(n_1623)
);

NOR2x1p5_ASAP7_75t_L g1624 ( 
.A(n_1355),
.B(n_1388),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1364),
.A2(n_503),
.B(n_502),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1388),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1393),
.Y(n_1627)
);

O2A1O1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1393),
.A2(n_110),
.B(n_108),
.C(n_109),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1408),
.B(n_111),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1408),
.B(n_112),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1322),
.A2(n_506),
.B(n_505),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_R g1632 ( 
.A(n_1396),
.B(n_112),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1361),
.B(n_113),
.Y(n_1633)
);

AOI21xp33_ASAP7_75t_L g1634 ( 
.A1(n_1408),
.A2(n_113),
.B(n_114),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1400),
.B(n_115),
.Y(n_1635)
);

OR2x6_ASAP7_75t_L g1636 ( 
.A(n_1396),
.B(n_1404),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1366),
.B(n_117),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1352),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1380),
.B(n_121),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1396),
.B(n_121),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1391),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_1641)
);

AOI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1406),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1378),
.Y(n_1643)
);

BUFx6f_ASAP7_75t_L g1644 ( 
.A(n_1376),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1368),
.A2(n_129),
.B1(n_126),
.B2(n_128),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1409),
.B(n_126),
.Y(n_1646)
);

BUFx12f_ASAP7_75t_L g1647 ( 
.A(n_1376),
.Y(n_1647)
);

BUFx2_ASAP7_75t_SL g1648 ( 
.A(n_1385),
.Y(n_1648)
);

BUFx4f_ASAP7_75t_L g1649 ( 
.A(n_1395),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1395),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1377),
.B(n_130),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1395),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1398),
.B(n_131),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1399),
.B(n_131),
.Y(n_1654)
);

OR2x6_ASAP7_75t_L g1655 ( 
.A(n_1390),
.B(n_132),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1401),
.A2(n_1410),
.B(n_1405),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1407),
.B(n_133),
.Y(n_1657)
);

NOR3xp33_ASAP7_75t_L g1658 ( 
.A(n_1365),
.B(n_133),
.C(n_134),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1387),
.B(n_134),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1207),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1207),
.B(n_137),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1207),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1190),
.B(n_138),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_SL g1664 ( 
.A1(n_1305),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1207),
.B(n_139),
.Y(n_1665)
);

INVx3_ASAP7_75t_L g1666 ( 
.A(n_1421),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1430),
.B(n_141),
.Y(n_1667)
);

BUFx6f_ASAP7_75t_L g1668 ( 
.A(n_1644),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1519),
.B(n_530),
.Y(n_1669)
);

A2O1A1Ixp33_ASAP7_75t_L g1670 ( 
.A1(n_1536),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_1670)
);

INVx5_ASAP7_75t_L g1671 ( 
.A(n_1421),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1415),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1421),
.B(n_142),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1422),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1560),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_1675)
);

AOI221x1_ASAP7_75t_L g1676 ( 
.A1(n_1449),
.A2(n_149),
.B1(n_145),
.B2(n_148),
.C(n_150),
.Y(n_1676)
);

OAI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1477),
.A2(n_533),
.B(n_532),
.Y(n_1677)
);

INVx3_ASAP7_75t_L g1678 ( 
.A(n_1600),
.Y(n_1678)
);

AOI21xp33_ASAP7_75t_L g1679 ( 
.A1(n_1605),
.A2(n_148),
.B(n_149),
.Y(n_1679)
);

NOR2x1_ASAP7_75t_L g1680 ( 
.A(n_1496),
.B(n_151),
.Y(n_1680)
);

INVx2_ASAP7_75t_SL g1681 ( 
.A(n_1422),
.Y(n_1681)
);

A2O1A1Ixp33_ASAP7_75t_L g1682 ( 
.A1(n_1583),
.A2(n_155),
.B(n_153),
.C(n_154),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1413),
.A2(n_156),
.B1(n_153),
.B2(n_154),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1535),
.B(n_1414),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1535),
.B(n_156),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_SL g1686 ( 
.A1(n_1544),
.A2(n_157),
.B(n_158),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1412),
.B(n_157),
.Y(n_1687)
);

OAI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1544),
.A2(n_540),
.B(n_539),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1537),
.B(n_158),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1547),
.B(n_159),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1441),
.Y(n_1691)
);

A2O1A1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1528),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1517),
.B(n_164),
.Y(n_1693)
);

NAND2x1_ASAP7_75t_L g1694 ( 
.A(n_1600),
.B(n_1416),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1627),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1540),
.A2(n_169),
.B(n_166),
.C(n_168),
.Y(n_1696)
);

NOR2x1_ASAP7_75t_SL g1697 ( 
.A(n_1496),
.B(n_168),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1502),
.A2(n_1510),
.B(n_1518),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1429),
.B(n_172),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1476),
.B(n_1465),
.Y(n_1700)
);

AO31x2_ASAP7_75t_L g1701 ( 
.A1(n_1562),
.A2(n_175),
.A3(n_173),
.B(n_174),
.Y(n_1701)
);

AND3x2_ASAP7_75t_L g1702 ( 
.A(n_1523),
.B(n_176),
.C(n_177),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1586),
.A2(n_178),
.B(n_179),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1656),
.A2(n_180),
.B(n_181),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1644),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1530),
.A2(n_182),
.B(n_180),
.C(n_181),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1622),
.A2(n_185),
.B(n_186),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1461),
.B(n_187),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1459),
.A2(n_188),
.B(n_189),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1525),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1571),
.A2(n_191),
.B(n_192),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1485),
.B(n_193),
.Y(n_1712)
);

A2O1A1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1531),
.A2(n_195),
.B(n_193),
.C(n_194),
.Y(n_1713)
);

AO21x1_ASAP7_75t_L g1714 ( 
.A1(n_1567),
.A2(n_194),
.B(n_196),
.Y(n_1714)
);

OAI21x1_ASAP7_75t_L g1715 ( 
.A1(n_1598),
.A2(n_196),
.B(n_197),
.Y(n_1715)
);

OAI21x1_ASAP7_75t_L g1716 ( 
.A1(n_1598),
.A2(n_199),
.B(n_200),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1444),
.A2(n_200),
.B(n_201),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1568),
.B(n_202),
.Y(n_1718)
);

AOI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1445),
.A2(n_1446),
.B(n_1433),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1494),
.Y(n_1720)
);

OAI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1447),
.A2(n_204),
.B(n_205),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1432),
.Y(n_1722)
);

NAND3x1_ASAP7_75t_L g1723 ( 
.A(n_1589),
.B(n_206),
.C(n_207),
.Y(n_1723)
);

OAI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1447),
.A2(n_206),
.B(n_209),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1437),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1609),
.A2(n_213),
.B1(n_210),
.B2(n_212),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1452),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1509),
.B(n_212),
.Y(n_1728)
);

OAI21x1_ASAP7_75t_L g1729 ( 
.A1(n_1611),
.A2(n_215),
.B(n_216),
.Y(n_1729)
);

O2A1O1Ixp5_ASAP7_75t_L g1730 ( 
.A1(n_1419),
.A2(n_218),
.B(n_216),
.C(n_217),
.Y(n_1730)
);

AOI221x1_ASAP7_75t_L g1731 ( 
.A1(n_1581),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.C(n_223),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1521),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1547),
.B(n_1539),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1499),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1548),
.B(n_224),
.Y(n_1735)
);

OAI21x1_ASAP7_75t_L g1736 ( 
.A1(n_1611),
.A2(n_226),
.B(n_227),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1471),
.B(n_228),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1643),
.A2(n_229),
.B(n_230),
.Y(n_1738)
);

AO31x2_ASAP7_75t_L g1739 ( 
.A1(n_1542),
.A2(n_234),
.A3(n_230),
.B(n_231),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1610),
.A2(n_235),
.B(n_236),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1454),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1475),
.B(n_1575),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1458),
.Y(n_1743)
);

BUFx8_ASAP7_75t_SL g1744 ( 
.A(n_1457),
.Y(n_1744)
);

OAI21x1_ASAP7_75t_SL g1745 ( 
.A1(n_1618),
.A2(n_239),
.B(n_240),
.Y(n_1745)
);

CKINVDCx20_ASAP7_75t_R g1746 ( 
.A(n_1439),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1551),
.B(n_241),
.Y(n_1747)
);

OAI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1555),
.A2(n_244),
.B(n_245),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1417),
.B(n_244),
.Y(n_1749)
);

BUFx6f_ASAP7_75t_L g1750 ( 
.A(n_1647),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1460),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1469),
.B(n_246),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1418),
.B(n_246),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1427),
.A2(n_247),
.B(n_248),
.Y(n_1754)
);

INVxp67_ASAP7_75t_L g1755 ( 
.A(n_1469),
.Y(n_1755)
);

NAND2x1p5_ASAP7_75t_L g1756 ( 
.A(n_1416),
.B(n_249),
.Y(n_1756)
);

AND2x2_ASAP7_75t_SL g1757 ( 
.A(n_1538),
.B(n_250),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1661),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1456),
.B(n_252),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1490),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1438),
.B(n_253),
.Y(n_1761)
);

AND2x2_ASAP7_75t_SL g1762 ( 
.A(n_1649),
.B(n_254),
.Y(n_1762)
);

NOR2xp67_ASAP7_75t_L g1763 ( 
.A(n_1596),
.B(n_254),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1443),
.B(n_1468),
.Y(n_1764)
);

OAI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1474),
.A2(n_255),
.B(n_256),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1636),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1470),
.B(n_261),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1588),
.Y(n_1768)
);

OAI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1503),
.A2(n_264),
.B(n_266),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1424),
.A2(n_1663),
.B1(n_1495),
.B2(n_1595),
.Y(n_1770)
);

CKINVDCx20_ASAP7_75t_R g1771 ( 
.A(n_1448),
.Y(n_1771)
);

OAI21x1_ASAP7_75t_L g1772 ( 
.A1(n_1618),
.A2(n_267),
.B(n_268),
.Y(n_1772)
);

OAI21xp33_ASAP7_75t_L g1773 ( 
.A1(n_1436),
.A2(n_268),
.B(n_270),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1423),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1425),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1442),
.A2(n_270),
.B(n_271),
.Y(n_1776)
);

OAI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1507),
.A2(n_273),
.B(n_274),
.Y(n_1777)
);

AO21x1_ASAP7_75t_L g1778 ( 
.A1(n_1619),
.A2(n_273),
.B(n_275),
.Y(n_1778)
);

OAI21x1_ASAP7_75t_L g1779 ( 
.A1(n_1619),
.A2(n_275),
.B(n_276),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1481),
.A2(n_278),
.B(n_279),
.Y(n_1780)
);

AO21x1_ASAP7_75t_L g1781 ( 
.A1(n_1541),
.A2(n_280),
.B(n_281),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1480),
.B(n_282),
.Y(n_1782)
);

OAI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1482),
.A2(n_283),
.B(n_284),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_SL g1784 ( 
.A1(n_1636),
.A2(n_285),
.B(n_286),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1549),
.B(n_287),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1636),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_1786)
);

INVxp67_ASAP7_75t_L g1787 ( 
.A(n_1616),
.Y(n_1787)
);

AOI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1486),
.A2(n_292),
.B(n_293),
.Y(n_1788)
);

OAI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1484),
.A2(n_292),
.B(n_294),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1480),
.B(n_294),
.Y(n_1790)
);

NAND2x1p5_ASAP7_75t_L g1791 ( 
.A(n_1588),
.B(n_295),
.Y(n_1791)
);

OAI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1489),
.A2(n_296),
.B(n_298),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1483),
.B(n_299),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1472),
.A2(n_301),
.B(n_302),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1473),
.B(n_301),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_SL g1796 ( 
.A(n_1578),
.B(n_302),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1501),
.B(n_303),
.Y(n_1797)
);

AOI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1520),
.A2(n_304),
.B(n_305),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1466),
.A2(n_304),
.B(n_308),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1488),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1462),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1582),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1434),
.B(n_310),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1561),
.B(n_312),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1549),
.B(n_313),
.Y(n_1805)
);

AOI221x1_ASAP7_75t_L g1806 ( 
.A1(n_1581),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.C(n_317),
.Y(n_1806)
);

OAI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1493),
.A2(n_315),
.B(n_316),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1587),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1526),
.A2(n_318),
.B(n_320),
.Y(n_1809)
);

OAI21x1_ASAP7_75t_SL g1810 ( 
.A1(n_1660),
.A2(n_325),
.B(n_326),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1592),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1558),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1532),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1435),
.B(n_326),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1428),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1501),
.B(n_327),
.Y(n_1816)
);

CKINVDCx8_ASAP7_75t_R g1817 ( 
.A(n_1529),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1561),
.B(n_1543),
.Y(n_1818)
);

BUFx12f_ASAP7_75t_L g1819 ( 
.A(n_1521),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1493),
.B(n_328),
.Y(n_1820)
);

OAI21x1_ASAP7_75t_L g1821 ( 
.A1(n_1625),
.A2(n_329),
.B(n_330),
.Y(n_1821)
);

OAI22x1_ASAP7_75t_L g1822 ( 
.A1(n_1541),
.A2(n_329),
.B1(n_330),
.B2(n_331),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1545),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1546),
.A2(n_1660),
.B1(n_1591),
.B2(n_1603),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1579),
.A2(n_331),
.B1(n_332),
.B2(n_333),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1506),
.A2(n_1577),
.B(n_1451),
.Y(n_1826)
);

INVx4_ASAP7_75t_L g1827 ( 
.A(n_1592),
.Y(n_1827)
);

INVxp67_ASAP7_75t_L g1828 ( 
.A(n_1455),
.Y(n_1828)
);

AOI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1450),
.A2(n_334),
.B(n_335),
.Y(n_1829)
);

AOI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1453),
.A2(n_336),
.B(n_337),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1665),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1504),
.B(n_336),
.Y(n_1832)
);

INVx1_ASAP7_75t_SL g1833 ( 
.A(n_1632),
.Y(n_1833)
);

A2O1A1Ixp33_ASAP7_75t_L g1834 ( 
.A1(n_1628),
.A2(n_338),
.B(n_339),
.C(n_340),
.Y(n_1834)
);

OR2x4_ASAP7_75t_L g1835 ( 
.A(n_1594),
.B(n_339),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1504),
.B(n_341),
.Y(n_1836)
);

NAND2x1p5_ASAP7_75t_L g1837 ( 
.A(n_1592),
.B(n_341),
.Y(n_1837)
);

OAI21x1_ASAP7_75t_SL g1838 ( 
.A1(n_1591),
.A2(n_343),
.B(n_344),
.Y(n_1838)
);

OA22x2_ASAP7_75t_L g1839 ( 
.A1(n_1561),
.A2(n_1505),
.B1(n_1664),
.B2(n_1590),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1552),
.B(n_344),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1553),
.B(n_345),
.Y(n_1841)
);

OAI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1584),
.A2(n_346),
.B(n_347),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1607),
.A2(n_346),
.B(n_348),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1500),
.B(n_1479),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1440),
.B(n_1527),
.Y(n_1845)
);

INVx2_ASAP7_75t_SL g1846 ( 
.A(n_1508),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1557),
.B(n_1467),
.Y(n_1847)
);

BUFx2_ASAP7_75t_SL g1848 ( 
.A(n_1566),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1479),
.B(n_348),
.Y(n_1849)
);

BUFx3_ASAP7_75t_L g1850 ( 
.A(n_1463),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1559),
.B(n_349),
.Y(n_1851)
);

O2A1O1Ixp5_ASAP7_75t_L g1852 ( 
.A1(n_1612),
.A2(n_350),
.B(n_351),
.C(n_352),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1585),
.B(n_355),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1585),
.B(n_1487),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1455),
.B(n_355),
.Y(n_1855)
);

OAI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1603),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1491),
.Y(n_1857)
);

A2O1A1Ixp33_ASAP7_75t_L g1858 ( 
.A1(n_1565),
.A2(n_360),
.B(n_361),
.C(n_362),
.Y(n_1858)
);

OAI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1608),
.A2(n_361),
.B(n_363),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1498),
.A2(n_363),
.B(n_364),
.Y(n_1860)
);

OAI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1617),
.A2(n_365),
.B(n_366),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1505),
.A2(n_365),
.B1(n_367),
.B2(n_368),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1597),
.B(n_367),
.Y(n_1863)
);

INVx1_ASAP7_75t_SL g1864 ( 
.A(n_1615),
.Y(n_1864)
);

OR2x6_ASAP7_75t_L g1865 ( 
.A(n_1574),
.B(n_1550),
.Y(n_1865)
);

AOI21xp5_ASAP7_75t_L g1866 ( 
.A1(n_1604),
.A2(n_369),
.B(n_371),
.Y(n_1866)
);

AOI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1650),
.A2(n_373),
.B(n_374),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1420),
.B(n_1478),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1652),
.A2(n_373),
.B(n_374),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1573),
.A2(n_375),
.B(n_377),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1641),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1524),
.B(n_378),
.Y(n_1872)
);

AND3x4_ASAP7_75t_L g1873 ( 
.A(n_1534),
.B(n_379),
.C(n_380),
.Y(n_1873)
);

AOI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1514),
.A2(n_379),
.B(n_381),
.Y(n_1874)
);

AOI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1533),
.A2(n_383),
.B(n_384),
.Y(n_1875)
);

AO21x2_ASAP7_75t_L g1876 ( 
.A1(n_1651),
.A2(n_384),
.B(n_387),
.Y(n_1876)
);

AOI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1554),
.A2(n_388),
.B(n_389),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1420),
.B(n_388),
.Y(n_1878)
);

OAI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1635),
.A2(n_389),
.B(n_390),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1614),
.B(n_393),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1626),
.A2(n_394),
.B1(n_395),
.B2(n_397),
.Y(n_1881)
);

NAND2xp33_ASAP7_75t_L g1882 ( 
.A(n_1566),
.B(n_395),
.Y(n_1882)
);

OAI21xp5_ASAP7_75t_L g1883 ( 
.A1(n_1497),
.A2(n_398),
.B(n_399),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1522),
.B(n_398),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1511),
.B(n_1621),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1512),
.B(n_399),
.Y(n_1886)
);

OA21x2_ASAP7_75t_L g1887 ( 
.A1(n_1620),
.A2(n_403),
.B(n_404),
.Y(n_1887)
);

INVxp67_ASAP7_75t_SL g1888 ( 
.A(n_1646),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1516),
.B(n_404),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1599),
.B(n_405),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1645),
.Y(n_1891)
);

NAND2x1p5_ASAP7_75t_L g1892 ( 
.A(n_1463),
.B(n_405),
.Y(n_1892)
);

OAI21x1_ASAP7_75t_L g1893 ( 
.A1(n_1631),
.A2(n_406),
.B(n_407),
.Y(n_1893)
);

OAI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1654),
.A2(n_1637),
.B(n_1576),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1638),
.A2(n_406),
.B(n_409),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1556),
.A2(n_409),
.B(n_411),
.Y(n_1896)
);

AO31x2_ASAP7_75t_L g1897 ( 
.A1(n_1564),
.A2(n_1602),
.A3(n_1593),
.B(n_1606),
.Y(n_1897)
);

OAI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1653),
.A2(n_411),
.B(n_412),
.Y(n_1898)
);

OAI21xp33_ASAP7_75t_SL g1899 ( 
.A1(n_1563),
.A2(n_1624),
.B(n_1569),
.Y(n_1899)
);

INVx5_ASAP7_75t_L g1900 ( 
.A(n_1566),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1645),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1492),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1570),
.B(n_413),
.Y(n_1903)
);

OAI21x1_ASAP7_75t_SL g1904 ( 
.A1(n_1640),
.A2(n_415),
.B(n_416),
.Y(n_1904)
);

OAI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1629),
.A2(n_1630),
.B1(n_1642),
.B2(n_1492),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1580),
.B(n_415),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1613),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1464),
.B(n_417),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1515),
.B(n_417),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1515),
.B(n_418),
.Y(n_1910)
);

BUFx6f_ASAP7_75t_L g1911 ( 
.A(n_1566),
.Y(n_1911)
);

AND2x6_ASAP7_75t_L g1912 ( 
.A(n_1639),
.B(n_418),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1623),
.B(n_419),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1655),
.Y(n_1914)
);

BUFx6f_ASAP7_75t_L g1915 ( 
.A(n_1655),
.Y(n_1915)
);

NAND2x1p5_ASAP7_75t_L g1916 ( 
.A(n_1601),
.B(n_1633),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1572),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1634),
.B(n_424),
.Y(n_1918)
);

OAI21x1_ASAP7_75t_L g1919 ( 
.A1(n_1659),
.A2(n_425),
.B(n_426),
.Y(n_1919)
);

BUFx2_ASAP7_75t_L g1920 ( 
.A(n_1655),
.Y(n_1920)
);

OAI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1658),
.A2(n_425),
.B(n_426),
.Y(n_1921)
);

OA21x2_ASAP7_75t_L g1922 ( 
.A1(n_1657),
.A2(n_428),
.B(n_429),
.Y(n_1922)
);

A2O1A1Ixp33_ASAP7_75t_L g1923 ( 
.A1(n_1648),
.A2(n_429),
.B(n_430),
.C(n_431),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1430),
.A2(n_430),
.B(n_431),
.Y(n_1924)
);

A2O1A1Ixp33_ASAP7_75t_L g1925 ( 
.A1(n_1662),
.A2(n_432),
.B(n_434),
.C(n_436),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1662),
.B(n_437),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1430),
.B(n_437),
.Y(n_1927)
);

AOI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1430),
.A2(n_439),
.B(n_440),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1430),
.A2(n_439),
.B(n_440),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1430),
.A2(n_441),
.B(n_442),
.Y(n_1930)
);

OAI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1662),
.A2(n_443),
.B1(n_444),
.B2(n_445),
.Y(n_1931)
);

AOI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1430),
.A2(n_444),
.B(n_446),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1662),
.B(n_448),
.Y(n_1933)
);

AOI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1430),
.A2(n_449),
.B(n_450),
.Y(n_1934)
);

AO31x2_ASAP7_75t_L g1935 ( 
.A1(n_1562),
.A2(n_449),
.A3(n_450),
.B(n_452),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1430),
.A2(n_452),
.B(n_453),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1662),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1662),
.B(n_454),
.Y(n_1938)
);

AOI21x1_ASAP7_75t_L g1939 ( 
.A1(n_1426),
.A2(n_455),
.B(n_456),
.Y(n_1939)
);

NOR2x1_ASAP7_75t_R g1940 ( 
.A(n_1457),
.B(n_1596),
.Y(n_1940)
);

INVx4_ASAP7_75t_SL g1941 ( 
.A(n_1566),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1662),
.B(n_1207),
.Y(n_1942)
);

BUFx4f_ASAP7_75t_L g1943 ( 
.A(n_1457),
.Y(n_1943)
);

OR2x6_ASAP7_75t_L g1944 ( 
.A(n_1421),
.B(n_1278),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1662),
.B(n_1207),
.Y(n_1945)
);

AOI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1430),
.A2(n_1092),
.B(n_1017),
.Y(n_1946)
);

AOI21xp33_ASAP7_75t_L g1947 ( 
.A1(n_1430),
.A2(n_1605),
.B(n_1662),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1430),
.B(n_1059),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1430),
.A2(n_1092),
.B(n_1017),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1662),
.B(n_1207),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1662),
.B(n_1207),
.Y(n_1951)
);

A2O1A1Ixp33_ASAP7_75t_L g1952 ( 
.A1(n_1662),
.A2(n_1430),
.B(n_1536),
.C(n_1449),
.Y(n_1952)
);

AOI22xp33_ASAP7_75t_L g1953 ( 
.A1(n_1517),
.A2(n_1662),
.B1(n_1539),
.B2(n_1430),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1662),
.B(n_1207),
.Y(n_1954)
);

OAI21xp5_ASAP7_75t_L g1955 ( 
.A1(n_1431),
.A2(n_1430),
.B(n_1536),
.Y(n_1955)
);

O2A1O1Ixp5_ASAP7_75t_L g1956 ( 
.A1(n_1449),
.A2(n_1419),
.B(n_1513),
.C(n_1562),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1519),
.B(n_1662),
.Y(n_1957)
);

INVx3_ASAP7_75t_L g1958 ( 
.A(n_1421),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1662),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1662),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1662),
.B(n_1192),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1662),
.B(n_1207),
.Y(n_1962)
);

BUFx3_ASAP7_75t_L g1963 ( 
.A(n_1421),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1430),
.B(n_1059),
.Y(n_1964)
);

O2A1O1Ixp5_ASAP7_75t_L g1965 ( 
.A1(n_1449),
.A2(n_1419),
.B(n_1513),
.C(n_1562),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_SL g1966 ( 
.A(n_1519),
.B(n_1662),
.Y(n_1966)
);

INVxp67_ASAP7_75t_L g1967 ( 
.A(n_1662),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1662),
.B(n_1207),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1662),
.Y(n_1969)
);

BUFx5_ASAP7_75t_L g1970 ( 
.A(n_1647),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1430),
.A2(n_1092),
.B(n_1017),
.Y(n_1971)
);

A2O1A1Ixp33_ASAP7_75t_L g1972 ( 
.A1(n_1662),
.A2(n_1430),
.B(n_1536),
.C(n_1449),
.Y(n_1972)
);

BUFx2_ASAP7_75t_L g1973 ( 
.A(n_1662),
.Y(n_1973)
);

AOI21xp5_ASAP7_75t_L g1974 ( 
.A1(n_1430),
.A2(n_1092),
.B(n_1017),
.Y(n_1974)
);

INVx1_ASAP7_75t_SL g1975 ( 
.A(n_1428),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_SL g1976 ( 
.A(n_1519),
.B(n_1662),
.Y(n_1976)
);

AOI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1430),
.A2(n_1092),
.B(n_1017),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1662),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1662),
.B(n_1207),
.Y(n_1979)
);

OAI22x1_ASAP7_75t_L g1980 ( 
.A1(n_1537),
.A2(n_1202),
.B1(n_1541),
.B2(n_1523),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1662),
.Y(n_1981)
);

AOI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1430),
.A2(n_1092),
.B(n_1017),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1662),
.B(n_1207),
.Y(n_1983)
);

A2O1A1Ixp33_ASAP7_75t_L g1984 ( 
.A1(n_1662),
.A2(n_1430),
.B(n_1536),
.C(n_1449),
.Y(n_1984)
);

OAI22x1_ASAP7_75t_L g1985 ( 
.A1(n_1537),
.A2(n_1202),
.B1(n_1541),
.B2(n_1523),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1662),
.Y(n_1986)
);

AO21x1_ASAP7_75t_L g1987 ( 
.A1(n_1567),
.A2(n_1619),
.B(n_1618),
.Y(n_1987)
);

AND2x2_ASAP7_75t_SL g1988 ( 
.A(n_1519),
.B(n_1341),
.Y(n_1988)
);

OR2x6_ASAP7_75t_L g1989 ( 
.A(n_1819),
.B(n_1944),
.Y(n_1989)
);

INVx2_ASAP7_75t_SL g1990 ( 
.A(n_1943),
.Y(n_1990)
);

INVx3_ASAP7_75t_SL g1991 ( 
.A(n_1750),
.Y(n_1991)
);

INVx2_ASAP7_75t_SL g1992 ( 
.A(n_1943),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1942),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1945),
.B(n_1950),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1960),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1668),
.Y(n_1996)
);

AO21x2_ASAP7_75t_L g1997 ( 
.A1(n_1987),
.A2(n_1745),
.B(n_1719),
.Y(n_1997)
);

AND2x4_ASAP7_75t_L g1998 ( 
.A(n_1951),
.B(n_1954),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1962),
.B(n_1968),
.Y(n_1999)
);

CKINVDCx11_ASAP7_75t_R g2000 ( 
.A(n_1817),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1937),
.Y(n_2001)
);

NOR2xp67_ASAP7_75t_L g2002 ( 
.A(n_1819),
.B(n_1671),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1979),
.B(n_1983),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1684),
.Y(n_2004)
);

NOR2xp67_ASAP7_75t_L g2005 ( 
.A(n_1671),
.B(n_1750),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_1672),
.B(n_1695),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1961),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1953),
.B(n_1960),
.Y(n_2008)
);

OA21x2_ASAP7_75t_L g2009 ( 
.A1(n_1715),
.A2(n_1729),
.B(n_1716),
.Y(n_2009)
);

NAND2x1p5_ASAP7_75t_L g2010 ( 
.A(n_1671),
.B(n_1750),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1953),
.B(n_1986),
.Y(n_2011)
);

OAI21x1_ASAP7_75t_SL g2012 ( 
.A1(n_1838),
.A2(n_1724),
.B(n_1721),
.Y(n_2012)
);

BUFx2_ASAP7_75t_L g2013 ( 
.A(n_1970),
.Y(n_2013)
);

INVx5_ASAP7_75t_L g2014 ( 
.A(n_1944),
.Y(n_2014)
);

INVx3_ASAP7_75t_L g2015 ( 
.A(n_1671),
.Y(n_2015)
);

INVxp67_ASAP7_75t_SL g2016 ( 
.A(n_1986),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1695),
.Y(n_2017)
);

AND2x4_ASAP7_75t_L g2018 ( 
.A(n_1967),
.B(n_1959),
.Y(n_2018)
);

AOI21x1_ASAP7_75t_L g2019 ( 
.A1(n_1957),
.A2(n_1976),
.B(n_1966),
.Y(n_2019)
);

AOI22xp33_ASAP7_75t_L g2020 ( 
.A1(n_1839),
.A2(n_1693),
.B1(n_1824),
.B2(n_1757),
.Y(n_2020)
);

OAI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_1967),
.A2(n_1988),
.B1(n_1888),
.B2(n_1973),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1959),
.Y(n_2022)
);

OA21x2_ASAP7_75t_L g2023 ( 
.A1(n_1715),
.A2(n_1729),
.B(n_1716),
.Y(n_2023)
);

OAI21x1_ASAP7_75t_SL g2024 ( 
.A1(n_1698),
.A2(n_1810),
.B(n_1697),
.Y(n_2024)
);

OA21x2_ASAP7_75t_L g2025 ( 
.A1(n_1736),
.A2(n_1779),
.B(n_1772),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_1744),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1981),
.Y(n_2027)
);

AOI21x1_ASAP7_75t_L g2028 ( 
.A1(n_1957),
.A2(n_1976),
.B(n_1966),
.Y(n_2028)
);

BUFx4f_ASAP7_75t_SL g2029 ( 
.A(n_1746),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_L g2030 ( 
.A(n_1733),
.B(n_1868),
.Y(n_2030)
);

OR2x2_ASAP7_75t_L g2031 ( 
.A(n_1787),
.B(n_1975),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1981),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1691),
.Y(n_2033)
);

CKINVDCx14_ASAP7_75t_R g2034 ( 
.A(n_1746),
.Y(n_2034)
);

BUFx8_ASAP7_75t_L g2035 ( 
.A(n_1970),
.Y(n_2035)
);

OAI21x1_ASAP7_75t_SL g2036 ( 
.A1(n_1807),
.A2(n_1879),
.B(n_1748),
.Y(n_2036)
);

OAI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_1956),
.A2(n_1965),
.B(n_1949),
.Y(n_2037)
);

INVx2_ASAP7_75t_SL g2038 ( 
.A(n_1970),
.Y(n_2038)
);

NAND2x1p5_ASAP7_75t_L g2039 ( 
.A(n_1827),
.B(n_1963),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1727),
.Y(n_2040)
);

BUFx3_ASAP7_75t_L g2041 ( 
.A(n_1970),
.Y(n_2041)
);

INVx2_ASAP7_75t_SL g2042 ( 
.A(n_1970),
.Y(n_2042)
);

OR2x2_ASAP7_75t_L g2043 ( 
.A(n_1787),
.B(n_1815),
.Y(n_2043)
);

BUFx3_ASAP7_75t_L g2044 ( 
.A(n_1970),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_SL g2045 ( 
.A(n_1940),
.B(n_1744),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1734),
.Y(n_2046)
);

AO21x2_ASAP7_75t_L g2047 ( 
.A1(n_1778),
.A2(n_1939),
.B(n_1686),
.Y(n_2047)
);

BUFx3_ASAP7_75t_L g2048 ( 
.A(n_1944),
.Y(n_2048)
);

BUFx2_ASAP7_75t_L g2049 ( 
.A(n_1771),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1969),
.Y(n_2050)
);

INVx6_ASAP7_75t_SL g2051 ( 
.A(n_1673),
.Y(n_2051)
);

BUFx2_ASAP7_75t_L g2052 ( 
.A(n_1771),
.Y(n_2052)
);

OAI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_1988),
.A2(n_1888),
.B1(n_1755),
.B2(n_1927),
.Y(n_2053)
);

CKINVDCx20_ASAP7_75t_R g2054 ( 
.A(n_1732),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1878),
.B(n_1757),
.Y(n_2055)
);

AO21x2_ASAP7_75t_L g2056 ( 
.A1(n_1688),
.A2(n_1901),
.B(n_1891),
.Y(n_2056)
);

OAI21xp5_ASAP7_75t_L g2057 ( 
.A1(n_1946),
.A2(n_1974),
.B(n_1971),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_SL g2058 ( 
.A(n_1762),
.B(n_1833),
.Y(n_2058)
);

AOI22x1_ASAP7_75t_L g2059 ( 
.A1(n_1980),
.A2(n_1985),
.B1(n_1848),
.B2(n_1826),
.Y(n_2059)
);

BUFx12f_ASAP7_75t_L g2060 ( 
.A(n_1846),
.Y(n_2060)
);

AOI22xp33_ASAP7_75t_L g2061 ( 
.A1(n_1839),
.A2(n_1871),
.B1(n_1903),
.B2(n_1947),
.Y(n_2061)
);

OAI21x1_ASAP7_75t_SL g2062 ( 
.A1(n_1898),
.A2(n_1781),
.B(n_1677),
.Y(n_2062)
);

CKINVDCx20_ASAP7_75t_R g2063 ( 
.A(n_1963),
.Y(n_2063)
);

OAI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_1977),
.A2(n_1982),
.B(n_1972),
.Y(n_2064)
);

O2A1O1Ixp33_ASAP7_75t_L g2065 ( 
.A1(n_1764),
.A2(n_1899),
.B(n_1972),
.C(n_1952),
.Y(n_2065)
);

INVx3_ASAP7_75t_L g2066 ( 
.A(n_1827),
.Y(n_2066)
);

BUFx4f_ASAP7_75t_L g2067 ( 
.A(n_1762),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_1673),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1720),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1700),
.B(n_1978),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_1948),
.B(n_1964),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1720),
.Y(n_2072)
);

INVxp67_ASAP7_75t_SL g2073 ( 
.A(n_1882),
.Y(n_2073)
);

NOR2x1_ASAP7_75t_SL g2074 ( 
.A(n_1900),
.B(n_1911),
.Y(n_2074)
);

BUFx2_ASAP7_75t_L g2075 ( 
.A(n_1674),
.Y(n_2075)
);

OA21x2_ASAP7_75t_L g2076 ( 
.A1(n_1821),
.A2(n_1984),
.B(n_1893),
.Y(n_2076)
);

AO21x2_ASAP7_75t_L g2077 ( 
.A1(n_1917),
.A2(n_1894),
.B(n_1870),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_1681),
.B(n_1790),
.Y(n_2078)
);

BUFx3_ASAP7_75t_L g2079 ( 
.A(n_1666),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_1678),
.Y(n_2080)
);

OR2x6_ASAP7_75t_L g2081 ( 
.A(n_1915),
.B(n_1756),
.Y(n_2081)
);

NOR2xp33_ASAP7_75t_L g2082 ( 
.A(n_1964),
.B(n_1847),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1818),
.B(n_1752),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_1673),
.Y(n_2084)
);

NOR2xp67_ASAP7_75t_SL g2085 ( 
.A(n_1900),
.B(n_1911),
.Y(n_2085)
);

OAI21x1_ASAP7_75t_SL g2086 ( 
.A1(n_1914),
.A2(n_1789),
.B(n_1783),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1774),
.Y(n_2087)
);

NOR2xp67_ASAP7_75t_L g2088 ( 
.A(n_1828),
.B(n_1678),
.Y(n_2088)
);

NAND2x1p5_ASAP7_75t_L g2089 ( 
.A(n_1900),
.B(n_1915),
.Y(n_2089)
);

OAI21x1_ASAP7_75t_SL g2090 ( 
.A1(n_1792),
.A2(n_1842),
.B(n_1843),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1775),
.Y(n_2091)
);

OAI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_1761),
.A2(n_1742),
.B(n_1718),
.Y(n_2092)
);

AOI22x1_ASAP7_75t_L g2093 ( 
.A1(n_1916),
.A2(n_1822),
.B1(n_1875),
.B2(n_1798),
.Y(n_2093)
);

AOI22xp5_ASAP7_75t_L g2094 ( 
.A1(n_1847),
.A2(n_1885),
.B1(n_1770),
.B2(n_1845),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1801),
.Y(n_2095)
);

OA21x2_ASAP7_75t_L g2096 ( 
.A1(n_1676),
.A2(n_1692),
.B(n_1670),
.Y(n_2096)
);

BUFx2_ASAP7_75t_R g2097 ( 
.A(n_1920),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1802),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1808),
.Y(n_2099)
);

INVx3_ASAP7_75t_L g2100 ( 
.A(n_1666),
.Y(n_2100)
);

NOR2xp33_ASAP7_75t_L g2101 ( 
.A(n_1854),
.B(n_1857),
.Y(n_2101)
);

AOI21xp5_ASAP7_75t_L g2102 ( 
.A1(n_1882),
.A2(n_1823),
.B(n_1812),
.Y(n_2102)
);

NOR2x1_ASAP7_75t_R g2103 ( 
.A(n_1915),
.B(n_1804),
.Y(n_2103)
);

AO21x2_ASAP7_75t_L g2104 ( 
.A1(n_1692),
.A2(n_1861),
.B(n_1859),
.Y(n_2104)
);

BUFx12f_ASAP7_75t_L g2105 ( 
.A(n_1759),
.Y(n_2105)
);

NAND2x1p5_ASAP7_75t_L g2106 ( 
.A(n_1900),
.B(n_1958),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1760),
.Y(n_2107)
);

CKINVDCx6p67_ASAP7_75t_R g2108 ( 
.A(n_1785),
.Y(n_2108)
);

OAI21x1_ASAP7_75t_SL g2109 ( 
.A1(n_1765),
.A2(n_1777),
.B(n_1769),
.Y(n_2109)
);

OAI21xp5_ASAP7_75t_L g2110 ( 
.A1(n_1761),
.A2(n_1718),
.B(n_1667),
.Y(n_2110)
);

AND2x4_ASAP7_75t_L g2111 ( 
.A(n_1941),
.B(n_1911),
.Y(n_2111)
);

OAI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_1844),
.A2(n_1905),
.B(n_1687),
.Y(n_2112)
);

OAI21x1_ASAP7_75t_SL g2113 ( 
.A1(n_1904),
.A2(n_1799),
.B(n_1941),
.Y(n_2113)
);

INVx4_ASAP7_75t_SL g2114 ( 
.A(n_1912),
.Y(n_2114)
);

NOR2xp33_ASAP7_75t_L g2115 ( 
.A(n_1864),
.B(n_1845),
.Y(n_2115)
);

BUFx2_ASAP7_75t_SL g2116 ( 
.A(n_1785),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_1668),
.Y(n_2117)
);

AO21x2_ASAP7_75t_L g2118 ( 
.A1(n_1670),
.A2(n_1669),
.B(n_1883),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1699),
.B(n_1712),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1911),
.B(n_1941),
.Y(n_2120)
);

AOI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_1840),
.A2(n_1851),
.B1(n_1906),
.B2(n_1814),
.Y(n_2121)
);

OR3x4_ASAP7_75t_SL g2122 ( 
.A(n_1723),
.B(n_1796),
.C(n_1835),
.Y(n_2122)
);

CKINVDCx20_ASAP7_75t_R g2123 ( 
.A(n_1828),
.Y(n_2123)
);

AO21x2_ASAP7_75t_L g2124 ( 
.A1(n_1841),
.A2(n_1834),
.B(n_1696),
.Y(n_2124)
);

INVx6_ASAP7_75t_L g2125 ( 
.A(n_1785),
.Y(n_2125)
);

BUFx8_ASAP7_75t_SL g2126 ( 
.A(n_1865),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1800),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1705),
.Y(n_2128)
);

INVx1_ASAP7_75t_SL g2129 ( 
.A(n_1805),
.Y(n_2129)
);

HB1xp67_ASAP7_75t_L g2130 ( 
.A(n_1805),
.Y(n_2130)
);

BUFx2_ASAP7_75t_L g2131 ( 
.A(n_1805),
.Y(n_2131)
);

OR2x2_ASAP7_75t_L g2132 ( 
.A(n_1685),
.B(n_1737),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1735),
.Y(n_2133)
);

NOR2xp33_ASAP7_75t_L g2134 ( 
.A(n_1728),
.B(n_1835),
.Y(n_2134)
);

OAI21xp5_ASAP7_75t_L g2135 ( 
.A1(n_1907),
.A2(n_1933),
.B(n_1926),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1938),
.Y(n_2136)
);

OA21x2_ASAP7_75t_L g2137 ( 
.A1(n_1919),
.A2(n_1806),
.B(n_1731),
.Y(n_2137)
);

INVx3_ASAP7_75t_L g2138 ( 
.A(n_1958),
.Y(n_2138)
);

HB1xp67_ASAP7_75t_L g2139 ( 
.A(n_1756),
.Y(n_2139)
);

OR2x2_ASAP7_75t_L g2140 ( 
.A(n_1689),
.B(n_1782),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1708),
.B(n_1863),
.Y(n_2141)
);

INVx4_ASAP7_75t_SL g2142 ( 
.A(n_1912),
.Y(n_2142)
);

CKINVDCx14_ASAP7_75t_R g2143 ( 
.A(n_1912),
.Y(n_2143)
);

OAI21xp5_ASAP7_75t_L g2144 ( 
.A1(n_1749),
.A2(n_1753),
.B(n_1747),
.Y(n_2144)
);

INVx3_ASAP7_75t_L g2145 ( 
.A(n_1694),
.Y(n_2145)
);

CKINVDCx20_ASAP7_75t_R g2146 ( 
.A(n_1768),
.Y(n_2146)
);

AO21x2_ASAP7_75t_L g2147 ( 
.A1(n_1834),
.A2(n_1696),
.B(n_1858),
.Y(n_2147)
);

CKINVDCx16_ASAP7_75t_R g2148 ( 
.A(n_1912),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1892),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1803),
.B(n_1853),
.Y(n_2150)
);

NAND2x1p5_ASAP7_75t_L g2151 ( 
.A(n_1768),
.B(n_1811),
.Y(n_2151)
);

AO21x2_ASAP7_75t_L g2152 ( 
.A1(n_1858),
.A2(n_1849),
.B(n_1682),
.Y(n_2152)
);

AOI22x1_ASAP7_75t_L g2153 ( 
.A1(n_1916),
.A2(n_1809),
.B1(n_1866),
.B2(n_1754),
.Y(n_2153)
);

INVx4_ASAP7_75t_L g2154 ( 
.A(n_1811),
.Y(n_2154)
);

OR2x6_ASAP7_75t_L g2155 ( 
.A(n_1784),
.B(n_1892),
.Y(n_2155)
);

OAI21x1_ASAP7_75t_L g2156 ( 
.A1(n_1717),
.A2(n_1791),
.B(n_1837),
.Y(n_2156)
);

OAI21x1_ASAP7_75t_L g2157 ( 
.A1(n_1791),
.A2(n_1837),
.B(n_1704),
.Y(n_2157)
);

OAI21x1_ASAP7_75t_L g2158 ( 
.A1(n_1922),
.A2(n_1852),
.B(n_1730),
.Y(n_2158)
);

BUFx2_ASAP7_75t_L g2159 ( 
.A(n_1912),
.Y(n_2159)
);

INVx1_ASAP7_75t_SL g2160 ( 
.A(n_1908),
.Y(n_2160)
);

OA21x2_ASAP7_75t_L g2161 ( 
.A1(n_1773),
.A2(n_1852),
.B(n_1921),
.Y(n_2161)
);

INVx6_ASAP7_75t_SL g2162 ( 
.A(n_1865),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_1850),
.B(n_1902),
.Y(n_2163)
);

AO21x2_ASAP7_75t_L g2164 ( 
.A1(n_1876),
.A2(n_1820),
.B(n_1836),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_1865),
.Y(n_2165)
);

AO21x2_ASAP7_75t_L g2166 ( 
.A1(n_1876),
.A2(n_1832),
.B(n_1713),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1690),
.Y(n_2167)
);

OAI221xp5_ASAP7_75t_L g2168 ( 
.A1(n_1825),
.A2(n_1797),
.B1(n_1816),
.B2(n_1814),
.C(n_1889),
.Y(n_2168)
);

NAND3xp33_ASAP7_75t_L g2169 ( 
.A(n_1825),
.B(n_1923),
.C(n_1713),
.Y(n_2169)
);

OA21x2_ASAP7_75t_L g2170 ( 
.A1(n_1706),
.A2(n_1925),
.B(n_1923),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_1862),
.B(n_1813),
.Y(n_2171)
);

OAI221xp5_ASAP7_75t_SL g2172 ( 
.A1(n_1683),
.A2(n_1710),
.B1(n_1925),
.B2(n_1706),
.C(n_1793),
.Y(n_2172)
);

CKINVDCx5p33_ASAP7_75t_R g2173 ( 
.A(n_1856),
.Y(n_2173)
);

OAI21x1_ASAP7_75t_L g2174 ( 
.A1(n_1722),
.A2(n_1725),
.B(n_1751),
.Y(n_2174)
);

BUFx3_ASAP7_75t_L g2175 ( 
.A(n_1705),
.Y(n_2175)
);

BUFx12f_ASAP7_75t_L g2176 ( 
.A(n_1886),
.Y(n_2176)
);

OAI21x1_ASAP7_75t_L g2177 ( 
.A1(n_1722),
.A2(n_1743),
.B(n_1741),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1680),
.Y(n_2178)
);

OAI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_1890),
.A2(n_1913),
.B(n_1831),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1910),
.Y(n_2180)
);

INVx4_ASAP7_75t_L g2181 ( 
.A(n_1873),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1726),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1767),
.B(n_1795),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1880),
.B(n_1897),
.Y(n_2184)
);

CKINVDCx5p33_ASAP7_75t_R g2185 ( 
.A(n_1766),
.Y(n_2185)
);

OAI21x1_ASAP7_75t_L g2186 ( 
.A1(n_1703),
.A2(n_1869),
.B(n_1867),
.Y(n_2186)
);

AO21x2_ASAP7_75t_L g2187 ( 
.A1(n_1918),
.A2(n_1707),
.B(n_1711),
.Y(n_2187)
);

BUFx2_ASAP7_75t_SL g2188 ( 
.A(n_1763),
.Y(n_2188)
);

NOR2x1_ASAP7_75t_SL g2189 ( 
.A(n_1855),
.B(n_1786),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1887),
.Y(n_2190)
);

OA21x2_ASAP7_75t_L g2191 ( 
.A1(n_1829),
.A2(n_1830),
.B(n_1860),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1931),
.Y(n_2192)
);

AND2x4_ASAP7_75t_L g2193 ( 
.A(n_1909),
.B(n_1897),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1887),
.Y(n_2194)
);

OAI21xp5_ASAP7_75t_L g2195 ( 
.A1(n_1794),
.A2(n_1788),
.B(n_1780),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1675),
.Y(n_2196)
);

OA21x2_ASAP7_75t_L g2197 ( 
.A1(n_1924),
.A2(n_1936),
.B(n_1934),
.Y(n_2197)
);

OAI21x1_ASAP7_75t_L g2198 ( 
.A1(n_1928),
.A2(n_1930),
.B(n_1929),
.Y(n_2198)
);

INVx6_ASAP7_75t_L g2199 ( 
.A(n_1873),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_1881),
.B(n_1739),
.Y(n_2200)
);

OAI21x1_ASAP7_75t_L g2201 ( 
.A1(n_1932),
.A2(n_1709),
.B(n_1740),
.Y(n_2201)
);

INVxp67_ASAP7_75t_SL g2202 ( 
.A(n_1855),
.Y(n_2202)
);

NOR2xp67_ASAP7_75t_L g2203 ( 
.A(n_1776),
.B(n_1896),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1758),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1887),
.Y(n_2205)
);

OAI21x1_ASAP7_75t_L g2206 ( 
.A1(n_1877),
.A2(n_1874),
.B(n_1895),
.Y(n_2206)
);

OAI21x1_ASAP7_75t_L g2207 ( 
.A1(n_1738),
.A2(n_1723),
.B(n_1897),
.Y(n_2207)
);

AO21x2_ASAP7_75t_L g2208 ( 
.A1(n_1679),
.A2(n_1897),
.B(n_1701),
.Y(n_2208)
);

OA21x2_ASAP7_75t_L g2209 ( 
.A1(n_1701),
.A2(n_1935),
.B(n_1739),
.Y(n_2209)
);

OAI21x1_ASAP7_75t_L g2210 ( 
.A1(n_1701),
.A2(n_1935),
.B(n_1739),
.Y(n_2210)
);

OAI21x1_ASAP7_75t_L g2211 ( 
.A1(n_1701),
.A2(n_1935),
.B(n_1739),
.Y(n_2211)
);

INVx6_ASAP7_75t_L g2212 ( 
.A(n_1702),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1942),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_1961),
.B(n_1192),
.Y(n_2214)
);

AO31x2_ASAP7_75t_L g2215 ( 
.A1(n_1987),
.A2(n_1778),
.A3(n_1714),
.B(n_1952),
.Y(n_2215)
);

AOI22x1_ASAP7_75t_L g2216 ( 
.A1(n_1980),
.A2(n_1985),
.B1(n_1624),
.B2(n_1955),
.Y(n_2216)
);

INVx3_ASAP7_75t_L g2217 ( 
.A(n_1671),
.Y(n_2217)
);

NOR2xp67_ASAP7_75t_L g2218 ( 
.A(n_1819),
.B(n_1246),
.Y(n_2218)
);

INVx5_ASAP7_75t_L g2219 ( 
.A(n_1944),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1942),
.Y(n_2220)
);

INVx4_ASAP7_75t_L g2221 ( 
.A(n_1819),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1937),
.Y(n_2222)
);

INVx3_ASAP7_75t_L g2223 ( 
.A(n_1671),
.Y(n_2223)
);

AOI21x1_ASAP7_75t_SL g2224 ( 
.A1(n_1889),
.A2(n_1872),
.B(n_1884),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_1961),
.B(n_1192),
.Y(n_2225)
);

NOR2xp67_ASAP7_75t_L g2226 ( 
.A(n_1819),
.B(n_1246),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1942),
.Y(n_2227)
);

OR2x2_ASAP7_75t_L g2228 ( 
.A(n_1684),
.B(n_1389),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1937),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1942),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1942),
.Y(n_2231)
);

HB1xp67_ASAP7_75t_L g2232 ( 
.A(n_1960),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1942),
.B(n_1662),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1942),
.Y(n_2234)
);

BUFx2_ASAP7_75t_R g2235 ( 
.A(n_1744),
.Y(n_2235)
);

HB1xp67_ASAP7_75t_L g2236 ( 
.A(n_1960),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_1961),
.B(n_1192),
.Y(n_2237)
);

BUFx6f_ASAP7_75t_L g2238 ( 
.A(n_1668),
.Y(n_2238)
);

INVx6_ASAP7_75t_L g2239 ( 
.A(n_1671),
.Y(n_2239)
);

OR2x2_ASAP7_75t_L g2240 ( 
.A(n_2006),
.B(n_1994),
.Y(n_2240)
);

AOI22xp33_ASAP7_75t_SL g2241 ( 
.A1(n_2199),
.A2(n_2143),
.B1(n_2181),
.B2(n_2067),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2007),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2050),
.Y(n_2243)
);

BUFx12f_ASAP7_75t_L g2244 ( 
.A(n_2000),
.Y(n_2244)
);

BUFx2_ASAP7_75t_L g2245 ( 
.A(n_2035),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2033),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2214),
.B(n_2225),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2040),
.Y(n_2248)
);

AOI22xp33_ASAP7_75t_SL g2249 ( 
.A1(n_2199),
.A2(n_2143),
.B1(n_2181),
.B2(n_2067),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2046),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2237),
.B(n_1994),
.Y(n_2251)
);

HB1xp67_ASAP7_75t_L g2252 ( 
.A(n_1995),
.Y(n_2252)
);

HB1xp67_ASAP7_75t_L g2253 ( 
.A(n_1995),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2087),
.Y(n_2254)
);

AOI22xp33_ASAP7_75t_L g2255 ( 
.A1(n_2199),
.A2(n_2020),
.B1(n_2055),
.B2(n_2061),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_1998),
.B(n_1999),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_1998),
.B(n_1999),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1998),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2091),
.Y(n_2259)
);

BUFx6f_ASAP7_75t_L g2260 ( 
.A(n_1996),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2003),
.Y(n_2261)
);

BUFx2_ASAP7_75t_L g2262 ( 
.A(n_2035),
.Y(n_2262)
);

AND2x4_ASAP7_75t_L g2263 ( 
.A(n_2114),
.B(n_2142),
.Y(n_2263)
);

INVx3_ASAP7_75t_L g2264 ( 
.A(n_2035),
.Y(n_2264)
);

HB1xp67_ASAP7_75t_L g2265 ( 
.A(n_2232),
.Y(n_2265)
);

INVx2_ASAP7_75t_SL g2266 ( 
.A(n_1991),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2017),
.Y(n_2267)
);

BUFx2_ASAP7_75t_SL g2268 ( 
.A(n_2002),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2107),
.Y(n_2269)
);

INVxp67_ASAP7_75t_L g2270 ( 
.A(n_2232),
.Y(n_2270)
);

AOI22xp33_ASAP7_75t_SL g2271 ( 
.A1(n_2148),
.A2(n_2116),
.B1(n_2058),
.B2(n_2212),
.Y(n_2271)
);

AO21x1_ASAP7_75t_SL g2272 ( 
.A1(n_2130),
.A2(n_2139),
.B(n_2084),
.Y(n_2272)
);

CKINVDCx20_ASAP7_75t_R g2273 ( 
.A(n_2029),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1993),
.Y(n_2274)
);

INVx3_ASAP7_75t_L g2275 ( 
.A(n_2041),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2213),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2220),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2227),
.Y(n_2278)
);

OAI22xp5_ASAP7_75t_L g2279 ( 
.A1(n_2108),
.A2(n_2020),
.B1(n_2061),
.B2(n_2125),
.Y(n_2279)
);

BUFx3_ASAP7_75t_L g2280 ( 
.A(n_2010),
.Y(n_2280)
);

BUFx4f_ASAP7_75t_SL g2281 ( 
.A(n_2221),
.Y(n_2281)
);

BUFx2_ASAP7_75t_R g2282 ( 
.A(n_2026),
.Y(n_2282)
);

AO21x1_ASAP7_75t_L g2283 ( 
.A1(n_2053),
.A2(n_2021),
.B(n_2102),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2230),
.Y(n_2284)
);

HB1xp67_ASAP7_75t_L g2285 ( 
.A(n_2236),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2231),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2234),
.B(n_2070),
.Y(n_2287)
);

BUFx8_ASAP7_75t_SL g2288 ( 
.A(n_2026),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2236),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2095),
.Y(n_2290)
);

AOI221xp5_ASAP7_75t_L g2291 ( 
.A1(n_2030),
.A2(n_2101),
.B1(n_2082),
.B2(n_2115),
.C(n_2092),
.Y(n_2291)
);

NOR2x1_ASAP7_75t_R g2292 ( 
.A(n_2000),
.B(n_2221),
.Y(n_2292)
);

BUFx3_ASAP7_75t_L g2293 ( 
.A(n_2010),
.Y(n_2293)
);

CKINVDCx20_ASAP7_75t_R g2294 ( 
.A(n_2029),
.Y(n_2294)
);

INVx3_ASAP7_75t_L g2295 ( 
.A(n_2041),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2098),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2099),
.Y(n_2297)
);

OR2x6_ASAP7_75t_L g2298 ( 
.A(n_2125),
.B(n_2159),
.Y(n_2298)
);

AOI221xp5_ASAP7_75t_L g2299 ( 
.A1(n_2030),
.A2(n_2101),
.B1(n_2082),
.B2(n_2115),
.C(n_2169),
.Y(n_2299)
);

AOI22xp33_ASAP7_75t_L g2300 ( 
.A1(n_2212),
.A2(n_2173),
.B1(n_2168),
.B2(n_2204),
.Y(n_2300)
);

BUFx12f_ASAP7_75t_L g2301 ( 
.A(n_1990),
.Y(n_2301)
);

NAND2xp33_ASAP7_75t_R g2302 ( 
.A(n_2131),
.B(n_2114),
.Y(n_2302)
);

INVx1_ASAP7_75t_SL g2303 ( 
.A(n_1991),
.Y(n_2303)
);

BUFx2_ASAP7_75t_L g2304 ( 
.A(n_2063),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2004),
.Y(n_2305)
);

OAI22xp5_ASAP7_75t_L g2306 ( 
.A1(n_2125),
.A2(n_2130),
.B1(n_2016),
.B2(n_2073),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2233),
.Y(n_2307)
);

INVx1_ASAP7_75t_SL g2308 ( 
.A(n_2054),
.Y(n_2308)
);

BUFx12f_ASAP7_75t_L g2309 ( 
.A(n_1992),
.Y(n_2309)
);

CKINVDCx11_ASAP7_75t_R g2310 ( 
.A(n_2054),
.Y(n_2310)
);

OAI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_2185),
.A2(n_2129),
.B1(n_2011),
.B2(n_2008),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2127),
.Y(n_2312)
);

INVx3_ASAP7_75t_L g2313 ( 
.A(n_2044),
.Y(n_2313)
);

AOI22xp33_ASAP7_75t_L g2314 ( 
.A1(n_2212),
.A2(n_2173),
.B1(n_2192),
.B2(n_2182),
.Y(n_2314)
);

AOI22xp33_ASAP7_75t_L g2315 ( 
.A1(n_2094),
.A2(n_2110),
.B1(n_2196),
.B2(n_2185),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2001),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2022),
.Y(n_2317)
);

INVxp67_ASAP7_75t_L g2318 ( 
.A(n_2013),
.Y(n_2318)
);

BUFx6f_ASAP7_75t_SL g2319 ( 
.A(n_1989),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2022),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2112),
.B(n_2065),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2027),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2032),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2032),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2222),
.Y(n_2325)
);

HB1xp67_ASAP7_75t_L g2326 ( 
.A(n_2068),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2083),
.B(n_2018),
.Y(n_2327)
);

AND2x4_ASAP7_75t_L g2328 ( 
.A(n_2114),
.B(n_2142),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2229),
.Y(n_2329)
);

INVx3_ASAP7_75t_L g2330 ( 
.A(n_2239),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2018),
.Y(n_2331)
);

HB1xp67_ASAP7_75t_L g2332 ( 
.A(n_2084),
.Y(n_2332)
);

OAI22xp5_ASAP7_75t_L g2333 ( 
.A1(n_2121),
.A2(n_2155),
.B1(n_2051),
.B2(n_2081),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2078),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2178),
.Y(n_2335)
);

OR2x2_ASAP7_75t_L g2336 ( 
.A(n_2228),
.B(n_2075),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2005),
.B(n_2160),
.Y(n_2337)
);

HB1xp67_ASAP7_75t_L g2338 ( 
.A(n_2174),
.Y(n_2338)
);

NAND2x1p5_ASAP7_75t_L g2339 ( 
.A(n_2014),
.B(n_2219),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2069),
.Y(n_2340)
);

AOI22xp33_ASAP7_75t_L g2341 ( 
.A1(n_2071),
.A2(n_2036),
.B1(n_2134),
.B2(n_2090),
.Y(n_2341)
);

AOI22xp33_ASAP7_75t_SL g2342 ( 
.A1(n_2139),
.A2(n_2012),
.B1(n_2109),
.B2(n_2165),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2069),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2072),
.Y(n_2344)
);

OAI22xp5_ASAP7_75t_L g2345 ( 
.A1(n_2155),
.A2(n_2051),
.B1(n_2081),
.B2(n_2123),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2072),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2134),
.B(n_2071),
.Y(n_2347)
);

OR2x6_ASAP7_75t_L g2348 ( 
.A(n_1989),
.B(n_2081),
.Y(n_2348)
);

HB1xp67_ASAP7_75t_L g2349 ( 
.A(n_2174),
.Y(n_2349)
);

INVxp67_ASAP7_75t_L g2350 ( 
.A(n_2038),
.Y(n_2350)
);

CKINVDCx9p33_ASAP7_75t_R g2351 ( 
.A(n_2142),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2180),
.Y(n_2352)
);

AOI22xp33_ASAP7_75t_L g2353 ( 
.A1(n_2136),
.A2(n_2147),
.B1(n_2133),
.B2(n_2170),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2171),
.B(n_2183),
.Y(n_2354)
);

NAND2x1p5_ASAP7_75t_L g2355 ( 
.A(n_2014),
.B(n_2219),
.Y(n_2355)
);

INVx2_ASAP7_75t_SL g2356 ( 
.A(n_1989),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2150),
.B(n_2141),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2042),
.Y(n_2358)
);

HB1xp67_ASAP7_75t_L g2359 ( 
.A(n_2177),
.Y(n_2359)
);

AO31x2_ASAP7_75t_L g2360 ( 
.A1(n_2190),
.A2(n_2205),
.A3(n_2194),
.B(n_2184),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2043),
.Y(n_2361)
);

INVx4_ASAP7_75t_SL g2362 ( 
.A(n_2239),
.Y(n_2362)
);

OAI22xp33_ASAP7_75t_L g2363 ( 
.A1(n_2155),
.A2(n_2165),
.B1(n_2051),
.B2(n_2162),
.Y(n_2363)
);

AND2x4_ASAP7_75t_L g2364 ( 
.A(n_2014),
.B(n_2219),
.Y(n_2364)
);

OAI22xp5_ASAP7_75t_L g2365 ( 
.A1(n_2123),
.A2(n_2172),
.B1(n_2119),
.B2(n_2149),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2218),
.B(n_2226),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2031),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2167),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2015),
.Y(n_2369)
);

AO21x1_ASAP7_75t_SL g2370 ( 
.A1(n_2162),
.A2(n_2074),
.B(n_2085),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2015),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2217),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2217),
.Y(n_2373)
);

INVx4_ASAP7_75t_L g2374 ( 
.A(n_2014),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2223),
.Y(n_2375)
);

BUFx2_ASAP7_75t_L g2376 ( 
.A(n_2063),
.Y(n_2376)
);

INVx3_ASAP7_75t_L g2377 ( 
.A(n_2239),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2223),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2088),
.Y(n_2379)
);

BUFx10_ASAP7_75t_L g2380 ( 
.A(n_2045),
.Y(n_2380)
);

BUFx3_ASAP7_75t_L g2381 ( 
.A(n_2146),
.Y(n_2381)
);

AOI21xp5_ASAP7_75t_L g2382 ( 
.A1(n_2037),
.A2(n_2064),
.B(n_2057),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2210),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2211),
.Y(n_2384)
);

OR2x6_ASAP7_75t_L g2385 ( 
.A(n_2120),
.B(n_2089),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_2146),
.B(n_2140),
.Y(n_2386)
);

OR2x2_ASAP7_75t_L g2387 ( 
.A(n_2049),
.B(n_2052),
.Y(n_2387)
);

INVx3_ASAP7_75t_L g2388 ( 
.A(n_2219),
.Y(n_2388)
);

OAI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_2211),
.A2(n_2158),
.B(n_2135),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2024),
.Y(n_2390)
);

OAI22xp5_ASAP7_75t_L g2391 ( 
.A1(n_2162),
.A2(n_2170),
.B1(n_2132),
.B2(n_2193),
.Y(n_2391)
);

AOI22xp33_ASAP7_75t_L g2392 ( 
.A1(n_2147),
.A2(n_2170),
.B1(n_2200),
.B2(n_2176),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2209),
.Y(n_2393)
);

CKINVDCx14_ASAP7_75t_R g2394 ( 
.A(n_2034),
.Y(n_2394)
);

INVx2_ASAP7_75t_SL g2395 ( 
.A(n_2060),
.Y(n_2395)
);

HB1xp67_ASAP7_75t_L g2396 ( 
.A(n_2175),
.Y(n_2396)
);

BUFx2_ASAP7_75t_L g2397 ( 
.A(n_2126),
.Y(n_2397)
);

OAI22xp5_ASAP7_75t_L g2398 ( 
.A1(n_2193),
.A2(n_2137),
.B1(n_2097),
.B2(n_2096),
.Y(n_2398)
);

AOI22xp5_ASAP7_75t_L g2399 ( 
.A1(n_2176),
.A2(n_2105),
.B1(n_2034),
.B2(n_2193),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2066),
.Y(n_2400)
);

HB1xp67_ASAP7_75t_L g2401 ( 
.A(n_2175),
.Y(n_2401)
);

INVx2_ASAP7_75t_SL g2402 ( 
.A(n_2060),
.Y(n_2402)
);

BUFx3_ASAP7_75t_L g2403 ( 
.A(n_2039),
.Y(n_2403)
);

AOI22xp33_ASAP7_75t_SL g2404 ( 
.A1(n_2189),
.A2(n_2062),
.B1(n_2086),
.B2(n_2216),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_2048),
.B(n_2105),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2080),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2080),
.Y(n_2407)
);

AOI22xp5_ASAP7_75t_L g2408 ( 
.A1(n_2124),
.A2(n_2144),
.B1(n_2179),
.B2(n_2187),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2188),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2103),
.Y(n_2410)
);

OAI22xp33_ASAP7_75t_L g2411 ( 
.A1(n_2122),
.A2(n_2137),
.B1(n_2096),
.B2(n_2089),
.Y(n_2411)
);

AOI22xp33_ASAP7_75t_L g2412 ( 
.A1(n_2124),
.A2(n_2104),
.B1(n_2152),
.B2(n_2153),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2100),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2307),
.B(n_2208),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2251),
.B(n_2039),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2247),
.B(n_2079),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2274),
.Y(n_2417)
);

OR2x2_ASAP7_75t_L g2418 ( 
.A(n_2240),
.B(n_2208),
.Y(n_2418)
);

BUFx3_ASAP7_75t_L g2419 ( 
.A(n_2245),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2392),
.B(n_2056),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2276),
.Y(n_2421)
);

HB1xp67_ASAP7_75t_L g2422 ( 
.A(n_2252),
.Y(n_2422)
);

HB1xp67_ASAP7_75t_L g2423 ( 
.A(n_2252),
.Y(n_2423)
);

BUFx4f_ASAP7_75t_L g2424 ( 
.A(n_2262),
.Y(n_2424)
);

INVx2_ASAP7_75t_SL g2425 ( 
.A(n_2264),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2287),
.B(n_2327),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2256),
.B(n_2079),
.Y(n_2427)
);

AOI22xp33_ASAP7_75t_L g2428 ( 
.A1(n_2299),
.A2(n_2104),
.B1(n_2187),
.B2(n_2118),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2277),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2299),
.B(n_2163),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2392),
.B(n_2056),
.Y(n_2431)
);

AND2x2_ASAP7_75t_L g2432 ( 
.A(n_2347),
.B(n_2154),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2386),
.B(n_2154),
.Y(n_2433)
);

AOI22xp33_ASAP7_75t_SL g2434 ( 
.A1(n_2365),
.A2(n_2113),
.B1(n_2059),
.B2(n_2093),
.Y(n_2434)
);

AND2x4_ASAP7_75t_SL g2435 ( 
.A(n_2264),
.B(n_2263),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2360),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2278),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2360),
.Y(n_2438)
);

OAI21xp5_ASAP7_75t_SL g2439 ( 
.A1(n_2241),
.A2(n_2111),
.B(n_2122),
.Y(n_2439)
);

BUFx3_ASAP7_75t_L g2440 ( 
.A(n_2280),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2357),
.B(n_2151),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2334),
.B(n_2151),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2360),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2284),
.Y(n_2444)
);

AND2x4_ASAP7_75t_L g2445 ( 
.A(n_2263),
.B(n_2111),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2286),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2243),
.Y(n_2447)
);

OR2x2_ASAP7_75t_L g2448 ( 
.A(n_2257),
.B(n_2215),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2291),
.B(n_2152),
.Y(n_2449)
);

AND2x2_ASAP7_75t_L g2450 ( 
.A(n_2361),
.B(n_2138),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2246),
.Y(n_2451)
);

INVx3_ASAP7_75t_L g2452 ( 
.A(n_2328),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2367),
.B(n_2207),
.Y(n_2453)
);

BUFx3_ASAP7_75t_L g2454 ( 
.A(n_2280),
.Y(n_2454)
);

OR2x2_ASAP7_75t_L g2455 ( 
.A(n_2257),
.B(n_2253),
.Y(n_2455)
);

HB1xp67_ASAP7_75t_L g2456 ( 
.A(n_2253),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2381),
.B(n_2207),
.Y(n_2457)
);

AND2x2_ASAP7_75t_L g2458 ( 
.A(n_2381),
.B(n_2077),
.Y(n_2458)
);

OR2x2_ASAP7_75t_L g2459 ( 
.A(n_2265),
.B(n_2215),
.Y(n_2459)
);

AND2x4_ASAP7_75t_SL g2460 ( 
.A(n_2328),
.B(n_2111),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2248),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2291),
.B(n_2077),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2393),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2303),
.B(n_2145),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2250),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2254),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2259),
.Y(n_2467)
);

HB1xp67_ASAP7_75t_L g2468 ( 
.A(n_2285),
.Y(n_2468)
);

AOI22xp33_ASAP7_75t_L g2469 ( 
.A1(n_2365),
.A2(n_2118),
.B1(n_2195),
.B2(n_2096),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2269),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2242),
.Y(n_2471)
);

INVx2_ASAP7_75t_SL g2472 ( 
.A(n_2293),
.Y(n_2472)
);

OAI21xp33_ASAP7_75t_L g2473 ( 
.A1(n_2255),
.A2(n_2341),
.B(n_2279),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2353),
.B(n_1997),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2267),
.Y(n_2475)
);

OAI222xp33_ASAP7_75t_L g2476 ( 
.A1(n_2333),
.A2(n_2120),
.B1(n_2202),
.B2(n_2028),
.C1(n_2019),
.C2(n_2106),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2352),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2304),
.B(n_2145),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2315),
.B(n_2166),
.Y(n_2479)
);

AND2x2_ASAP7_75t_L g2480 ( 
.A(n_2376),
.B(n_2266),
.Y(n_2480)
);

AND2x4_ASAP7_75t_L g2481 ( 
.A(n_2390),
.B(n_1997),
.Y(n_2481)
);

BUFx3_ASAP7_75t_L g2482 ( 
.A(n_2293),
.Y(n_2482)
);

NAND3xp33_ASAP7_75t_L g2483 ( 
.A(n_2341),
.B(n_2203),
.C(n_2191),
.Y(n_2483)
);

AOI22xp33_ASAP7_75t_L g2484 ( 
.A1(n_2255),
.A2(n_2161),
.B1(n_2197),
.B2(n_2191),
.Y(n_2484)
);

OR2x2_ASAP7_75t_L g2485 ( 
.A(n_2270),
.B(n_2164),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2368),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2305),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2315),
.B(n_2354),
.Y(n_2488)
);

INVx2_ASAP7_75t_SL g2489 ( 
.A(n_2403),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2289),
.Y(n_2490)
);

BUFx3_ASAP7_75t_L g2491 ( 
.A(n_2403),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2290),
.Y(n_2492)
);

AOI22xp33_ASAP7_75t_SL g2493 ( 
.A1(n_2333),
.A2(n_2279),
.B1(n_2345),
.B2(n_2319),
.Y(n_2493)
);

AOI22xp33_ASAP7_75t_L g2494 ( 
.A1(n_2300),
.A2(n_2161),
.B1(n_2197),
.B2(n_2191),
.Y(n_2494)
);

AND2x2_ASAP7_75t_L g2495 ( 
.A(n_2337),
.B(n_2197),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2336),
.B(n_2258),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2296),
.Y(n_2497)
);

BUFx2_ASAP7_75t_L g2498 ( 
.A(n_2351),
.Y(n_2498)
);

HB1xp67_ASAP7_75t_L g2499 ( 
.A(n_2338),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2297),
.Y(n_2500)
);

AND2x2_ASAP7_75t_L g2501 ( 
.A(n_2261),
.B(n_2164),
.Y(n_2501)
);

BUFx6f_ASAP7_75t_L g2502 ( 
.A(n_2260),
.Y(n_2502)
);

HB1xp67_ASAP7_75t_L g2503 ( 
.A(n_2349),
.Y(n_2503)
);

BUFx3_ASAP7_75t_L g2504 ( 
.A(n_2339),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2312),
.Y(n_2505)
);

HB1xp67_ASAP7_75t_L g2506 ( 
.A(n_2349),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2335),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2353),
.B(n_2076),
.Y(n_2508)
);

HB1xp67_ASAP7_75t_L g2509 ( 
.A(n_2359),
.Y(n_2509)
);

AOI22xp33_ASAP7_75t_L g2510 ( 
.A1(n_2300),
.A2(n_2249),
.B1(n_2241),
.B2(n_2314),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2316),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2317),
.Y(n_2512)
);

CKINVDCx11_ASAP7_75t_R g2513 ( 
.A(n_2310),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_2405),
.B(n_2047),
.Y(n_2514)
);

OR2x2_ASAP7_75t_L g2515 ( 
.A(n_2308),
.B(n_2128),
.Y(n_2515)
);

AND4x1_ASAP7_75t_L g2516 ( 
.A(n_2281),
.B(n_2235),
.C(n_2224),
.D(n_2106),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2322),
.Y(n_2517)
);

AND2x2_ASAP7_75t_L g2518 ( 
.A(n_2323),
.B(n_2076),
.Y(n_2518)
);

AOI222xp33_ASAP7_75t_L g2519 ( 
.A1(n_2292),
.A2(n_2158),
.B1(n_2156),
.B2(n_2157),
.C1(n_2201),
.C2(n_2186),
.Y(n_2519)
);

AOI22xp33_ASAP7_75t_SL g2520 ( 
.A1(n_2345),
.A2(n_2023),
.B1(n_2025),
.B2(n_2009),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2324),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2325),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2399),
.B(n_2268),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2329),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2366),
.B(n_2198),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2356),
.B(n_2201),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2340),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2387),
.B(n_2198),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2272),
.B(n_2397),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2343),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2344),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2346),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2379),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2320),
.B(n_2076),
.Y(n_2534)
);

NOR2x1_ASAP7_75t_SL g2535 ( 
.A(n_2370),
.B(n_2238),
.Y(n_2535)
);

OR2x2_ASAP7_75t_L g2536 ( 
.A(n_2318),
.B(n_2311),
.Y(n_2536)
);

OAI21xp5_ASAP7_75t_SL g2537 ( 
.A1(n_2271),
.A2(n_2238),
.B(n_2117),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2350),
.B(n_2186),
.Y(n_2538)
);

AOI22xp33_ASAP7_75t_SL g2539 ( 
.A1(n_2319),
.A2(n_2025),
.B1(n_2009),
.B2(n_2023),
.Y(n_2539)
);

INVx1_ASAP7_75t_SL g2540 ( 
.A(n_2310),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2369),
.Y(n_2541)
);

OR2x2_ASAP7_75t_SL g2542 ( 
.A(n_2394),
.B(n_2025),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2371),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2488),
.B(n_2331),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2426),
.B(n_2396),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2463),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2417),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2421),
.B(n_2321),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2429),
.Y(n_2549)
);

INVx2_ASAP7_75t_SL g2550 ( 
.A(n_2435),
.Y(n_2550)
);

HB1xp67_ASAP7_75t_L g2551 ( 
.A(n_2499),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2437),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2444),
.Y(n_2553)
);

OAI21xp33_ASAP7_75t_L g2554 ( 
.A1(n_2473),
.A2(n_2493),
.B(n_2469),
.Y(n_2554)
);

NOR2xp67_ASAP7_75t_L g2555 ( 
.A(n_2529),
.B(n_2409),
.Y(n_2555)
);

INVx3_ASAP7_75t_L g2556 ( 
.A(n_2481),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2446),
.Y(n_2557)
);

AND2x2_ASAP7_75t_L g2558 ( 
.A(n_2416),
.B(n_2401),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2486),
.Y(n_2559)
);

BUFx2_ASAP7_75t_L g2560 ( 
.A(n_2419),
.Y(n_2560)
);

AND2x2_ASAP7_75t_L g2561 ( 
.A(n_2496),
.B(n_2401),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2487),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2447),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2477),
.B(n_2321),
.Y(n_2564)
);

INVx1_ASAP7_75t_SL g2565 ( 
.A(n_2513),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2471),
.B(n_2326),
.Y(n_2566)
);

OAI22xp5_ASAP7_75t_L g2567 ( 
.A1(n_2493),
.A2(n_2271),
.B1(n_2363),
.B2(n_2394),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2451),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2461),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2433),
.B(n_2326),
.Y(n_2570)
);

CKINVDCx5p33_ASAP7_75t_R g2571 ( 
.A(n_2513),
.Y(n_2571)
);

INVx3_ASAP7_75t_L g2572 ( 
.A(n_2481),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2490),
.B(n_2332),
.Y(n_2573)
);

INVxp67_ASAP7_75t_SL g2574 ( 
.A(n_2499),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2465),
.Y(n_2575)
);

OR2x2_ASAP7_75t_L g2576 ( 
.A(n_2455),
.B(n_2332),
.Y(n_2576)
);

AND2x4_ASAP7_75t_L g2577 ( 
.A(n_2525),
.B(n_2528),
.Y(n_2577)
);

AND2x2_ASAP7_75t_L g2578 ( 
.A(n_2432),
.B(n_2350),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2466),
.Y(n_2579)
);

AND2x4_ASAP7_75t_L g2580 ( 
.A(n_2495),
.B(n_2383),
.Y(n_2580)
);

AOI22xp33_ASAP7_75t_L g2581 ( 
.A1(n_2510),
.A2(n_2283),
.B1(n_2391),
.B2(n_2348),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2467),
.Y(n_2582)
);

BUFx2_ASAP7_75t_L g2583 ( 
.A(n_2419),
.Y(n_2583)
);

AND2x2_ASAP7_75t_L g2584 ( 
.A(n_2415),
.B(n_2372),
.Y(n_2584)
);

INVx2_ASAP7_75t_SL g2585 ( 
.A(n_2435),
.Y(n_2585)
);

AND2x2_ASAP7_75t_L g2586 ( 
.A(n_2441),
.B(n_2373),
.Y(n_2586)
);

HB1xp67_ASAP7_75t_L g2587 ( 
.A(n_2503),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2470),
.Y(n_2588)
);

INVxp67_ASAP7_75t_L g2589 ( 
.A(n_2422),
.Y(n_2589)
);

BUFx6f_ASAP7_75t_L g2590 ( 
.A(n_2502),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2507),
.Y(n_2591)
);

AOI22xp33_ASAP7_75t_L g2592 ( 
.A1(n_2510),
.A2(n_2391),
.B1(n_2348),
.B2(n_2380),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2475),
.B(n_2382),
.Y(n_2593)
);

OR2x2_ASAP7_75t_L g2594 ( 
.A(n_2422),
.B(n_2306),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2492),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2497),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_2427),
.B(n_2478),
.Y(n_2597)
);

BUFx2_ASAP7_75t_L g2598 ( 
.A(n_2491),
.Y(n_2598)
);

BUFx3_ASAP7_75t_L g2599 ( 
.A(n_2424),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2500),
.B(n_2382),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2505),
.Y(n_2601)
);

NAND2xp33_ASAP7_75t_SL g2602 ( 
.A(n_2498),
.B(n_2302),
.Y(n_2602)
);

HB1xp67_ASAP7_75t_L g2603 ( 
.A(n_2506),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2450),
.B(n_2408),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2533),
.Y(n_2605)
);

OR2x2_ASAP7_75t_L g2606 ( 
.A(n_2423),
.B(n_2306),
.Y(n_2606)
);

AOI21xp5_ASAP7_75t_R g2607 ( 
.A1(n_2445),
.A2(n_2398),
.B(n_2380),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2541),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2543),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2515),
.B(n_2375),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2480),
.B(n_2378),
.Y(n_2611)
);

AND2x4_ASAP7_75t_L g2612 ( 
.A(n_2457),
.B(n_2384),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2423),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2456),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2514),
.B(n_2275),
.Y(n_2615)
);

AND2x2_ASAP7_75t_L g2616 ( 
.A(n_2464),
.B(n_2295),
.Y(n_2616)
);

BUFx8_ASAP7_75t_L g2617 ( 
.A(n_2489),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2442),
.B(n_2313),
.Y(n_2618)
);

AOI222xp33_ASAP7_75t_L g2619 ( 
.A1(n_2424),
.A2(n_2281),
.B1(n_2244),
.B2(n_2398),
.C1(n_2411),
.C2(n_2410),
.Y(n_2619)
);

AND2x2_ASAP7_75t_L g2620 ( 
.A(n_2453),
.B(n_2458),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2468),
.Y(n_2621)
);

AOI22xp33_ASAP7_75t_L g2622 ( 
.A1(n_2430),
.A2(n_2348),
.B1(n_2342),
.B2(n_2411),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2511),
.Y(n_2623)
);

AND2x2_ASAP7_75t_L g2624 ( 
.A(n_2489),
.B(n_2400),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2512),
.Y(n_2625)
);

INVx3_ASAP7_75t_L g2626 ( 
.A(n_2481),
.Y(n_2626)
);

OAI22xp5_ASAP7_75t_L g2627 ( 
.A1(n_2439),
.A2(n_2342),
.B1(n_2355),
.B2(n_2339),
.Y(n_2627)
);

NAND2xp33_ASAP7_75t_R g2628 ( 
.A(n_2452),
.B(n_2351),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2436),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2438),
.Y(n_2630)
);

INVx4_ASAP7_75t_L g2631 ( 
.A(n_2504),
.Y(n_2631)
);

INVxp67_ASAP7_75t_SL g2632 ( 
.A(n_2509),
.Y(n_2632)
);

NOR2x1_ASAP7_75t_L g2633 ( 
.A(n_2504),
.B(n_2491),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2517),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2521),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2438),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2522),
.B(n_2406),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2523),
.B(n_2407),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2443),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2524),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_L g2641 ( 
.A(n_2516),
.B(n_2358),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2443),
.Y(n_2642)
);

AND2x4_ASAP7_75t_L g2643 ( 
.A(n_2538),
.B(n_2389),
.Y(n_2643)
);

INVx3_ASAP7_75t_L g2644 ( 
.A(n_2556),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2546),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2620),
.B(n_2474),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2545),
.B(n_2449),
.Y(n_2647)
);

NAND4xp25_ASAP7_75t_L g2648 ( 
.A(n_2554),
.B(n_2469),
.C(n_2540),
.D(n_2484),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2620),
.B(n_2474),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2560),
.B(n_2418),
.Y(n_2650)
);

HB1xp67_ASAP7_75t_L g2651 ( 
.A(n_2583),
.Y(n_2651)
);

AND2x4_ASAP7_75t_L g2652 ( 
.A(n_2556),
.B(n_2572),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2561),
.B(n_2448),
.Y(n_2653)
);

NOR2xp67_ASAP7_75t_L g2654 ( 
.A(n_2631),
.B(n_2555),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2577),
.B(n_2508),
.Y(n_2655)
);

AND2x2_ASAP7_75t_L g2656 ( 
.A(n_2577),
.B(n_2580),
.Y(n_2656)
);

AND2x4_ASAP7_75t_L g2657 ( 
.A(n_2556),
.B(n_2483),
.Y(n_2657)
);

AND2x2_ASAP7_75t_L g2658 ( 
.A(n_2577),
.B(n_2508),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2580),
.B(n_2420),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2580),
.B(n_2420),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2643),
.B(n_2431),
.Y(n_2661)
);

NOR2xp33_ASAP7_75t_L g2662 ( 
.A(n_2565),
.B(n_2395),
.Y(n_2662)
);

OR2x2_ASAP7_75t_L g2663 ( 
.A(n_2593),
.B(n_2485),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2643),
.B(n_2431),
.Y(n_2664)
);

AND2x2_ASAP7_75t_L g2665 ( 
.A(n_2643),
.B(n_2518),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2605),
.B(n_2527),
.Y(n_2666)
);

AND2x4_ASAP7_75t_L g2667 ( 
.A(n_2572),
.B(n_2626),
.Y(n_2667)
);

INVxp67_ASAP7_75t_SL g2668 ( 
.A(n_2551),
.Y(n_2668)
);

AND2x2_ASAP7_75t_L g2669 ( 
.A(n_2612),
.B(n_2518),
.Y(n_2669)
);

INVxp67_ASAP7_75t_L g2670 ( 
.A(n_2598),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2600),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2612),
.B(n_2501),
.Y(n_2672)
);

NOR2xp33_ASAP7_75t_R g2673 ( 
.A(n_2617),
.B(n_2273),
.Y(n_2673)
);

OR2x6_ASAP7_75t_L g2674 ( 
.A(n_2594),
.B(n_2537),
.Y(n_2674)
);

OR2x2_ASAP7_75t_L g2675 ( 
.A(n_2576),
.B(n_2459),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2623),
.Y(n_2676)
);

AND2x4_ASAP7_75t_SL g2677 ( 
.A(n_2631),
.B(n_2452),
.Y(n_2677)
);

HB1xp67_ASAP7_75t_L g2678 ( 
.A(n_2551),
.Y(n_2678)
);

HB1xp67_ASAP7_75t_L g2679 ( 
.A(n_2587),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2615),
.B(n_2534),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2625),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2613),
.B(n_2530),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2614),
.B(n_2531),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2621),
.B(n_2532),
.Y(n_2684)
);

AND2x2_ASAP7_75t_L g2685 ( 
.A(n_2626),
.B(n_2539),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2626),
.B(n_2539),
.Y(n_2686)
);

INVx3_ASAP7_75t_L g2687 ( 
.A(n_2590),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2547),
.B(n_2549),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2634),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2635),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2640),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2552),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2676),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2676),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2681),
.Y(n_2695)
);

NAND2x1_ASAP7_75t_L g2696 ( 
.A(n_2654),
.B(n_2631),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2661),
.B(n_2664),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2681),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2661),
.B(n_2520),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2689),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2689),
.Y(n_2701)
);

NOR2xp67_ASAP7_75t_L g2702 ( 
.A(n_2654),
.B(n_2571),
.Y(n_2702)
);

AND2x2_ASAP7_75t_L g2703 ( 
.A(n_2664),
.B(n_2520),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2690),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2646),
.B(n_2604),
.Y(n_2705)
);

INVx1_ASAP7_75t_SL g2706 ( 
.A(n_2673),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2690),
.Y(n_2707)
);

OR2x2_ASAP7_75t_L g2708 ( 
.A(n_2663),
.B(n_2606),
.Y(n_2708)
);

AND2x2_ASAP7_75t_L g2709 ( 
.A(n_2646),
.B(n_2629),
.Y(n_2709)
);

HB1xp67_ASAP7_75t_L g2710 ( 
.A(n_2678),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2691),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2649),
.B(n_2630),
.Y(n_2712)
);

OR2x2_ASAP7_75t_L g2713 ( 
.A(n_2663),
.B(n_2675),
.Y(n_2713)
);

AND2x4_ASAP7_75t_SL g2714 ( 
.A(n_2656),
.B(n_2550),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_SL g2715 ( 
.A(n_2677),
.B(n_2567),
.Y(n_2715)
);

OAI21xp33_ASAP7_75t_SL g2716 ( 
.A1(n_2656),
.A2(n_2619),
.B(n_2585),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2649),
.B(n_2630),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2665),
.B(n_2636),
.Y(n_2718)
);

OR2x2_ASAP7_75t_L g2719 ( 
.A(n_2675),
.B(n_2589),
.Y(n_2719)
);

NOR3x1_ASAP7_75t_L g2720 ( 
.A(n_2648),
.B(n_2585),
.C(n_2550),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2691),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2671),
.B(n_2589),
.Y(n_2722)
);

AOI21x1_ASAP7_75t_SL g2723 ( 
.A1(n_2651),
.A2(n_2607),
.B(n_2462),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2692),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2692),
.Y(n_2725)
);

AND2x2_ASAP7_75t_L g2726 ( 
.A(n_2665),
.B(n_2636),
.Y(n_2726)
);

OR2x2_ASAP7_75t_L g2727 ( 
.A(n_2650),
.B(n_2587),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2655),
.B(n_2658),
.Y(n_2728)
);

INVx1_ASAP7_75t_SL g2729 ( 
.A(n_2677),
.Y(n_2729)
);

INVx2_ASAP7_75t_SL g2730 ( 
.A(n_2677),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2655),
.B(n_2639),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2645),
.Y(n_2732)
);

NOR2xp33_ASAP7_75t_L g2733 ( 
.A(n_2662),
.B(n_2571),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2645),
.Y(n_2734)
);

AND2x2_ASAP7_75t_L g2735 ( 
.A(n_2658),
.B(n_2639),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2659),
.B(n_2642),
.Y(n_2736)
);

AND2x2_ASAP7_75t_L g2737 ( 
.A(n_2659),
.B(n_2642),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2671),
.B(n_2553),
.Y(n_2738)
);

HB1xp67_ASAP7_75t_L g2739 ( 
.A(n_2679),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2713),
.Y(n_2740)
);

INVxp67_ASAP7_75t_L g2741 ( 
.A(n_2710),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2713),
.Y(n_2742)
);

OR2x2_ASAP7_75t_L g2743 ( 
.A(n_2708),
.B(n_2647),
.Y(n_2743)
);

HB1xp67_ASAP7_75t_L g2744 ( 
.A(n_2739),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2719),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2705),
.B(n_2668),
.Y(n_2746)
);

HB1xp67_ASAP7_75t_L g2747 ( 
.A(n_2727),
.Y(n_2747)
);

BUFx3_ASAP7_75t_L g2748 ( 
.A(n_2696),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2719),
.Y(n_2749)
);

OR2x2_ASAP7_75t_L g2750 ( 
.A(n_2708),
.B(n_2653),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2727),
.Y(n_2751)
);

OR2x2_ASAP7_75t_L g2752 ( 
.A(n_2709),
.B(n_2660),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2738),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2705),
.B(n_2648),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2693),
.Y(n_2755)
);

OAI21xp5_ASAP7_75t_L g2756 ( 
.A1(n_2716),
.A2(n_2627),
.B(n_2670),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2693),
.Y(n_2757)
);

OR2x2_ASAP7_75t_L g2758 ( 
.A(n_2709),
.B(n_2660),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2704),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2732),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2699),
.B(n_2680),
.Y(n_2761)
);

INVx2_ASAP7_75t_SL g2762 ( 
.A(n_2696),
.Y(n_2762)
);

INVx1_ASAP7_75t_SL g2763 ( 
.A(n_2706),
.Y(n_2763)
);

AND2x2_ASAP7_75t_L g2764 ( 
.A(n_2728),
.B(n_2669),
.Y(n_2764)
);

OAI21xp33_ASAP7_75t_L g2765 ( 
.A1(n_2715),
.A2(n_2581),
.B(n_2685),
.Y(n_2765)
);

OR2x2_ASAP7_75t_L g2766 ( 
.A(n_2712),
.B(n_2680),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2728),
.B(n_2669),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2697),
.B(n_2685),
.Y(n_2768)
);

OAI21xp5_ASAP7_75t_L g2769 ( 
.A1(n_2702),
.A2(n_2581),
.B(n_2622),
.Y(n_2769)
);

INVx2_ASAP7_75t_SL g2770 ( 
.A(n_2714),
.Y(n_2770)
);

INVx3_ASAP7_75t_L g2771 ( 
.A(n_2730),
.Y(n_2771)
);

OR2x2_ASAP7_75t_L g2772 ( 
.A(n_2712),
.B(n_2717),
.Y(n_2772)
);

INVx1_ASAP7_75t_SL g2773 ( 
.A(n_2714),
.Y(n_2773)
);

INVxp67_ASAP7_75t_SL g2774 ( 
.A(n_2720),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2704),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2707),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2732),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2707),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2699),
.B(n_2686),
.Y(n_2779)
);

OAI21xp5_ASAP7_75t_L g2780 ( 
.A1(n_2730),
.A2(n_2622),
.B(n_2592),
.Y(n_2780)
);

OAI32xp33_ASAP7_75t_L g2781 ( 
.A1(n_2729),
.A2(n_2599),
.A3(n_2602),
.B1(n_2628),
.B2(n_2644),
.Y(n_2781)
);

AOI22xp5_ASAP7_75t_L g2782 ( 
.A1(n_2703),
.A2(n_2592),
.B1(n_2674),
.B2(n_2686),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2703),
.B(n_2672),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2747),
.Y(n_2784)
);

AOI21xp33_ASAP7_75t_L g2785 ( 
.A1(n_2774),
.A2(n_2641),
.B(n_2733),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2747),
.Y(n_2786)
);

AOI22xp5_ASAP7_75t_L g2787 ( 
.A1(n_2765),
.A2(n_2674),
.B1(n_2722),
.B2(n_2697),
.Y(n_2787)
);

OAI21xp5_ASAP7_75t_L g2788 ( 
.A1(n_2756),
.A2(n_2774),
.B(n_2769),
.Y(n_2788)
);

OAI32xp33_ASAP7_75t_L g2789 ( 
.A1(n_2773),
.A2(n_2599),
.A3(n_2602),
.B1(n_2628),
.B2(n_2641),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2771),
.B(n_2731),
.Y(n_2790)
);

OAI32xp33_ASAP7_75t_L g2791 ( 
.A1(n_2771),
.A2(n_2754),
.A3(n_2770),
.B1(n_2748),
.B2(n_2763),
.Y(n_2791)
);

O2A1O1Ixp33_ASAP7_75t_L g2792 ( 
.A1(n_2762),
.A2(n_2402),
.B(n_2273),
.C(n_2294),
.Y(n_2792)
);

OAI22xp5_ASAP7_75t_L g2793 ( 
.A1(n_2770),
.A2(n_2674),
.B1(n_2542),
.B2(n_2633),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2744),
.B(n_2717),
.Y(n_2794)
);

O2A1O1Ixp33_ASAP7_75t_L g2795 ( 
.A1(n_2762),
.A2(n_2294),
.B(n_2425),
.C(n_2674),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2744),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2755),
.Y(n_2797)
);

NOR2xp33_ASAP7_75t_L g2798 ( 
.A(n_2753),
.B(n_2282),
.Y(n_2798)
);

O2A1O1Ixp33_ASAP7_75t_L g2799 ( 
.A1(n_2780),
.A2(n_2425),
.B(n_2674),
.C(n_2476),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2757),
.Y(n_2800)
);

OAI32xp33_ASAP7_75t_L g2801 ( 
.A1(n_2771),
.A2(n_2644),
.A3(n_2536),
.B1(n_2302),
.B2(n_2694),
.Y(n_2801)
);

AO221x1_ASAP7_75t_L g2802 ( 
.A1(n_2741),
.A2(n_2644),
.B1(n_2452),
.B2(n_2723),
.C(n_2617),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2759),
.Y(n_2803)
);

AOI22xp5_ASAP7_75t_L g2804 ( 
.A1(n_2782),
.A2(n_2638),
.B1(n_2737),
.B2(n_2736),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_SL g2805 ( 
.A(n_2748),
.B(n_2617),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2775),
.Y(n_2806)
);

AOI22xp5_ASAP7_75t_L g2807 ( 
.A1(n_2745),
.A2(n_2737),
.B1(n_2736),
.B2(n_2726),
.Y(n_2807)
);

O2A1O1Ixp5_ASAP7_75t_L g2808 ( 
.A1(n_2781),
.A2(n_2695),
.B(n_2700),
.C(n_2698),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2772),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2796),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_SL g2811 ( 
.A(n_2792),
.B(n_2741),
.Y(n_2811)
);

NAND2x1_ASAP7_75t_SL g2812 ( 
.A(n_2787),
.B(n_2768),
.Y(n_2812)
);

OAI21xp33_ASAP7_75t_L g2813 ( 
.A1(n_2788),
.A2(n_2779),
.B(n_2751),
.Y(n_2813)
);

AOI21xp33_ASAP7_75t_L g2814 ( 
.A1(n_2792),
.A2(n_2564),
.B(n_2548),
.Y(n_2814)
);

AOI21xp33_ASAP7_75t_SL g2815 ( 
.A1(n_2791),
.A2(n_2749),
.B(n_2742),
.Y(n_2815)
);

AOI21xp5_ASAP7_75t_L g2816 ( 
.A1(n_2795),
.A2(n_2746),
.B(n_2740),
.Y(n_2816)
);

OAI22xp5_ASAP7_75t_L g2817 ( 
.A1(n_2795),
.A2(n_2750),
.B1(n_2766),
.B2(n_2743),
.Y(n_2817)
);

OAI211xp5_ASAP7_75t_SL g2818 ( 
.A1(n_2785),
.A2(n_2434),
.B(n_2783),
.C(n_2519),
.Y(n_2818)
);

XOR2x2_ASAP7_75t_L g2819 ( 
.A(n_2798),
.B(n_2805),
.Y(n_2819)
);

AOI22xp5_ASAP7_75t_L g2820 ( 
.A1(n_2793),
.A2(n_2768),
.B1(n_2761),
.B2(n_2652),
.Y(n_2820)
);

OAI221xp5_ASAP7_75t_L g2821 ( 
.A1(n_2808),
.A2(n_2434),
.B1(n_2778),
.B2(n_2776),
.C(n_2404),
.Y(n_2821)
);

AOI22xp5_ASAP7_75t_L g2822 ( 
.A1(n_2804),
.A2(n_2667),
.B1(n_2652),
.B2(n_2657),
.Y(n_2822)
);

O2A1O1Ixp33_ASAP7_75t_L g2823 ( 
.A1(n_2799),
.A2(n_2789),
.B(n_2801),
.C(n_2786),
.Y(n_2823)
);

AOI21xp5_ASAP7_75t_L g2824 ( 
.A1(n_2802),
.A2(n_2535),
.B(n_2688),
.Y(n_2824)
);

OAI22xp5_ASAP7_75t_L g2825 ( 
.A1(n_2807),
.A2(n_2758),
.B1(n_2752),
.B2(n_2764),
.Y(n_2825)
);

OAI322xp33_ASAP7_75t_L g2826 ( 
.A1(n_2784),
.A2(n_2711),
.A3(n_2721),
.B1(n_2724),
.B2(n_2725),
.C1(n_2701),
.C2(n_2666),
.Y(n_2826)
);

NAND2xp33_ASAP7_75t_L g2827 ( 
.A(n_2794),
.B(n_2767),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2809),
.Y(n_2828)
);

AOI21xp33_ASAP7_75t_L g2829 ( 
.A1(n_2799),
.A2(n_2683),
.B(n_2682),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2797),
.Y(n_2830)
);

OAI22xp5_ASAP7_75t_L g2831 ( 
.A1(n_2790),
.A2(n_2726),
.B1(n_2718),
.B2(n_2731),
.Y(n_2831)
);

AOI21xp33_ASAP7_75t_L g2832 ( 
.A1(n_2800),
.A2(n_2684),
.B(n_2414),
.Y(n_2832)
);

AOI311xp33_ASAP7_75t_L g2833 ( 
.A1(n_2803),
.A2(n_2568),
.A3(n_2601),
.B(n_2596),
.C(n_2595),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2806),
.B(n_2760),
.Y(n_2834)
);

OAI21xp33_ASAP7_75t_L g2835 ( 
.A1(n_2788),
.A2(n_2777),
.B(n_2760),
.Y(n_2835)
);

NAND4xp25_ASAP7_75t_L g2836 ( 
.A(n_2788),
.B(n_2404),
.C(n_2484),
.D(n_2428),
.Y(n_2836)
);

A2O1A1Ixp33_ASAP7_75t_L g2837 ( 
.A1(n_2792),
.A2(n_2718),
.B(n_2735),
.C(n_2652),
.Y(n_2837)
);

NOR3xp33_ASAP7_75t_L g2838 ( 
.A(n_2823),
.B(n_2374),
.C(n_2330),
.Y(n_2838)
);

NOR2x1_ASAP7_75t_L g2839 ( 
.A(n_2811),
.B(n_2374),
.Y(n_2839)
);

NAND4xp25_ASAP7_75t_L g2840 ( 
.A(n_2818),
.B(n_2813),
.C(n_2815),
.D(n_2821),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2830),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2816),
.B(n_2777),
.Y(n_2842)
);

NOR2xp33_ASAP7_75t_L g2843 ( 
.A(n_2817),
.B(n_2288),
.Y(n_2843)
);

OA22x2_ASAP7_75t_L g2844 ( 
.A1(n_2835),
.A2(n_2611),
.B1(n_2657),
.B2(n_2652),
.Y(n_2844)
);

AOI221xp5_ASAP7_75t_L g2845 ( 
.A1(n_2817),
.A2(n_2575),
.B1(n_2591),
.B2(n_2557),
.C(n_2559),
.Y(n_2845)
);

NOR2xp33_ASAP7_75t_SL g2846 ( 
.A(n_2824),
.B(n_2282),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2829),
.B(n_2735),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_SL g2848 ( 
.A(n_2833),
.B(n_2657),
.Y(n_2848)
);

NAND3xp33_ASAP7_75t_L g2849 ( 
.A(n_2810),
.B(n_2428),
.C(n_2494),
.Y(n_2849)
);

AOI21xp5_ASAP7_75t_L g2850 ( 
.A1(n_2819),
.A2(n_2632),
.B(n_2574),
.Y(n_2850)
);

NOR2xp33_ASAP7_75t_L g2851 ( 
.A(n_2826),
.B(n_2288),
.Y(n_2851)
);

NOR2xp33_ASAP7_75t_L g2852 ( 
.A(n_2825),
.B(n_2301),
.Y(n_2852)
);

AOI21xp5_ASAP7_75t_L g2853 ( 
.A1(n_2837),
.A2(n_2827),
.B(n_2834),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_SL g2854 ( 
.A(n_2820),
.B(n_2657),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2828),
.B(n_2597),
.Y(n_2855)
);

INVxp33_ASAP7_75t_SL g2856 ( 
.A(n_2822),
.Y(n_2856)
);

NAND4xp25_ASAP7_75t_L g2857 ( 
.A(n_2836),
.B(n_2494),
.C(n_2440),
.D(n_2482),
.Y(n_2857)
);

AND2x2_ASAP7_75t_L g2858 ( 
.A(n_2831),
.B(n_2672),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2845),
.B(n_2814),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2851),
.B(n_2847),
.Y(n_2860)
);

AOI22xp5_ASAP7_75t_L g2861 ( 
.A1(n_2840),
.A2(n_2832),
.B1(n_2616),
.B2(n_2578),
.Y(n_2861)
);

NOR2xp33_ASAP7_75t_L g2862 ( 
.A(n_2843),
.B(n_2812),
.Y(n_2862)
);

NOR2xp33_ASAP7_75t_L g2863 ( 
.A(n_2856),
.B(n_2852),
.Y(n_2863)
);

NAND3xp33_ASAP7_75t_L g2864 ( 
.A(n_2838),
.B(n_2413),
.C(n_2734),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_SL g2865 ( 
.A(n_2846),
.B(n_2309),
.Y(n_2865)
);

NOR2x1_ASAP7_75t_L g2866 ( 
.A(n_2839),
.B(n_2364),
.Y(n_2866)
);

NOR4xp25_ASAP7_75t_L g2867 ( 
.A(n_2841),
.B(n_2848),
.C(n_2857),
.D(n_2842),
.Y(n_2867)
);

NOR2x1_ASAP7_75t_L g2868 ( 
.A(n_2850),
.B(n_2364),
.Y(n_2868)
);

NOR2xp67_ASAP7_75t_SL g2869 ( 
.A(n_2853),
.B(n_2388),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2855),
.Y(n_2870)
);

NAND3xp33_ASAP7_75t_L g2871 ( 
.A(n_2849),
.B(n_2734),
.C(n_2563),
.Y(n_2871)
);

AOI22xp5_ASAP7_75t_L g2872 ( 
.A1(n_2854),
.A2(n_2667),
.B1(n_2644),
.B2(n_2624),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2858),
.B(n_2562),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2844),
.B(n_2569),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2844),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2870),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2873),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2859),
.B(n_2579),
.Y(n_2878)
);

NAND3xp33_ASAP7_75t_SL g2879 ( 
.A(n_2867),
.B(n_2355),
.C(n_2412),
.Y(n_2879)
);

NOR2xp67_ASAP7_75t_SL g2880 ( 
.A(n_2865),
.B(n_2440),
.Y(n_2880)
);

NAND4xp75_ASAP7_75t_L g2881 ( 
.A(n_2875),
.B(n_2472),
.C(n_2479),
.D(n_2544),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2861),
.Y(n_2882)
);

NAND4xp75_ASAP7_75t_L g2883 ( 
.A(n_2863),
.B(n_2862),
.C(n_2868),
.D(n_2860),
.Y(n_2883)
);

NAND4xp75_ASAP7_75t_L g2884 ( 
.A(n_2866),
.B(n_2472),
.C(n_2526),
.D(n_2586),
.Y(n_2884)
);

NOR4xp75_ASAP7_75t_L g2885 ( 
.A(n_2874),
.B(n_2388),
.C(n_2377),
.D(n_2330),
.Y(n_2885)
);

NOR2x1_ASAP7_75t_L g2886 ( 
.A(n_2871),
.B(n_2454),
.Y(n_2886)
);

NOR3xp33_ASAP7_75t_L g2887 ( 
.A(n_2864),
.B(n_2377),
.C(n_2566),
.Y(n_2887)
);

NOR2x1_ASAP7_75t_L g2888 ( 
.A(n_2869),
.B(n_2454),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2872),
.Y(n_2889)
);

NOR2x1_ASAP7_75t_L g2890 ( 
.A(n_2863),
.B(n_2482),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2876),
.Y(n_2891)
);

AO22x1_ASAP7_75t_L g2892 ( 
.A1(n_2890),
.A2(n_2582),
.B1(n_2588),
.B2(n_2608),
.Y(n_2892)
);

AOI22xp5_ASAP7_75t_L g2893 ( 
.A1(n_2879),
.A2(n_2667),
.B1(n_2618),
.B2(n_2609),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2877),
.Y(n_2894)
);

INVx1_ASAP7_75t_SL g2895 ( 
.A(n_2883),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2878),
.Y(n_2896)
);

NOR2x1_ASAP7_75t_L g2897 ( 
.A(n_2882),
.B(n_2385),
.Y(n_2897)
);

HB1xp67_ASAP7_75t_L g2898 ( 
.A(n_2889),
.Y(n_2898)
);

NOR2x1_ASAP7_75t_L g2899 ( 
.A(n_2888),
.B(n_2385),
.Y(n_2899)
);

NAND2x1p5_ASAP7_75t_SL g2900 ( 
.A(n_2886),
.B(n_2570),
.Y(n_2900)
);

NOR2xp67_ASAP7_75t_L g2901 ( 
.A(n_2878),
.B(n_2687),
.Y(n_2901)
);

AND2x2_ASAP7_75t_L g2902 ( 
.A(n_2880),
.B(n_2667),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2898),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2891),
.Y(n_2904)
);

AOI22xp5_ASAP7_75t_L g2905 ( 
.A1(n_2895),
.A2(n_2884),
.B1(n_2881),
.B2(n_2887),
.Y(n_2905)
);

AOI22xp5_ASAP7_75t_L g2906 ( 
.A1(n_2897),
.A2(n_2885),
.B1(n_2584),
.B2(n_2298),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2894),
.Y(n_2907)
);

INVx2_ASAP7_75t_SL g2908 ( 
.A(n_2902),
.Y(n_2908)
);

INVx2_ASAP7_75t_SL g2909 ( 
.A(n_2899),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2896),
.Y(n_2910)
);

CKINVDCx5p33_ASAP7_75t_R g2911 ( 
.A(n_2892),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2901),
.Y(n_2912)
);

AOI22x1_ASAP7_75t_L g2913 ( 
.A1(n_2900),
.A2(n_2901),
.B1(n_2893),
.B2(n_2603),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2898),
.Y(n_2914)
);

XNOR2x1_ASAP7_75t_L g2915 ( 
.A(n_2895),
.B(n_2445),
.Y(n_2915)
);

AOI22xp5_ASAP7_75t_L g2916 ( 
.A1(n_2908),
.A2(n_2362),
.B1(n_2445),
.B2(n_2298),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2903),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2903),
.Y(n_2918)
);

XNOR2xp5_ASAP7_75t_L g2919 ( 
.A(n_2915),
.B(n_2905),
.Y(n_2919)
);

AOI22xp5_ASAP7_75t_L g2920 ( 
.A1(n_2914),
.A2(n_2362),
.B1(n_2298),
.B2(n_2610),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2904),
.Y(n_2921)
);

NOR2xp33_ASAP7_75t_L g2922 ( 
.A(n_2911),
.B(n_2637),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2921),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2917),
.Y(n_2924)
);

INVxp67_ASAP7_75t_SL g2925 ( 
.A(n_2918),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2919),
.Y(n_2926)
);

NOR2xp33_ASAP7_75t_L g2927 ( 
.A(n_2922),
.B(n_2907),
.Y(n_2927)
);

AOI21xp5_ASAP7_75t_L g2928 ( 
.A1(n_2925),
.A2(n_2910),
.B(n_2909),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2925),
.Y(n_2929)
);

OAI22xp5_ASAP7_75t_SL g2930 ( 
.A1(n_2926),
.A2(n_2912),
.B1(n_2920),
.B2(n_2916),
.Y(n_2930)
);

AOI22xp5_ASAP7_75t_L g2931 ( 
.A1(n_2927),
.A2(n_2906),
.B1(n_2913),
.B2(n_2362),
.Y(n_2931)
);

OAI21xp5_ASAP7_75t_L g2932 ( 
.A1(n_2923),
.A2(n_2206),
.B(n_2156),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2929),
.Y(n_2933)
);

OAI22xp5_ASAP7_75t_SL g2934 ( 
.A1(n_2930),
.A2(n_2924),
.B1(n_2385),
.B2(n_2573),
.Y(n_2934)
);

NOR3xp33_ASAP7_75t_L g2935 ( 
.A(n_2928),
.B(n_2157),
.C(n_2687),
.Y(n_2935)
);

AOI31xp33_ASAP7_75t_L g2936 ( 
.A1(n_2933),
.A2(n_2931),
.A3(n_2934),
.B(n_2932),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2936),
.B(n_2935),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2937),
.B(n_2206),
.Y(n_2938)
);

AOI22xp5_ASAP7_75t_L g2939 ( 
.A1(n_2938),
.A2(n_2460),
.B1(n_2558),
.B2(n_2687),
.Y(n_2939)
);


endmodule