module fake_netlist_6_2669_n_1072 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1072);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1072;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_1008;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_875;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_341;
wire n_362;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_544;
wire n_372;
wire n_468;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_758;
wire n_525;
wire n_720;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_723;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_189),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_120),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_108),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_188),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_213),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_95),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_187),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_13),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_55),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_138),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_147),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_8),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_242),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_208),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_203),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_103),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_173),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_247),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_215),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_198),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_47),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_230),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_71),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_127),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_36),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_72),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_231),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_52),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_206),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_245),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_60),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_130),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_182),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_177),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_248),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_57),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_186),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_93),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_100),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_226),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_44),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_162),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_167),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_222),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_78),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_53),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_70),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_212),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_228),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_204),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_122),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_59),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_104),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_13),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_134),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_64),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_45),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_110),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_98),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_202),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_154),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_168),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_29),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_80),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_161),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_252),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_265),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_261),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_278),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_307),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_270),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_293),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_256),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_256),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_306),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_268),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_260),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_284),
.B(n_0),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_268),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_276),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_291),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_255),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_294),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_297),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_274),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_306),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_254),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_300),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_257),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_312),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_255),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_312),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_259),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_255),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_255),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_262),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_263),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_315),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_264),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_266),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_315),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_267),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_315),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_315),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_L g361 ( 
.A(n_269),
.B(n_0),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_361),
.B(n_335),
.Y(n_362)
);

CKINVDCx8_ASAP7_75t_R g363 ( 
.A(n_328),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_334),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_337),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_347),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_338),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_330),
.B(n_258),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_339),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_336),
.Y(n_370)
);

AND2x4_ASAP7_75t_SL g371 ( 
.A(n_352),
.B(n_281),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_320),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_350),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_336),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_333),
.B(n_288),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_351),
.Y(n_376)
);

NAND2x1p5_ASAP7_75t_L g377 ( 
.A(n_332),
.B(n_340),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_351),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_345),
.B(n_271),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_354),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_357),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_324),
.B(n_272),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_322),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_320),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_359),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_360),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_323),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_325),
.Y(n_388)
);

INVxp33_ASAP7_75t_SL g389 ( 
.A(n_349),
.Y(n_389)
);

OAI21x1_ASAP7_75t_L g390 ( 
.A1(n_343),
.A2(n_275),
.B(n_273),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_344),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_341),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g393 ( 
.A1(n_326),
.A2(n_279),
.B(n_277),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_327),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_355),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_358),
.B(n_280),
.Y(n_397)
);

CKINVDCx8_ASAP7_75t_R g398 ( 
.A(n_328),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_355),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_349),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_353),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_329),
.A2(n_283),
.B1(n_285),
.B2(n_282),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_356),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_331),
.Y(n_405)
);

CKINVDCx6p67_ASAP7_75t_R g406 ( 
.A(n_352),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_321),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_356),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_358),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_405),
.B(n_329),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_286),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_370),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_366),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_383),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_387),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_374),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_287),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_374),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_378),
.Y(n_419)
);

NAND2xp33_ASAP7_75t_SL g420 ( 
.A(n_375),
.B(n_289),
.Y(n_420)
);

BUFx10_ASAP7_75t_L g421 ( 
.A(n_362),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_378),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_290),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_403),
.A2(n_295),
.B1(n_298),
.B2(n_292),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_370),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_399),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_370),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_388),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_364),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_373),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_370),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_370),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_365),
.Y(n_433)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

BUFx4f_ASAP7_75t_L g435 ( 
.A(n_393),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_376),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_367),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_369),
.B(n_299),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_362),
.B(n_301),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_376),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_362),
.B(n_302),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_393),
.A2(n_305),
.B1(n_308),
.B2(n_303),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_373),
.Y(n_443)
);

AO22x2_ASAP7_75t_L g444 ( 
.A1(n_409),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_380),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_371),
.B(n_342),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_L g447 ( 
.A1(n_393),
.A2(n_310),
.B1(n_311),
.B2(n_309),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_391),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_391),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_405),
.B(n_313),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_392),
.Y(n_451)
);

NAND3xp33_ASAP7_75t_L g452 ( 
.A(n_368),
.B(n_317),
.C(n_314),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_380),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_401),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_381),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_385),
.B(n_318),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_385),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_386),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_375),
.B(n_342),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_386),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_392),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_377),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_379),
.B(n_319),
.Y(n_464)
);

AND2x6_ASAP7_75t_L g465 ( 
.A(n_401),
.B(n_42),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_368),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_377),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_390),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_401),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_363),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_377),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_390),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_401),
.B(n_346),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_393),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_466),
.A2(n_389),
.B1(n_404),
.B2(n_401),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_466),
.B(n_394),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_451),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_448),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_389),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_413),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_413),
.Y(n_481)
);

AO22x2_ASAP7_75t_L g482 ( 
.A1(n_474),
.A2(n_408),
.B1(n_382),
.B2(n_397),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_436),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_426),
.B(n_408),
.Y(n_484)
);

NAND2x1p5_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_404),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_460),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_404),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_414),
.B(n_404),
.Y(n_488)
);

BUFx6f_ASAP7_75t_SL g489 ( 
.A(n_451),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_430),
.Y(n_490)
);

NAND2x1p5_ASAP7_75t_L g491 ( 
.A(n_454),
.B(n_404),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_430),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_443),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_436),
.Y(n_494)
);

AO22x2_ASAP7_75t_L g495 ( 
.A1(n_474),
.A2(n_398),
.B1(n_363),
.B2(n_348),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_443),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_445),
.Y(n_497)
);

OAI221xp5_ASAP7_75t_L g498 ( 
.A1(n_442),
.A2(n_407),
.B1(n_395),
.B2(n_384),
.C(n_372),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_470),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_445),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_458),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_458),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_461),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_464),
.B(n_400),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_461),
.Y(n_505)
);

BUFx8_ASAP7_75t_L g506 ( 
.A(n_450),
.Y(n_506)
);

OAI221xp5_ASAP7_75t_L g507 ( 
.A1(n_447),
.A2(n_407),
.B1(n_395),
.B2(n_384),
.C(n_402),
.Y(n_507)
);

NAND2x1p5_ASAP7_75t_L g508 ( 
.A(n_454),
.B(n_398),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_415),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_428),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_429),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_440),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_433),
.Y(n_513)
);

AO22x2_ASAP7_75t_L g514 ( 
.A1(n_444),
.A2(n_348),
.B1(n_346),
.B2(n_371),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_440),
.Y(n_515)
);

AO22x2_ASAP7_75t_L g516 ( 
.A1(n_444),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_437),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_450),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_423),
.Y(n_519)
);

OA22x2_ASAP7_75t_L g520 ( 
.A1(n_410),
.A2(n_406),
.B1(n_6),
.B2(n_4),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_462),
.B(n_43),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_453),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_453),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_421),
.B(n_406),
.Y(n_524)
);

OAI221xp5_ASAP7_75t_L g525 ( 
.A1(n_424),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_469),
.B(n_46),
.Y(n_526)
);

NAND3xp33_ASAP7_75t_L g527 ( 
.A(n_420),
.B(n_5),
.C(n_7),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_416),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_446),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_455),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_455),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_467),
.A2(n_49),
.B1(n_50),
.B2(n_48),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_421),
.B(n_8),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_448),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_416),
.Y(n_535)
);

AO22x2_ASAP7_75t_L g536 ( 
.A1(n_444),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_449),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_439),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_449),
.Y(n_539)
);

AO22x2_ASAP7_75t_L g540 ( 
.A1(n_444),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_540)
);

AO22x2_ASAP7_75t_L g541 ( 
.A1(n_473),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_456),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_476),
.B(n_421),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_475),
.B(n_469),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_518),
.B(n_470),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_488),
.B(n_439),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_488),
.B(n_439),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_504),
.B(n_452),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_477),
.B(n_423),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_479),
.B(n_435),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_484),
.B(n_435),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_519),
.B(n_420),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_480),
.B(n_423),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_R g554 ( 
.A(n_533),
.B(n_468),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_487),
.B(n_411),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_521),
.B(n_417),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_521),
.B(n_441),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_SL g558 ( 
.A(n_489),
.B(n_446),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_SL g559 ( 
.A(n_489),
.B(n_438),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_508),
.B(n_438),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_486),
.B(n_438),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_485),
.B(n_457),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_SL g563 ( 
.A(n_538),
.B(n_457),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_481),
.B(n_456),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_SL g565 ( 
.A(n_524),
.B(n_457),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_491),
.B(n_459),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_509),
.B(n_459),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_510),
.B(n_434),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_511),
.B(n_513),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_517),
.B(n_434),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_490),
.B(n_434),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_492),
.B(n_468),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_493),
.B(n_496),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_SL g574 ( 
.A(n_499),
.B(n_468),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_497),
.B(n_472),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_500),
.B(n_472),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_501),
.B(n_472),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_502),
.B(n_432),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_SL g579 ( 
.A(n_503),
.B(n_432),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_505),
.B(n_427),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_522),
.B(n_427),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_523),
.B(n_530),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_531),
.B(n_427),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_542),
.B(n_506),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_506),
.B(n_431),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_527),
.B(n_431),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_478),
.B(n_534),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_478),
.B(n_412),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_534),
.B(n_537),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_537),
.B(n_539),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_539),
.B(n_418),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_520),
.B(n_412),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_SL g593 ( 
.A(n_526),
.B(n_465),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_532),
.B(n_412),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_483),
.B(n_425),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_528),
.B(n_418),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_494),
.B(n_425),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_512),
.B(n_425),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_535),
.B(n_419),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_515),
.B(n_419),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_529),
.B(n_422),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_498),
.B(n_422),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_577),
.A2(n_465),
.B(n_482),
.Y(n_603)
);

AOI221xp5_ASAP7_75t_L g604 ( 
.A1(n_548),
.A2(n_507),
.B1(n_495),
.B2(n_525),
.C(n_514),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_543),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_589),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_545),
.B(n_495),
.Y(n_607)
);

NOR2xp67_ASAP7_75t_L g608 ( 
.A(n_553),
.B(n_51),
.Y(n_608)
);

AO32x2_ASAP7_75t_L g609 ( 
.A1(n_554),
.A2(n_482),
.A3(n_514),
.B1(n_536),
.B2(n_516),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_549),
.B(n_465),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_573),
.B(n_541),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_601),
.Y(n_612)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_587),
.A2(n_465),
.B(n_56),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_549),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_551),
.A2(n_541),
.B(n_536),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_589),
.Y(n_616)
);

AOI21xp33_ASAP7_75t_L g617 ( 
.A1(n_561),
.A2(n_540),
.B(n_516),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_573),
.B(n_540),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_569),
.B(n_560),
.Y(n_619)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_572),
.A2(n_58),
.B(n_54),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_557),
.B(n_12),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_SL g622 ( 
.A1(n_544),
.A2(n_62),
.B(n_61),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_584),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_564),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_552),
.B(n_14),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_L g626 ( 
.A1(n_550),
.A2(n_576),
.B(n_575),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_591),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_602),
.A2(n_253),
.B(n_63),
.Y(n_628)
);

A2O1A1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_563),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_629)
);

OAI21x1_ASAP7_75t_L g630 ( 
.A1(n_590),
.A2(n_588),
.B(n_578),
.Y(n_630)
);

O2A1O1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_546),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_547),
.A2(n_143),
.B1(n_250),
.B2(n_249),
.Y(n_632)
);

A2O1A1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_565),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_592),
.B(n_19),
.Y(n_634)
);

AO21x1_ASAP7_75t_L g635 ( 
.A1(n_593),
.A2(n_20),
.B(n_21),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_559),
.B(n_65),
.Y(n_636)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_581),
.A2(n_67),
.B(n_66),
.Y(n_637)
);

OAI21x1_ASAP7_75t_L g638 ( 
.A1(n_583),
.A2(n_566),
.B(n_580),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_585),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_L g640 ( 
.A(n_556),
.B(n_21),
.C(n_22),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_586),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_555),
.A2(n_251),
.B(n_69),
.Y(n_642)
);

AO31x2_ASAP7_75t_L g643 ( 
.A1(n_596),
.A2(n_23),
.A3(n_24),
.B(n_25),
.Y(n_643)
);

NAND2x1p5_ASAP7_75t_L g644 ( 
.A(n_562),
.B(n_68),
.Y(n_644)
);

OAI21x1_ASAP7_75t_SL g645 ( 
.A1(n_599),
.A2(n_74),
.B(n_73),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_567),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_582),
.B(n_25),
.Y(n_647)
);

OAI21x1_ASAP7_75t_L g648 ( 
.A1(n_595),
.A2(n_76),
.B(n_75),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_568),
.B(n_26),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_594),
.A2(n_151),
.B1(n_244),
.B2(n_243),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_600),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_571),
.A2(n_79),
.B(n_77),
.Y(n_652)
);

A2O1A1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_574),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_597),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_558),
.Y(n_655)
);

O2A1O1Ixp33_ASAP7_75t_L g656 ( 
.A1(n_570),
.A2(n_598),
.B(n_579),
.C(n_29),
.Y(n_656)
);

O2A1O1Ixp5_ASAP7_75t_L g657 ( 
.A1(n_550),
.A2(n_156),
.B(n_241),
.C(n_240),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_548),
.B(n_27),
.Y(n_658)
);

OAI21xp5_ASAP7_75t_L g659 ( 
.A1(n_577),
.A2(n_82),
.B(n_81),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_606),
.Y(n_660)
);

AO32x2_ASAP7_75t_L g661 ( 
.A1(n_650),
.A2(n_28),
.A3(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_661)
);

AO21x2_ASAP7_75t_L g662 ( 
.A1(n_603),
.A2(n_628),
.B(n_626),
.Y(n_662)
);

O2A1O1Ixp33_ASAP7_75t_SL g663 ( 
.A1(n_658),
.A2(n_158),
.B(n_239),
.C(n_238),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_651),
.Y(n_664)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_638),
.A2(n_630),
.B(n_620),
.Y(n_665)
);

OAI21x1_ASAP7_75t_L g666 ( 
.A1(n_613),
.A2(n_648),
.B(n_637),
.Y(n_666)
);

BUFx12f_ASAP7_75t_L g667 ( 
.A(n_639),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_615),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_668)
);

A2O1A1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_604),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_639),
.Y(n_670)
);

A2O1A1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_625),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_671)
);

BUFx12f_ASAP7_75t_L g672 ( 
.A(n_639),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_SL g673 ( 
.A(n_623),
.B(n_36),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_616),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_614),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_646),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_605),
.B(n_37),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_612),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_607),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_679)
);

NOR2xp67_ASAP7_75t_SL g680 ( 
.A(n_622),
.B(n_38),
.Y(n_680)
);

OAI21x1_ASAP7_75t_L g681 ( 
.A1(n_657),
.A2(n_163),
.B(n_237),
.Y(n_681)
);

BUFx12f_ASAP7_75t_L g682 ( 
.A(n_655),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_659),
.A2(n_246),
.B(n_160),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_659),
.A2(n_236),
.B(n_159),
.Y(n_684)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_656),
.A2(n_157),
.B(n_234),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_642),
.A2(n_155),
.B(n_233),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_617),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_611),
.Y(n_688)
);

OAI21x1_ASAP7_75t_L g689 ( 
.A1(n_642),
.A2(n_164),
.B(n_232),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_634),
.Y(n_690)
);

A2O1A1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_619),
.A2(n_40),
.B(n_41),
.C(n_83),
.Y(n_691)
);

O2A1O1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_633),
.A2(n_84),
.B(n_85),
.C(n_86),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_610),
.B(n_87),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_624),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_L g695 ( 
.A1(n_640),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_647),
.Y(n_696)
);

NAND2x1p5_ASAP7_75t_L g697 ( 
.A(n_610),
.B(n_91),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_608),
.A2(n_235),
.B(n_94),
.Y(n_698)
);

OAI22xp33_ASAP7_75t_L g699 ( 
.A1(n_618),
.A2(n_92),
.B1(n_96),
.B2(n_97),
.Y(n_699)
);

AOI22x1_ASAP7_75t_L g700 ( 
.A1(n_645),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_621),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_652),
.A2(n_105),
.B(n_106),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_627),
.A2(n_107),
.B(n_109),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_608),
.B(n_111),
.Y(n_704)
);

AOI21x1_ASAP7_75t_L g705 ( 
.A1(n_649),
.A2(n_112),
.B(n_113),
.Y(n_705)
);

O2A1O1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_629),
.A2(n_114),
.B(n_115),
.C(n_116),
.Y(n_706)
);

BUFx12f_ASAP7_75t_L g707 ( 
.A(n_644),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_654),
.A2(n_117),
.B(n_118),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_640),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_636),
.A2(n_119),
.B(n_121),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_635),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_643),
.Y(n_712)
);

NAND3xp33_ASAP7_75t_L g713 ( 
.A(n_641),
.B(n_123),
.C(n_124),
.Y(n_713)
);

OAI21x1_ASAP7_75t_L g714 ( 
.A1(n_632),
.A2(n_125),
.B(n_126),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_678),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_712),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_694),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_688),
.B(n_609),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_664),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_688),
.B(n_609),
.Y(n_720)
);

INVxp67_ASAP7_75t_R g721 ( 
.A(n_677),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_701),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_670),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_696),
.B(n_609),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_711),
.Y(n_725)
);

OAI21x1_ASAP7_75t_L g726 ( 
.A1(n_665),
.A2(n_631),
.B(n_632),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_682),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_667),
.Y(n_728)
);

BUFx4f_ASAP7_75t_SL g729 ( 
.A(n_672),
.Y(n_729)
);

OAI21x1_ASAP7_75t_L g730 ( 
.A1(n_666),
.A2(n_643),
.B(n_653),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_675),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_662),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_693),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_709),
.B(n_643),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_676),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_662),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_708),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_686),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_693),
.B(n_128),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_660),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_674),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_661),
.Y(n_742)
);

OAI21xp33_ASAP7_75t_SL g743 ( 
.A1(n_683),
.A2(n_129),
.B(n_131),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_690),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_702),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_689),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_669),
.B(n_132),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_681),
.Y(n_748)
);

AOI21x1_ASAP7_75t_L g749 ( 
.A1(n_705),
.A2(n_133),
.B(n_135),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_687),
.B(n_229),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_685),
.Y(n_751)
);

HB1xp67_ASAP7_75t_SL g752 ( 
.A(n_668),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_661),
.B(n_136),
.Y(n_753)
);

OA21x2_ASAP7_75t_L g754 ( 
.A1(n_683),
.A2(n_137),
.B(n_139),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_679),
.B(n_227),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_661),
.B(n_140),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_697),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_684),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_714),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_684),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_697),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_707),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_668),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_704),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_700),
.Y(n_765)
);

OA21x2_ASAP7_75t_L g766 ( 
.A1(n_698),
.A2(n_141),
.B(n_142),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_704),
.Y(n_767)
);

OAI21x1_ASAP7_75t_L g768 ( 
.A1(n_703),
.A2(n_144),
.B(n_145),
.Y(n_768)
);

AO21x1_ASAP7_75t_SL g769 ( 
.A1(n_698),
.A2(n_146),
.B(n_148),
.Y(n_769)
);

BUFx8_ASAP7_75t_SL g770 ( 
.A(n_673),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_713),
.Y(n_771)
);

BUFx4_ASAP7_75t_R g772 ( 
.A(n_680),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_663),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_706),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_671),
.B(n_225),
.Y(n_775)
);

OA21x2_ASAP7_75t_L g776 ( 
.A1(n_703),
.A2(n_149),
.B(n_150),
.Y(n_776)
);

AO21x2_ASAP7_75t_L g777 ( 
.A1(n_695),
.A2(n_152),
.B(n_153),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_R g778 ( 
.A(n_729),
.B(n_165),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_728),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_744),
.B(n_691),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_728),
.Y(n_781)
);

OR2x6_ASAP7_75t_L g782 ( 
.A(n_739),
.B(n_710),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_722),
.B(n_695),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_R g784 ( 
.A(n_727),
.B(n_710),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_721),
.B(n_713),
.Y(n_785)
);

CKINVDCx11_ASAP7_75t_R g786 ( 
.A(n_728),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_715),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_716),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_723),
.Y(n_789)
);

NAND2xp33_ASAP7_75t_R g790 ( 
.A(n_762),
.B(n_166),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_731),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_733),
.B(n_169),
.Y(n_792)
);

CKINVDCx8_ASAP7_75t_R g793 ( 
.A(n_739),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_R g794 ( 
.A(n_762),
.B(n_170),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_733),
.B(n_171),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_761),
.B(n_172),
.Y(n_796)
);

BUFx8_ASAP7_75t_SL g797 ( 
.A(n_770),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_744),
.B(n_699),
.Y(n_798)
);

NOR2x1_ASAP7_75t_L g799 ( 
.A(n_762),
.B(n_706),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_767),
.B(n_692),
.Y(n_800)
);

BUFx10_ASAP7_75t_L g801 ( 
.A(n_731),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_762),
.Y(n_802)
);

BUFx10_ASAP7_75t_L g803 ( 
.A(n_739),
.Y(n_803)
);

NAND2x1p5_ASAP7_75t_L g804 ( 
.A(n_739),
.B(n_692),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_719),
.B(n_174),
.Y(n_805)
);

NAND2xp33_ASAP7_75t_R g806 ( 
.A(n_766),
.B(n_175),
.Y(n_806)
);

OR2x6_ASAP7_75t_L g807 ( 
.A(n_757),
.B(n_176),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_721),
.B(n_178),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_761),
.B(n_179),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_R g810 ( 
.A(n_766),
.B(n_754),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_R g811 ( 
.A(n_752),
.B(n_224),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_719),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_757),
.B(n_180),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_772),
.B(n_764),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_757),
.B(n_181),
.Y(n_815)
);

NAND2x1p5_ASAP7_75t_L g816 ( 
.A(n_757),
.B(n_183),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_767),
.B(n_184),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_740),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_740),
.B(n_185),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_724),
.B(n_190),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_716),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_767),
.B(n_191),
.Y(n_822)
);

NAND2xp33_ASAP7_75t_R g823 ( 
.A(n_766),
.B(n_192),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_741),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_717),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_741),
.B(n_193),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_R g827 ( 
.A(n_764),
.B(n_223),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_717),
.B(n_194),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_R g829 ( 
.A(n_766),
.B(n_195),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_735),
.Y(n_830)
);

XOR2xp5_ASAP7_75t_L g831 ( 
.A(n_755),
.B(n_196),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_735),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_788),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_830),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_791),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_821),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_825),
.Y(n_837)
);

NOR2x1_ASAP7_75t_SL g838 ( 
.A(n_782),
.B(n_777),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_832),
.Y(n_839)
);

NAND2x1p5_ASAP7_75t_L g840 ( 
.A(n_799),
.B(n_760),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_812),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_818),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_824),
.B(n_718),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_785),
.B(n_718),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_787),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_789),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_800),
.Y(n_847)
);

AND2x4_ASAP7_75t_SL g848 ( 
.A(n_782),
.B(n_759),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_805),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_780),
.Y(n_850)
);

BUFx4f_ASAP7_75t_SL g851 ( 
.A(n_779),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_783),
.A2(n_760),
.B1(n_777),
.B2(n_758),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_804),
.A2(n_777),
.B1(n_758),
.B2(n_747),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_820),
.B(n_742),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_814),
.B(n_742),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_817),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_806),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_801),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_813),
.B(n_759),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_798),
.B(n_720),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_831),
.A2(n_747),
.B1(n_771),
.B2(n_775),
.Y(n_861)
);

OAI221xp5_ASAP7_75t_L g862 ( 
.A1(n_790),
.A2(n_743),
.B1(n_750),
.B2(n_771),
.C(n_774),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_828),
.B(n_753),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_828),
.B(n_753),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_822),
.Y(n_865)
);

OAI221xp5_ASAP7_75t_L g866 ( 
.A1(n_823),
.A2(n_743),
.B1(n_774),
.B2(n_763),
.C(n_765),
.Y(n_866)
);

NOR2x1_ASAP7_75t_L g867 ( 
.A(n_781),
.B(n_734),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_807),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_813),
.B(n_759),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_808),
.B(n_720),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_796),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_807),
.B(n_736),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_815),
.B(n_738),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_796),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_809),
.B(n_756),
.Y(n_875)
);

INVxp67_ASAP7_75t_SL g876 ( 
.A(n_829),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_810),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_809),
.B(n_724),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_815),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_819),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_793),
.B(n_756),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_819),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_784),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_826),
.B(n_736),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_811),
.A2(n_769),
.B1(n_763),
.B2(n_754),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_802),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_826),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_803),
.B(n_732),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_833),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_883),
.B(n_734),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_877),
.B(n_732),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_833),
.Y(n_892)
);

OAI31xp33_ASAP7_75t_L g893 ( 
.A1(n_862),
.A2(n_816),
.A3(n_792),
.B(n_795),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_837),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_837),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_867),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_836),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_836),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_839),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_839),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_867),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_839),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_853),
.A2(n_754),
.B(n_776),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_855),
.B(n_732),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_855),
.B(n_751),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_847),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_847),
.B(n_725),
.Y(n_907)
);

OAI33xp33_ASAP7_75t_L g908 ( 
.A1(n_850),
.A2(n_725),
.A3(n_765),
.B1(n_773),
.B2(n_737),
.B3(n_738),
.Y(n_908)
);

NAND4xp25_ASAP7_75t_L g909 ( 
.A(n_852),
.B(n_773),
.C(n_795),
.D(n_792),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_850),
.B(n_751),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_846),
.B(n_738),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_860),
.B(n_746),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_L g913 ( 
.A(n_861),
.B(n_754),
.C(n_776),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_841),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_841),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_854),
.B(n_746),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_834),
.Y(n_917)
);

OAI33xp33_ASAP7_75t_L g918 ( 
.A1(n_843),
.A2(n_737),
.A3(n_746),
.B1(n_748),
.B2(n_745),
.B3(n_786),
.Y(n_918)
);

NOR2x1_ASAP7_75t_L g919 ( 
.A(n_842),
.B(n_776),
.Y(n_919)
);

AOI221xp5_ASAP7_75t_L g920 ( 
.A1(n_866),
.A2(n_794),
.B1(n_827),
.B2(n_778),
.C(n_748),
.Y(n_920)
);

OAI31xp33_ASAP7_75t_L g921 ( 
.A1(n_857),
.A2(n_769),
.A3(n_745),
.B(n_776),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_849),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_849),
.Y(n_923)
);

AOI21xp33_ASAP7_75t_L g924 ( 
.A1(n_876),
.A2(n_768),
.B(n_730),
.Y(n_924)
);

OAI33xp33_ASAP7_75t_L g925 ( 
.A1(n_844),
.A2(n_835),
.A3(n_870),
.B1(n_882),
.B2(n_880),
.B3(n_878),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_854),
.B(n_730),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_838),
.B(n_726),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_926),
.B(n_838),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_917),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_926),
.B(n_848),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_889),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_911),
.B(n_849),
.Y(n_932)
);

OR2x2_ASAP7_75t_L g933 ( 
.A(n_922),
.B(n_840),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_892),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_905),
.B(n_848),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_897),
.B(n_848),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_898),
.B(n_834),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_905),
.B(n_891),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_891),
.B(n_840),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_896),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_899),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_922),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_896),
.B(n_916),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_916),
.B(n_840),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_894),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_920),
.A2(n_868),
.B1(n_879),
.B2(n_885),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_901),
.B(n_881),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_906),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_890),
.B(n_865),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_895),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_890),
.B(n_865),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_904),
.B(n_923),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_900),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_914),
.B(n_842),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_925),
.B(n_845),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_902),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_915),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_907),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_955),
.B(n_910),
.Y(n_959)
);

AO221x2_ASAP7_75t_L g960 ( 
.A1(n_949),
.A2(n_913),
.B1(n_880),
.B2(n_882),
.C(n_879),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_931),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_958),
.B(n_910),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_946),
.A2(n_868),
.B1(n_909),
.B2(n_918),
.Y(n_963)
);

INVxp67_ASAP7_75t_L g964 ( 
.A(n_947),
.Y(n_964)
);

OAI22xp33_ASAP7_75t_L g965 ( 
.A1(n_951),
.A2(n_868),
.B1(n_903),
.B2(n_872),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_948),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_932),
.B(n_912),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_929),
.B(n_904),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_947),
.A2(n_868),
.B1(n_908),
.B2(n_881),
.Y(n_969)
);

OAI22xp33_ASAP7_75t_L g970 ( 
.A1(n_940),
.A2(n_872),
.B1(n_887),
.B2(n_874),
.Y(n_970)
);

NOR4xp25_ASAP7_75t_SL g971 ( 
.A(n_957),
.B(n_924),
.C(n_893),
.D(n_921),
.Y(n_971)
);

NAND2xp33_ASAP7_75t_SL g972 ( 
.A(n_939),
.B(n_886),
.Y(n_972)
);

INVxp67_ASAP7_75t_SL g973 ( 
.A(n_933),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_937),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_964),
.B(n_939),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_959),
.B(n_934),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_966),
.B(n_944),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_974),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_968),
.B(n_933),
.Y(n_979)
);

NOR2x1_ASAP7_75t_L g980 ( 
.A(n_961),
.B(n_940),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_962),
.B(n_945),
.Y(n_981)
);

NAND3x1_ASAP7_75t_L g982 ( 
.A(n_963),
.B(n_943),
.C(n_928),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_973),
.B(n_944),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_967),
.B(n_928),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_960),
.B(n_938),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_960),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_972),
.B(n_937),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_SL g988 ( 
.A1(n_986),
.A2(n_969),
.B(n_965),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_978),
.Y(n_989)
);

OAI221xp5_ASAP7_75t_L g990 ( 
.A1(n_987),
.A2(n_971),
.B1(n_858),
.B2(n_950),
.C(n_957),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_981),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_976),
.A2(n_927),
.B1(n_856),
.B2(n_865),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_981),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_976),
.B(n_943),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_977),
.Y(n_995)
);

OAI211xp5_ASAP7_75t_L g996 ( 
.A1(n_980),
.A2(n_927),
.B(n_919),
.C(n_858),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_989),
.B(n_975),
.Y(n_997)
);

NAND2xp33_ASAP7_75t_L g998 ( 
.A(n_989),
.B(n_982),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_995),
.B(n_985),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_991),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_993),
.B(n_983),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_997),
.B(n_1000),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_1001),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_999),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_998),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_1000),
.Y(n_1006)
);

NOR2x1_ASAP7_75t_L g1007 ( 
.A(n_1005),
.B(n_990),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_1002),
.B(n_994),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_1006),
.B(n_984),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1004),
.Y(n_1010)
);

NOR2x1_ASAP7_75t_L g1011 ( 
.A(n_1003),
.B(n_988),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_1006),
.B(n_988),
.Y(n_1012)
);

NOR3xp33_ASAP7_75t_L g1013 ( 
.A(n_1005),
.B(n_996),
.C(n_970),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1010),
.Y(n_1014)
);

AOI222xp33_ASAP7_75t_L g1015 ( 
.A1(n_1011),
.A2(n_992),
.B1(n_851),
.B2(n_863),
.C1(n_864),
.C2(n_937),
.Y(n_1015)
);

AOI211x1_ASAP7_75t_L g1016 ( 
.A1(n_1012),
.A2(n_956),
.B(n_941),
.C(n_953),
.Y(n_1016)
);

OAI211xp5_ASAP7_75t_L g1017 ( 
.A1(n_1007),
.A2(n_979),
.B(n_797),
.C(n_856),
.Y(n_1017)
);

AOI211xp5_ASAP7_75t_L g1018 ( 
.A1(n_1013),
.A2(n_936),
.B(n_768),
.C(n_874),
.Y(n_1018)
);

AOI221xp5_ASAP7_75t_L g1019 ( 
.A1(n_1009),
.A2(n_954),
.B1(n_956),
.B2(n_941),
.C(n_942),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_1014),
.B(n_1008),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_1017),
.B(n_938),
.Y(n_1021)
);

XOR2xp5_ASAP7_75t_L g1022 ( 
.A(n_1018),
.B(n_871),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_1015),
.A2(n_1019),
.B1(n_936),
.B2(n_1016),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_1014),
.Y(n_1024)
);

NAND4xp75_ASAP7_75t_L g1025 ( 
.A(n_1014),
.B(n_930),
.C(n_935),
.D(n_863),
.Y(n_1025)
);

NAND4xp75_ASAP7_75t_L g1026 ( 
.A(n_1014),
.B(n_930),
.C(n_935),
.D(n_864),
.Y(n_1026)
);

XNOR2xp5_ASAP7_75t_L g1027 ( 
.A(n_1020),
.B(n_936),
.Y(n_1027)
);

XNOR2xp5_ASAP7_75t_L g1028 ( 
.A(n_1021),
.B(n_871),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_1024),
.B(n_954),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_1023),
.B(n_954),
.Y(n_1030)
);

XNOR2x1_ASAP7_75t_L g1031 ( 
.A(n_1025),
.B(n_197),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1026),
.B(n_952),
.Y(n_1032)
);

NAND2xp33_ASAP7_75t_SL g1033 ( 
.A(n_1022),
.B(n_942),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_1020),
.B(n_952),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_R g1035 ( 
.A(n_1020),
.B(n_199),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_1035),
.Y(n_1036)
);

AO22x1_ASAP7_75t_L g1037 ( 
.A1(n_1029),
.A2(n_887),
.B1(n_875),
.B2(n_873),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_1027),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1034),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_1030),
.A2(n_873),
.B1(n_884),
.B2(n_859),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_1031),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_1033),
.A2(n_873),
.B1(n_884),
.B2(n_859),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_1028),
.Y(n_1043)
);

OR2x2_ASAP7_75t_L g1044 ( 
.A(n_1032),
.B(n_875),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_1035),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_1032),
.B(n_888),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1034),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1034),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1041),
.B(n_888),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1045),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1039),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1047),
.Y(n_1052)
);

CKINVDCx16_ASAP7_75t_R g1053 ( 
.A(n_1043),
.Y(n_1053)
);

BUFx4f_ASAP7_75t_L g1054 ( 
.A(n_1036),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1048),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1053),
.B(n_1038),
.Y(n_1056)
);

NOR2xp67_ASAP7_75t_L g1057 ( 
.A(n_1051),
.B(n_1046),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1052),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1055),
.B(n_1044),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1050),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_1060),
.A2(n_1054),
.B1(n_1049),
.B2(n_1042),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_SL g1062 ( 
.A1(n_1056),
.A2(n_1040),
.B1(n_1037),
.B2(n_873),
.Y(n_1062)
);

AOI31xp33_ASAP7_75t_L g1063 ( 
.A1(n_1059),
.A2(n_200),
.A3(n_201),
.B(n_205),
.Y(n_1063)
);

AOI31xp33_ASAP7_75t_L g1064 ( 
.A1(n_1058),
.A2(n_207),
.A3(n_209),
.B(n_210),
.Y(n_1064)
);

OAI222xp33_ASAP7_75t_L g1065 ( 
.A1(n_1061),
.A2(n_1057),
.B1(n_749),
.B2(n_869),
.C1(n_859),
.C2(n_217),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_1063),
.A2(n_211),
.B(n_214),
.C(n_216),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1066),
.Y(n_1067)
);

BUFx4_ASAP7_75t_R g1068 ( 
.A(n_1065),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1068),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1067),
.Y(n_1070)
);

OAI221xp5_ASAP7_75t_R g1071 ( 
.A1(n_1069),
.A2(n_1062),
.B1(n_1064),
.B2(n_219),
.C(n_220),
.Y(n_1071)
);

AOI211xp5_ASAP7_75t_L g1072 ( 
.A1(n_1071),
.A2(n_1070),
.B(n_218),
.C(n_221),
.Y(n_1072)
);


endmodule