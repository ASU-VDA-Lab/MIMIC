module fake_jpeg_12274_n_171 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_171);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_12),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_20),
.B(n_31),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_16),
.B(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_5),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

BUFx4f_ASAP7_75t_SL g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_1),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_2),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_2),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_68),
.B1(n_64),
.B2(n_51),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_74),
.B1(n_78),
.B2(n_68),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_80),
.A2(n_59),
.B1(n_60),
.B2(n_57),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_55),
.B1(n_68),
.B2(n_57),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_93),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_50),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_98),
.B(n_99),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_29),
.B1(n_47),
.B2(n_46),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_72),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_73),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_112),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g105 ( 
.A(n_93),
.B(n_64),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_105),
.A2(n_117),
.B(n_118),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_78),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_108),
.C(n_111),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_65),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_62),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_51),
.B1(n_52),
.B2(n_70),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_9),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_89),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_87),
.B(n_67),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_116),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_69),
.C(n_66),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_121),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_55),
.B(n_66),
.C(n_6),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_3),
.B(n_4),
.C(n_7),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_3),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_123),
.A2(n_128),
.B1(n_136),
.B2(n_142),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_130),
.B1(n_33),
.B2(n_35),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_28),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_129),
.B(n_139),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_130)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_11),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_134),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_48),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_110),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_13),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_138),
.A2(n_30),
.B(n_32),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_115),
.B(n_19),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_22),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_141),
.B(n_36),
.Y(n_154)
);

AO21x2_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_110),
.B(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_24),
.C(n_26),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_139),
.C(n_129),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_155),
.B(n_135),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_152),
.Y(n_161)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

AOI322xp5_ASAP7_75t_SL g157 ( 
.A1(n_153),
.A2(n_154),
.A3(n_125),
.B1(n_122),
.B2(n_141),
.C1(n_42),
.C2(n_41),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_157),
.B(n_158),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_147),
.B1(n_145),
.B2(n_151),
.Y(n_164)
);

AO221x1_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_144),
.B1(n_155),
.B2(n_132),
.C(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_163),
.B(n_156),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_161),
.C(n_138),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_166),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_163),
.B(n_162),
.Y(n_168)
);

XOR2x1_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_143),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_143),
.B(n_157),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_37),
.Y(n_171)
);


endmodule