module fake_jpeg_3499_n_425 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_425);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_425;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_8),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_56),
.B(n_70),
.Y(n_166)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_19),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_58),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_60),
.Y(n_207)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_61),
.Y(n_178)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_62),
.Y(n_191)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_21),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_64),
.B(n_66),
.Y(n_129)
);

BUFx2_ASAP7_75t_R g65 ( 
.A(n_21),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_65),
.Y(n_148)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_67),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_21),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_68),
.B(n_82),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_23),
.B(n_8),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_69),
.B(n_75),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_27),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_23),
.B(n_9),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_77),
.Y(n_173)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_78),
.Y(n_196)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_22),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_83),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_24),
.B(n_7),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_84),
.B(n_89),
.Y(n_153)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_86),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_87),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_32),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_88),
.B(n_96),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_41),
.B(n_18),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_24),
.B(n_7),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_91),
.B(n_95),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_93),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_94),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_25),
.B(n_12),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g96 ( 
.A(n_28),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_97),
.Y(n_181)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_106),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_99),
.Y(n_193)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_100),
.Y(n_200)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_105),
.Y(n_124)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_103),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_25),
.B(n_12),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_104),
.B(n_113),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_107),
.B(n_109),
.Y(n_162)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

AO22x1_ASAP7_75t_L g160 ( 
.A1(n_108),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_32),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_110),
.B(n_111),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_112),
.B(n_115),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_27),
.B(n_6),
.Y(n_113)
);

BUFx6f_ASAP7_75t_SL g114 ( 
.A(n_55),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_114),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_42),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_28),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_116),
.B(n_121),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_42),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_42),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_120),
.B(n_122),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_42),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_40),
.B(n_6),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_29),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_123),
.B(n_100),
.Y(n_190)
);

OAI22x1_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_36),
.B1(n_26),
.B2(n_53),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_125),
.B(n_205),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_52),
.B1(n_54),
.B2(n_49),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_126),
.A2(n_137),
.B1(n_138),
.B2(n_144),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_79),
.A2(n_55),
.B1(n_34),
.B2(n_51),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_127),
.A2(n_132),
.B1(n_140),
.B2(n_141),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_53),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_131),
.B(n_135),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_78),
.A2(n_31),
.B1(n_37),
.B2(n_51),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_37),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_80),
.A2(n_52),
.B1(n_118),
.B2(n_117),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_83),
.A2(n_54),
.B1(n_46),
.B2(n_49),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_60),
.A2(n_31),
.B1(n_50),
.B2(n_48),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_74),
.A2(n_40),
.B1(n_50),
.B2(n_48),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_87),
.A2(n_99),
.B1(n_97),
.B2(n_58),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_L g146 ( 
.A1(n_81),
.A2(n_54),
.B1(n_49),
.B2(n_46),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_146),
.A2(n_172),
.B1(n_174),
.B2(n_197),
.Y(n_210)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_59),
.A2(n_54),
.B1(n_49),
.B2(n_46),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g217 ( 
.A1(n_147),
.A2(n_146),
.A3(n_160),
.B1(n_187),
.B2(n_149),
.Y(n_217)
);

AO22x1_ASAP7_75t_SL g149 ( 
.A1(n_101),
.A2(n_46),
.B1(n_2),
.B2(n_3),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_149),
.B(n_182),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_45),
.B1(n_43),
.B2(n_15),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_150),
.A2(n_184),
.B1(n_186),
.B2(n_208),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_43),
.B1(n_45),
.B2(n_3),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_151),
.A2(n_161),
.B1(n_164),
.B2(n_170),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_65),
.B(n_14),
.C(n_16),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_155),
.B(n_172),
.C(n_149),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_108),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_57),
.A2(n_1),
.B1(n_4),
.B2(n_16),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_77),
.A2(n_4),
.B1(n_18),
.B2(n_90),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_93),
.A2(n_67),
.B1(n_103),
.B2(n_86),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_86),
.A2(n_18),
.B1(n_116),
.B2(n_94),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_94),
.A2(n_105),
.B1(n_116),
.B2(n_56),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_105),
.A2(n_36),
.B1(n_55),
.B2(n_35),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_176),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_56),
.B(n_70),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_70),
.A2(n_56),
.B1(n_115),
.B2(n_121),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_56),
.B(n_70),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_185),
.B(n_187),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_70),
.A2(n_56),
.B1(n_122),
.B2(n_89),
.Y(n_186)
);

AO22x1_ASAP7_75t_SL g187 ( 
.A1(n_63),
.A2(n_58),
.B1(n_76),
.B2(n_78),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_148),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_122),
.B(n_69),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_194),
.B(n_199),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_56),
.B(n_70),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_195),
.B(n_155),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_70),
.A2(n_56),
.B1(n_68),
.B2(n_121),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_122),
.B(n_69),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_122),
.B(n_69),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_201),
.B(n_206),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_70),
.A2(n_56),
.B1(n_68),
.B2(n_121),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_203),
.A2(n_166),
.B1(n_195),
.B2(n_188),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_70),
.A2(n_122),
.B1(n_47),
.B2(n_121),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_204),
.A2(n_203),
.B1(n_147),
.B2(n_187),
.Y(n_237)
);

OR2x2_ASAP7_75t_SL g205 ( 
.A(n_70),
.B(n_35),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_122),
.B(n_69),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_70),
.A2(n_56),
.B1(n_115),
.B2(n_121),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_202),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_212),
.B(n_217),
.Y(n_287)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_213),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_133),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_125),
.A2(n_135),
.B(n_124),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_216),
.A2(n_244),
.B(n_241),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_124),
.B(n_131),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_218),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_158),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_219),
.B(n_224),
.Y(n_279)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_134),
.B(n_168),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_222),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_153),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_129),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_124),
.B(n_136),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_225),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_191),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_227),
.B(n_228),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_159),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_230),
.Y(n_295)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_133),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_152),
.B(n_189),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_235),
.B(n_243),
.Y(n_280)
);

AND2x4_ASAP7_75t_SL g236 ( 
.A(n_205),
.B(n_197),
.Y(n_236)
);

NAND2x1_ASAP7_75t_SL g281 ( 
.A(n_236),
.B(n_245),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_237),
.A2(n_254),
.B1(n_239),
.B2(n_210),
.Y(n_288)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_165),
.B(n_130),
.Y(n_243)
);

AND2x2_ASAP7_75t_SL g245 ( 
.A(n_174),
.B(n_142),
.Y(n_245)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_173),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_175),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_145),
.B(n_128),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_251),
.Y(n_306)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_181),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_147),
.B(n_162),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_266),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_147),
.A2(n_160),
.B1(n_139),
.B2(n_128),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_139),
.B(n_145),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_256),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_169),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_196),
.B(n_163),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_257),
.A2(n_216),
.B(n_251),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_177),
.B(n_196),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_259),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_177),
.B(n_143),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_143),
.B(n_180),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_260),
.B(n_261),
.Y(n_300)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_175),
.Y(n_261)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_169),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_154),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_265),
.Y(n_302)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_154),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_267),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_163),
.B(n_207),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_193),
.B(n_192),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_193),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_192),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_157),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_270),
.Y(n_305)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_156),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_157),
.Y(n_272)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_167),
.B(n_134),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_274),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_182),
.B(n_185),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_240),
.A2(n_253),
.B1(n_241),
.B2(n_244),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_282),
.A2(n_288),
.B1(n_298),
.B2(n_242),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_234),
.A2(n_226),
.B1(n_210),
.B2(n_225),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_283),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_284),
.Y(n_319)
);

AND2x6_ASAP7_75t_L g285 ( 
.A(n_236),
.B(n_247),
.Y(n_285)
);

AOI21xp33_ASAP7_75t_L g325 ( 
.A1(n_285),
.A2(n_233),
.B(n_272),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_223),
.B(n_274),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_290),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_223),
.B(n_240),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_292),
.A2(n_307),
.B(n_215),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_212),
.B(n_218),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_303),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_245),
.A2(n_248),
.B1(n_217),
.B2(n_236),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_246),
.A2(n_218),
.B1(n_245),
.B2(n_234),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_229),
.B1(n_269),
.B2(n_266),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_214),
.B(n_225),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_226),
.A2(n_214),
.B1(n_257),
.B2(n_251),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_276),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_309),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_211),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_310),
.Y(n_344)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_294),
.Y(n_311)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_311),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_312),
.B(n_314),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_289),
.B(n_230),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_315),
.B(n_316),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_290),
.B(n_213),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_280),
.B(n_209),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_317),
.B(n_318),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_264),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_304),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_320),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_302),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_324),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_257),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_322),
.A2(n_334),
.B(n_339),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_263),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_281),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_270),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_326),
.B(n_330),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_292),
.A2(n_249),
.B(n_220),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_327),
.A2(n_340),
.B(n_284),
.Y(n_362)
);

INVx13_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_329),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_278),
.B(n_282),
.Y(n_330)
);

AND2x2_ASAP7_75t_SL g331 ( 
.A(n_278),
.B(n_250),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_295),
.Y(n_332)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_332),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_288),
.A2(n_267),
.B1(n_252),
.B2(n_231),
.Y(n_333)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_333),
.Y(n_351)
);

NOR2x1_ASAP7_75t_L g334 ( 
.A(n_299),
.B(n_238),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_304),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_295),
.Y(n_336)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_336),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_298),
.A2(n_262),
.B1(n_268),
.B2(n_232),
.Y(n_337)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_337),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_304),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_300),
.B(n_271),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_324),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_346),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_330),
.B(n_285),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_319),
.Y(n_366)
);

A2O1A1Ixp33_ASAP7_75t_L g358 ( 
.A1(n_328),
.A2(n_287),
.B(n_275),
.C(n_281),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_339),
.Y(n_359)
);

INVx13_ASAP7_75t_L g365 ( 
.A(n_359),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_313),
.B(n_287),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_320),
.A2(n_306),
.B1(n_296),
.B2(n_291),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_361),
.A2(n_296),
.B1(n_303),
.B2(n_338),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_362),
.A2(n_281),
.B(n_314),
.Y(n_378)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_310),
.Y(n_363)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_363),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_366),
.B(n_347),
.Y(n_396)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_344),
.Y(n_368)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_368),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_362),
.A2(n_323),
.B(n_340),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_369),
.A2(n_376),
.B(n_377),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_357),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_344),
.Y(n_372)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_372),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_373),
.A2(n_380),
.B1(n_381),
.B2(n_387),
.Y(n_390)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_345),
.Y(n_374)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_374),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_342),
.B(n_308),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_375),
.B(n_384),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_353),
.A2(n_327),
.B(n_334),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_353),
.A2(n_334),
.B(n_319),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_378),
.A2(n_352),
.B(n_356),
.Y(n_395)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_345),
.Y(n_379)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_379),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_364),
.A2(n_312),
.B1(n_337),
.B2(n_313),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_364),
.A2(n_316),
.B1(n_333),
.B2(n_315),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_349),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_349),
.Y(n_383)
);

INVxp33_ASAP7_75t_SL g400 ( 
.A(n_383),
.Y(n_400)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_354),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_354),
.Y(n_385)
);

INVx13_ASAP7_75t_L g386 ( 
.A(n_341),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_346),
.B(n_321),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_380),
.A2(n_355),
.B1(n_358),
.B2(n_348),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_395),
.A2(n_341),
.B(n_385),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_396),
.B(n_378),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_371),
.A2(n_355),
.B1(n_351),
.B2(n_343),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_381),
.A2(n_351),
.B1(n_331),
.B2(n_360),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_398),
.A2(n_401),
.B1(n_367),
.B2(n_384),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_369),
.A2(n_331),
.B1(n_335),
.B2(n_350),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_388),
.A2(n_397),
.B1(n_393),
.B2(n_390),
.Y(n_402)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_402),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_389),
.Y(n_403)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_403),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_404),
.B(n_407),
.Y(n_409)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_400),
.Y(n_405)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_405),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_393),
.A2(n_370),
.B1(n_365),
.B2(n_331),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_408),
.A2(n_399),
.B1(n_394),
.B2(n_392),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_413),
.B(n_406),
.Y(n_414)
);

OAI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_414),
.A2(n_415),
.B1(n_412),
.B2(n_411),
.Y(n_418)
);

INVx11_ASAP7_75t_L g415 ( 
.A(n_410),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_409),
.B(n_404),
.C(n_405),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_416),
.B(n_412),
.C(n_413),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_417),
.B(n_418),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_418),
.Y(n_420)
);

AOI322xp5_ASAP7_75t_L g421 ( 
.A1(n_419),
.A2(n_415),
.A3(n_391),
.B1(n_392),
.B2(n_379),
.C1(n_368),
.C2(n_367),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_421),
.B(n_383),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_422),
.A2(n_372),
.B(n_382),
.Y(n_423)
);

A2O1A1Ixp33_ASAP7_75t_L g424 ( 
.A1(n_423),
.A2(n_420),
.B(n_374),
.C(n_386),
.Y(n_424)
);

HAxp5_ASAP7_75t_SL g425 ( 
.A(n_424),
.B(n_329),
.CON(n_425),
.SN(n_425)
);


endmodule