module fake_jpeg_9721_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx10_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_13),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx11_ASAP7_75t_SL g67 ( 
.A(n_2),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_0),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_1),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_1),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_57),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx5_ASAP7_75t_SL g91 ( 
.A(n_77),
.Y(n_91)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_78),
.A2(n_63),
.B1(n_66),
.B2(n_60),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_58),
.B1(n_50),
.B2(n_61),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_79),
.A2(n_90),
.B1(n_95),
.B2(n_96),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_55),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_87),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_98),
.B1(n_80),
.B2(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_4),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_94),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_48),
.B1(n_46),
.B2(n_45),
.Y(n_90)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_51),
.B1(n_52),
.B2(n_67),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_68),
.A2(n_26),
.B1(n_8),
.B2(n_10),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_97),
.B1(n_91),
.B2(n_83),
.Y(n_102)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_96),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_86),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_100),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_115),
.B(n_116),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_113),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_112),
.B1(n_106),
.B2(n_103),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_118),
.A2(n_100),
.B1(n_104),
.B2(n_111),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_107),
.C(n_110),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_109),
.B1(n_108),
.B2(n_101),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_16),
.B(n_17),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_19),
.C(n_20),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_21),
.Y(n_127)
);

AO21x1_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_22),
.B(n_24),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_128),
.A2(n_29),
.B(n_32),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_33),
.B(n_34),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_35),
.C(n_39),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_131),
.Y(n_132)
);


endmodule