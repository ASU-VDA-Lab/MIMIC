module fake_ibex_1080_n_2960 (n_151, n_85, n_507, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_114, n_236, n_34, n_376, n_377, n_531, n_15, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_527, n_465, n_48, n_325, n_57, n_301, n_496, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_13, n_122, n_523, n_116, n_370, n_431, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_490, n_52, n_448, n_99, n_466, n_269, n_156, n_126, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_514, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_484, n_480, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_516, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_199, n_495, n_410, n_308, n_463, n_411, n_135, n_520, n_512, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_517, n_211, n_218, n_314, n_132, n_277, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_382, n_502, n_532, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_476, n_461, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_311, n_406, n_97, n_197, n_528, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_425, n_2960);

input n_151;
input n_85;
input n_507;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_531;
input n_15;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_523;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_490;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_126;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_514;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_480;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_516;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_199;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_520;
input n_512;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_476;
input n_461;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2960;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_1079;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1954;
wire n_1859;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_2955;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_1308;
wire n_556;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2391;
wire n_2151;
wire n_1391;
wire n_667;
wire n_884;
wire n_2396;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2724;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2605;
wire n_2343;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_641;
wire n_557;
wire n_1937;
wire n_2311;
wire n_893;
wire n_1654;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_538;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_852;
wire n_1427;
wire n_1133;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2814;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_1955;
wire n_917;
wire n_2413;
wire n_2249;
wire n_2362;
wire n_968;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_2906;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_553;
wire n_554;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_2373;
wire n_630;
wire n_1869;
wire n_567;
wire n_2275;
wire n_1853;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_971;
wire n_1326;
wire n_702;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_2541;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_2723;
wire n_1616;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_1281;
wire n_1447;
wire n_2451;
wire n_2166;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_2256;
wire n_606;
wire n_737;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2879;
wire n_2958;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_864;
wire n_608;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_2821;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_591;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_2838;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_594;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_660;
wire n_2590;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_576;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_607;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_2954;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2823;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_2905;
wire n_803;
wire n_2570;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_2095;
wire n_555;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_2903;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_2463;
wire n_2654;
wire n_717;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_668;
wire n_871;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_588;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_2298;
wire n_2771;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_545;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_2862;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2683;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_598;
wire n_2141;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_2566;
wire n_1991;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_2180;
wire n_1952;
wire n_2087;
wire n_2920;
wire n_604;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2555;
wire n_2639;
wire n_2330;
wire n_636;
wire n_1259;
wire n_2108;
wire n_2535;
wire n_595;
wire n_1001;
wire n_2945;
wire n_570;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2709;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2437;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_2665;
wire n_1124;
wire n_611;
wire n_1690;
wire n_2688;
wire n_2881;
wire n_1673;
wire n_2018;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2320;
wire n_2237;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_2758;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_571;
wire n_648;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_2447;
wire n_2818;
wire n_1057;
wire n_1473;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_775;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_535;
wire n_1956;
wire n_681;
wire n_2608;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2861;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2576;
wire n_786;
wire n_2348;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_1256;
wire n_2798;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_1961;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_688;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_2518;
wire n_2784;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2574;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_1029;
wire n_2394;
wire n_770;
wire n_1635;
wire n_1572;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_2323;
wire n_740;
wire n_549;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_1986;
wire n_2882;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_569;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_2734;
wire n_2870;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_543;
wire n_580;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2928;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_999;
wire n_2634;
wire n_1092;
wire n_1808;
wire n_560;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_2931;
wire n_2492;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2104;
wire n_949;
wire n_704;
wire n_2357;
wire n_2148;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_924;
wire n_2937;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_2092;
wire n_566;
wire n_581;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2704;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_2907;
wire n_1160;
wire n_1442;
wire n_658;
wire n_2168;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2749;
wire n_888;
wire n_2378;
wire n_1325;
wire n_2754;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_908;
wire n_1346;
wire n_565;
wire n_2834;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_415),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_105),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_226),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_491),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_236),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_195),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_449),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_48),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_83),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_452),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_221),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_152),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_366),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_533),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_48),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_8),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_32),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_23),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_44),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_266),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_132),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_18),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_317),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_376),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_339),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_414),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_52),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_441),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_59),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_352),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_309),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_422),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_354),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_458),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_381),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_530),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_461),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_21),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_144),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_118),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_203),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_435),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_49),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_142),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_108),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_113),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_479),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_289),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_114),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_258),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_336),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_84),
.Y(n_586)
);

CKINVDCx16_ASAP7_75t_R g587 ( 
.A(n_63),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_394),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_59),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_241),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_55),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_234),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_403),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_138),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_77),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_47),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_521),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_427),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_335),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_375),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_42),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_308),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_301),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_176),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_319),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_180),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_325),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_210),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_235),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_1),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_160),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_177),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_362),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_343),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_98),
.Y(n_615)
);

INVx4_ASAP7_75t_R g616 ( 
.A(n_443),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_57),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_401),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_164),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_341),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_342),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_40),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_237),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_275),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_159),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_37),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_478),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_347),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_68),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_502),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_510),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_225),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_222),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_97),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_368),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_423),
.Y(n_636)
);

BUFx8_ASAP7_75t_SL g637 ( 
.A(n_97),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_395),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_82),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_299),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_141),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_346),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_108),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_531),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_72),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_113),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_103),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_310),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_437),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_215),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_239),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_163),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_331),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_390),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_0),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_72),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_137),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_330),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_214),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_3),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_197),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_43),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_228),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_432),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_87),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_104),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_35),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_212),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_188),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_384),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_205),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_278),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_320),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_233),
.Y(n_674)
);

BUFx10_ASAP7_75t_L g675 ( 
.A(n_123),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_178),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_125),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_24),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g679 ( 
.A(n_216),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_364),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_160),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_246),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_248),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_439),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_125),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_11),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_280),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_143),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_306),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_207),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_447),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_454),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_349),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_508),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_281),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_337),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_409),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_23),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_497),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_359),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_146),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_492),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_360),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_2),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_147),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_282),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_103),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_297),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_249),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_351),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_60),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_60),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_52),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_493),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_298),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_380),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_136),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_498),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_1),
.Y(n_719)
);

CKINVDCx16_ASAP7_75t_R g720 ( 
.A(n_145),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_122),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_198),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_377),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_250),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_448),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_270),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_29),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_175),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_92),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_407),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_38),
.Y(n_731)
);

BUFx2_ASAP7_75t_SL g732 ( 
.A(n_204),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_50),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_334),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_505),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_251),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_286),
.Y(n_737)
);

BUFx10_ASAP7_75t_L g738 ( 
.A(n_173),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_527),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_393),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_119),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_18),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_149),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_220),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_481),
.Y(n_745)
);

CKINVDCx16_ASAP7_75t_R g746 ( 
.A(n_257),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_183),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_243),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_285),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_116),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_506),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_68),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_344),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_503),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_353),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_357),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_369),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_158),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_480),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_92),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_350),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_525),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_141),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_176),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_94),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_400),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_383),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_158),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_524),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_67),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_512),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_382),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_277),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_199),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_93),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_16),
.Y(n_776)
);

BUFx5_ASAP7_75t_L g777 ( 
.A(n_283),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_17),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_370),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_71),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_513),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_467),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_46),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_6),
.Y(n_784)
);

BUFx10_ASAP7_75t_L g785 ( 
.A(n_402),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_40),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_87),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_37),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_408),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_420),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_62),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_50),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_316),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_77),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_279),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_304),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_509),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_22),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_28),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_326),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_118),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_515),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_413),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_32),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_245),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_385),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_240),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_418),
.Y(n_808)
);

CKINVDCx16_ASAP7_75t_R g809 ( 
.A(n_440),
.Y(n_809)
);

BUFx10_ASAP7_75t_L g810 ( 
.A(n_71),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_230),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_6),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_80),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_96),
.Y(n_814)
);

INVxp33_ASAP7_75t_L g815 ( 
.A(n_518),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_522),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_486),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_122),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_500),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_101),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_177),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_69),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_8),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_332),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_21),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_28),
.Y(n_826)
);

BUFx8_ASAP7_75t_SL g827 ( 
.A(n_488),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_302),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_157),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_169),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_174),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_39),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_345),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_252),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_504),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_102),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_371),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_262),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_406),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_477),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_63),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_293),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_192),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_305),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_232),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_499),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_472),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_528),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_47),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_496),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_273),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_126),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_321),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_200),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_156),
.Y(n_855)
);

BUFx10_ASAP7_75t_L g856 ( 
.A(n_19),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_315),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_201),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_78),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_288),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_147),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_397),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_815),
.B(n_0),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_637),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_611),
.B(n_2),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_542),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_560),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_542),
.Y(n_868)
);

INVx4_ASAP7_75t_L g869 ( 
.A(n_785),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_550),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_587),
.B(n_3),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_720),
.B(n_4),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_619),
.B(n_4),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_611),
.B(n_5),
.Y(n_874)
);

INVx6_ASAP7_75t_L g875 ( 
.A(n_785),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_625),
.B(n_5),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_550),
.Y(n_877)
);

AND2x6_ASAP7_75t_L g878 ( 
.A(n_642),
.B(n_534),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_551),
.Y(n_879)
);

NOR2x1_ASAP7_75t_L g880 ( 
.A(n_551),
.B(n_7),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_578),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_644),
.B(n_7),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_560),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_785),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_815),
.B(n_9),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_675),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_827),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_679),
.B(n_9),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_560),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_705),
.B(n_10),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_SL g891 ( 
.A(n_618),
.B(n_182),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_560),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_684),
.B(n_10),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_600),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_827),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_578),
.B(n_11),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_675),
.Y(n_897)
);

INVx5_ASAP7_75t_L g898 ( 
.A(n_585),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_734),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_789),
.Y(n_900)
);

NOR2x1_ASAP7_75t_L g901 ( 
.A(n_586),
.B(n_12),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_675),
.B(n_12),
.Y(n_902)
);

BUFx12f_ASAP7_75t_L g903 ( 
.A(n_738),
.Y(n_903)
);

INVx5_ASAP7_75t_L g904 ( 
.A(n_585),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_738),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_585),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_585),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_590),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_586),
.Y(n_909)
);

AND2x6_ASAP7_75t_L g910 ( 
.A(n_642),
.B(n_184),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_858),
.Y(n_911)
);

INVx5_ASAP7_75t_L g912 ( 
.A(n_590),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_569),
.B(n_13),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_704),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_704),
.Y(n_915)
);

INVx5_ASAP7_75t_L g916 ( 
.A(n_590),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_659),
.B(n_13),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_728),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_738),
.B(n_14),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_728),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_590),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_810),
.Y(n_922)
);

INVx6_ASAP7_75t_L g923 ( 
.A(n_810),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_692),
.B(n_14),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_537),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_731),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_731),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_536),
.B(n_15),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_703),
.B(n_15),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_780),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_780),
.B(n_16),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_795),
.Y(n_932)
);

INVx5_ASAP7_75t_L g933 ( 
.A(n_795),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_553),
.B(n_17),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_730),
.B(n_19),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_559),
.B(n_20),
.Y(n_936)
);

INVx4_ASAP7_75t_L g937 ( 
.A(n_538),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_858),
.Y(n_938)
);

BUFx12f_ASAP7_75t_L g939 ( 
.A(n_810),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_749),
.B(n_20),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_856),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_856),
.B(n_22),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_746),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_SL g944 ( 
.A(n_809),
.B(n_532),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_856),
.B(n_553),
.Y(n_945)
);

INVx5_ASAP7_75t_L g946 ( 
.A(n_795),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_546),
.B(n_24),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_777),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_583),
.B(n_25),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_795),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_667),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_667),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_667),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_583),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_561),
.B(n_25),
.Y(n_955)
);

INVx5_ASAP7_75t_L g956 ( 
.A(n_667),
.Y(n_956)
);

BUFx12f_ASAP7_75t_L g957 ( 
.A(n_543),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_606),
.B(n_26),
.Y(n_958)
);

BUFx8_ASAP7_75t_L g959 ( 
.A(n_606),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_752),
.Y(n_960)
);

BUFx12f_ASAP7_75t_L g961 ( 
.A(n_549),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_777),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_752),
.Y(n_963)
);

BUFx12f_ASAP7_75t_L g964 ( 
.A(n_552),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_656),
.B(n_26),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_752),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_656),
.B(n_27),
.Y(n_967)
);

BUFx8_ASAP7_75t_L g968 ( 
.A(n_786),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_786),
.B(n_27),
.Y(n_969)
);

BUFx12f_ASAP7_75t_L g970 ( 
.A(n_555),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_572),
.B(n_29),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_637),
.Y(n_972)
);

BUFx8_ASAP7_75t_SL g973 ( 
.A(n_563),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_556),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_573),
.B(n_30),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_791),
.B(n_30),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_777),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_791),
.B(n_31),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_869),
.B(n_799),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_894),
.A2(n_597),
.B1(n_602),
.B2(n_535),
.Y(n_980)
);

AO22x2_ASAP7_75t_L g981 ( 
.A1(n_871),
.A2(n_743),
.B1(n_855),
.B2(n_852),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_866),
.Y(n_982)
);

AO22x2_ASAP7_75t_L g983 ( 
.A1(n_872),
.A2(n_861),
.B1(n_574),
.B2(n_615),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_865),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_974),
.Y(n_985)
);

OAI22xp33_ASAP7_75t_L g986 ( 
.A1(n_928),
.A2(n_859),
.B1(n_563),
.B2(n_595),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_899),
.A2(n_597),
.B1(n_602),
.B2(n_535),
.Y(n_987)
);

NOR2x1p5_ASAP7_75t_L g988 ( 
.A(n_903),
.B(n_764),
.Y(n_988)
);

OR2x6_ASAP7_75t_L g989 ( 
.A(n_939),
.B(n_732),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_865),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_874),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_900),
.A2(n_669),
.B1(n_708),
.B2(n_631),
.Y(n_992)
);

AND2x2_ASAP7_75t_SL g993 ( 
.A(n_891),
.B(n_944),
.Y(n_993)
);

AO22x2_ASAP7_75t_L g994 ( 
.A1(n_874),
.A2(n_617),
.B1(n_643),
.B2(n_604),
.Y(n_994)
);

OA22x2_ASAP7_75t_L g995 ( 
.A1(n_887),
.A2(n_641),
.B1(n_652),
.B2(n_610),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_870),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_882),
.A2(n_669),
.B1(n_708),
.B2(n_631),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_869),
.B(n_875),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_877),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_909),
.Y(n_1000)
);

AOI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_888),
.A2(n_772),
.B1(n_773),
.B2(n_715),
.Y(n_1001)
);

OAI22xp33_ASAP7_75t_SL g1002 ( 
.A1(n_891),
.A2(n_579),
.B1(n_580),
.B2(n_577),
.Y(n_1002)
);

OAI22xp33_ASAP7_75t_R g1003 ( 
.A1(n_973),
.A2(n_678),
.B1(n_685),
.B2(n_657),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_905),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_896),
.A2(n_772),
.B1(n_773),
.B2(n_715),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_925),
.B(n_589),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_934),
.Y(n_1007)
);

AO22x2_ASAP7_75t_L g1008 ( 
.A1(n_896),
.A2(n_688),
.B1(n_698),
.B2(n_686),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_SL g1009 ( 
.A1(n_864),
.A2(n_594),
.B1(n_666),
.B2(n_595),
.Y(n_1009)
);

AO22x2_ASAP7_75t_L g1010 ( 
.A1(n_931),
.A2(n_719),
.B1(n_721),
.B2(n_713),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_915),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_931),
.A2(n_844),
.B1(n_850),
.B2(n_802),
.Y(n_1012)
);

OAI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_947),
.A2(n_594),
.B1(n_741),
.B2(n_666),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_920),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_925),
.B(n_591),
.Y(n_1015)
);

OA22x2_ASAP7_75t_L g1016 ( 
.A1(n_895),
.A2(n_601),
.B1(n_612),
.B2(n_596),
.Y(n_1016)
);

OAI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_972),
.A2(n_784),
.B1(n_792),
.B2(n_741),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_923),
.A2(n_844),
.B1(n_850),
.B2(n_802),
.Y(n_1018)
);

AO22x2_ASAP7_75t_L g1019 ( 
.A1(n_945),
.A2(n_758),
.B1(n_768),
.B2(n_742),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_923),
.A2(n_853),
.B1(n_626),
.B2(n_629),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_926),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_875),
.B(n_540),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_863),
.A2(n_853),
.B1(n_634),
.B2(n_639),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_937),
.B(n_622),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_863),
.A2(n_646),
.B1(n_647),
.B2(n_645),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_885),
.A2(n_660),
.B1(n_662),
.B2(n_655),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_957),
.Y(n_1027)
);

AO22x2_ASAP7_75t_L g1028 ( 
.A1(n_934),
.A2(n_775),
.B1(n_787),
.B2(n_770),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_885),
.A2(n_676),
.B1(n_677),
.B2(n_665),
.Y(n_1029)
);

AO22x2_ASAP7_75t_L g1030 ( 
.A1(n_958),
.A2(n_788),
.B1(n_812),
.B2(n_794),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_943),
.A2(n_897),
.B1(n_886),
.B2(n_905),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_944),
.A2(n_701),
.B1(n_707),
.B2(n_681),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_922),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_893),
.A2(n_712),
.B1(n_717),
.B2(n_711),
.Y(n_1034)
);

NAND2xp33_ASAP7_75t_SL g1035 ( 
.A(n_902),
.B(n_784),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_922),
.A2(n_729),
.B1(n_733),
.B2(n_727),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_958),
.Y(n_1037)
);

AO22x2_ASAP7_75t_L g1038 ( 
.A1(n_965),
.A2(n_821),
.B1(n_841),
.B2(n_813),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_941),
.Y(n_1039)
);

OAI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_893),
.A2(n_836),
.B1(n_859),
.B2(n_792),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_941),
.B(n_799),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_868),
.A2(n_760),
.B1(n_763),
.B2(n_750),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_881),
.B(n_822),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_965),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_919),
.A2(n_765),
.B1(n_778),
.B2(n_776),
.Y(n_1045)
);

OA22x2_ASAP7_75t_L g1046 ( 
.A1(n_879),
.A2(n_930),
.B1(n_976),
.B2(n_967),
.Y(n_1046)
);

OR2x6_ASAP7_75t_L g1047 ( 
.A(n_961),
.B(n_822),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_911),
.Y(n_1048)
);

AO22x2_ASAP7_75t_L g1049 ( 
.A1(n_967),
.A2(n_976),
.B1(n_942),
.B2(n_969),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_879),
.B(n_930),
.Y(n_1050)
);

OAI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_955),
.A2(n_836),
.B1(n_783),
.B2(n_801),
.Y(n_1051)
);

OAI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_955),
.A2(n_798),
.B1(n_814),
.B2(n_804),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_884),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_938),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_949),
.A2(n_818),
.B1(n_823),
.B2(n_820),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_956),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_956),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_978),
.A2(n_825),
.B1(n_829),
.B2(n_826),
.Y(n_1058)
);

XOR2xp5_ASAP7_75t_L g1059 ( 
.A(n_864),
.B(n_830),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_913),
.A2(n_831),
.B1(n_849),
.B2(n_832),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_937),
.B(n_752),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_913),
.A2(n_571),
.B1(n_575),
.B2(n_547),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_917),
.A2(n_620),
.B1(n_627),
.B2(n_592),
.Y(n_1063)
);

NAND3x1_ASAP7_75t_L g1064 ( 
.A(n_880),
.B(n_633),
.C(n_632),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_914),
.B(n_638),
.Y(n_1065)
);

OAI22xp33_ASAP7_75t_SL g1066 ( 
.A1(n_873),
.A2(n_648),
.B1(n_649),
.B2(n_640),
.Y(n_1066)
);

OAI22xp33_ASAP7_75t_SL g1067 ( 
.A1(n_873),
.A2(n_653),
.B1(n_658),
.B2(n_650),
.Y(n_1067)
);

AO22x2_ASAP7_75t_L g1068 ( 
.A1(n_876),
.A2(n_671),
.B1(n_672),
.B2(n_661),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_964),
.B(n_539),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_956),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_948),
.Y(n_1071)
);

AND2x2_ASAP7_75t_SL g1072 ( 
.A(n_936),
.B(n_680),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_962),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_867),
.Y(n_1074)
);

OAI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_971),
.A2(n_689),
.B1(n_694),
.B2(n_683),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_917),
.A2(n_706),
.B1(n_709),
.B2(n_700),
.Y(n_1076)
);

OAI22xp33_ASAP7_75t_SL g1077 ( 
.A1(n_876),
.A2(n_722),
.B1(n_726),
.B2(n_716),
.Y(n_1077)
);

AOI22x1_ASAP7_75t_L g1078 ( 
.A1(n_977),
.A2(n_607),
.B1(n_636),
.B2(n_548),
.Y(n_1078)
);

OAI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_971),
.A2(n_740),
.B1(n_751),
.B2(n_735),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_959),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_918),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_927),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_935),
.A2(n_767),
.B1(n_774),
.B2(n_757),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_970),
.B(n_544),
.Y(n_1084)
);

INVxp67_ASAP7_75t_SL g1085 ( 
.A(n_959),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_890),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_973),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_890),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_968),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_898),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_954),
.B(n_545),
.Y(n_1091)
);

AO22x2_ASAP7_75t_L g1092 ( 
.A1(n_975),
.A2(n_782),
.B1(n_800),
.B2(n_779),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_924),
.Y(n_1093)
);

XNOR2xp5_ASAP7_75t_L g1094 ( 
.A(n_880),
.B(n_31),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_935),
.A2(n_824),
.B1(n_828),
.B2(n_819),
.Y(n_1095)
);

AO22x2_ASAP7_75t_L g1096 ( 
.A1(n_975),
.A2(n_839),
.B1(n_842),
.B2(n_835),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_924),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_898),
.Y(n_1098)
);

OR2x6_ASAP7_75t_L g1099 ( 
.A(n_901),
.B(n_845),
.Y(n_1099)
);

OAI22xp33_ASAP7_75t_SL g1100 ( 
.A1(n_929),
.A2(n_854),
.B1(n_847),
.B2(n_554),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_SL g1101 ( 
.A1(n_901),
.A2(n_548),
.B1(n_636),
.B2(n_607),
.Y(n_1101)
);

BUFx10_ASAP7_75t_L g1102 ( 
.A(n_936),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_968),
.A2(n_557),
.B1(n_562),
.B2(n_558),
.Y(n_1103)
);

AND2x2_ASAP7_75t_SL g1104 ( 
.A(n_940),
.B(n_687),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_929),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_940),
.B(n_564),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_904),
.B(n_565),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_904),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_904),
.Y(n_1109)
);

AO22x2_ASAP7_75t_L g1110 ( 
.A1(n_878),
.A2(n_687),
.B1(n_808),
.B2(n_739),
.Y(n_1110)
);

OA22x2_ASAP7_75t_L g1111 ( 
.A1(n_878),
.A2(n_699),
.B1(n_710),
.B2(n_541),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_912),
.Y(n_1112)
);

AO22x2_ASAP7_75t_L g1113 ( 
.A1(n_878),
.A2(n_808),
.B1(n_739),
.B2(n_762),
.Y(n_1113)
);

NOR2x1p5_ASAP7_75t_L g1114 ( 
.A(n_951),
.B(n_566),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_912),
.B(n_567),
.Y(n_1115)
);

NAND2xp33_ASAP7_75t_SL g1116 ( 
.A(n_951),
.B(n_568),
.Y(n_1116)
);

AOI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_878),
.A2(n_576),
.B1(n_581),
.B2(n_570),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_912),
.Y(n_1118)
);

AO22x2_ASAP7_75t_L g1119 ( 
.A1(n_910),
.A2(n_862),
.B1(n_761),
.B2(n_35),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_910),
.B(n_582),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_916),
.B(n_946),
.Y(n_1121)
);

AO22x2_ASAP7_75t_L g1122 ( 
.A1(n_910),
.A2(n_36),
.B1(n_33),
.B2(n_34),
.Y(n_1122)
);

OR2x6_ASAP7_75t_L g1123 ( 
.A(n_951),
.B(n_952),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_SL g1124 ( 
.A1(n_952),
.A2(n_588),
.B1(n_593),
.B2(n_584),
.Y(n_1124)
);

OAI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_916),
.A2(n_599),
.B1(n_603),
.B2(n_598),
.Y(n_1125)
);

INVxp67_ASAP7_75t_L g1126 ( 
.A(n_910),
.Y(n_1126)
);

AO22x2_ASAP7_75t_L g1127 ( 
.A1(n_916),
.A2(n_36),
.B1(n_33),
.B2(n_34),
.Y(n_1127)
);

OAI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_946),
.A2(n_608),
.B1(n_609),
.B2(n_605),
.Y(n_1128)
);

OAI22xp33_ASAP7_75t_SL g1129 ( 
.A1(n_946),
.A2(n_860),
.B1(n_614),
.B2(n_621),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_933),
.B(n_613),
.Y(n_1130)
);

AO22x2_ASAP7_75t_L g1131 ( 
.A1(n_933),
.A2(n_41),
.B1(n_38),
.B2(n_39),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_933),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_952),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_SL g1134 ( 
.A1(n_953),
.A2(n_624),
.B1(n_628),
.B2(n_623),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_933),
.B(n_630),
.Y(n_1135)
);

AO22x2_ASAP7_75t_L g1136 ( 
.A1(n_953),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1136)
);

AND2x2_ASAP7_75t_SL g1137 ( 
.A(n_953),
.B(n_616),
.Y(n_1137)
);

OAI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_960),
.A2(n_651),
.B1(n_654),
.B2(n_635),
.Y(n_1138)
);

OAI22xp33_ASAP7_75t_SL g1139 ( 
.A1(n_960),
.A2(n_664),
.B1(n_668),
.B2(n_663),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_960),
.A2(n_857),
.B1(n_673),
.B2(n_674),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_963),
.B(n_670),
.Y(n_1141)
);

AO22x2_ASAP7_75t_L g1142 ( 
.A1(n_963),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_963),
.B(n_682),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_966),
.B(n_690),
.Y(n_1144)
);

AO22x2_ASAP7_75t_L g1145 ( 
.A1(n_966),
.A2(n_51),
.B1(n_45),
.B2(n_49),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_966),
.B(n_691),
.Y(n_1146)
);

AO22x2_ASAP7_75t_L g1147 ( 
.A1(n_867),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_867),
.A2(n_851),
.B1(n_695),
.B2(n_696),
.Y(n_1148)
);

NAND2xp33_ASAP7_75t_SL g1149 ( 
.A(n_883),
.B(n_693),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_883),
.B(n_53),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_950),
.B(n_697),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_950),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_950),
.B(n_702),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_883),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_889),
.A2(n_718),
.B1(n_723),
.B2(n_714),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_889),
.B(n_724),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_889),
.Y(n_1157)
);

INVx1_ASAP7_75t_SL g1158 ( 
.A(n_892),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_892),
.A2(n_736),
.B1(n_737),
.B2(n_725),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_892),
.A2(n_848),
.B1(n_745),
.B2(n_747),
.Y(n_1160)
);

INVx8_ASAP7_75t_L g1161 ( 
.A(n_906),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_906),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_906),
.Y(n_1163)
);

OAI22xp33_ASAP7_75t_SL g1164 ( 
.A1(n_907),
.A2(n_748),
.B1(n_753),
.B2(n_744),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_907),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_907),
.Y(n_1166)
);

OR2x6_ASAP7_75t_L g1167 ( 
.A(n_908),
.B(n_54),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_932),
.B(n_754),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_908),
.A2(n_846),
.B1(n_756),
.B2(n_759),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_932),
.B(n_755),
.Y(n_1170)
);

NAND3x1_ASAP7_75t_L g1171 ( 
.A(n_908),
.B(n_55),
.C(n_56),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_921),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_921),
.A2(n_769),
.B1(n_771),
.B2(n_766),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_921),
.B(n_781),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_932),
.A2(n_790),
.B1(n_796),
.B2(n_793),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_869),
.B(n_797),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_869),
.B(n_803),
.Y(n_1177)
);

OAI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_928),
.A2(n_806),
.B1(n_807),
.B2(n_805),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_974),
.Y(n_1179)
);

NAND2xp33_ASAP7_75t_SL g1180 ( 
.A(n_943),
.B(n_811),
.Y(n_1180)
);

AO22x2_ASAP7_75t_L g1181 ( 
.A1(n_871),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1181)
);

AO22x2_ASAP7_75t_L g1182 ( 
.A1(n_871),
.A2(n_62),
.B1(n_58),
.B2(n_61),
.Y(n_1182)
);

OAI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_928),
.A2(n_817),
.B1(n_833),
.B2(n_816),
.Y(n_1183)
);

OA22x2_ASAP7_75t_L g1184 ( 
.A1(n_900),
.A2(n_837),
.B1(n_838),
.B2(n_834),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_894),
.A2(n_843),
.B1(n_840),
.B2(n_777),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_894),
.A2(n_777),
.B1(n_65),
.B2(n_61),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_894),
.A2(n_777),
.B1(n_66),
.B2(n_64),
.Y(n_1187)
);

AO22x2_ASAP7_75t_L g1188 ( 
.A1(n_871),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_869),
.B(n_777),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1086),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1093),
.B(n_185),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1088),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1041),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1097),
.B(n_186),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1080),
.Y(n_1195)
);

INVxp67_ASAP7_75t_SL g1196 ( 
.A(n_1105),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1044),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1104),
.B(n_187),
.Y(n_1198)
);

INVxp33_ASAP7_75t_L g1199 ( 
.A(n_1179),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1061),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_984),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_990),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_985),
.B(n_67),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1150),
.Y(n_1204)
);

NAND2xp33_ASAP7_75t_R g1205 ( 
.A(n_1089),
.B(n_1047),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_991),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1004),
.B(n_189),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1050),
.B(n_190),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1081),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1033),
.B(n_191),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_1009),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1082),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1189),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_982),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_996),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_999),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1087),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1000),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1011),
.Y(n_1219)
);

AND2x6_ASAP7_75t_L g1220 ( 
.A(n_1120),
.B(n_1007),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1014),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1039),
.B(n_193),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1021),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_979),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1075),
.B(n_194),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1028),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1028),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1079),
.B(n_196),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_998),
.B(n_202),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1030),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1030),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1047),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_986),
.B(n_69),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1053),
.B(n_206),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1038),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1038),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1027),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_994),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1048),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_994),
.Y(n_1240)
);

XOR2xp5_ASAP7_75t_L g1241 ( 
.A(n_1059),
.B(n_70),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1037),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_989),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1177),
.B(n_208),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1046),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1006),
.B(n_1015),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1049),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1013),
.B(n_70),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1049),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1126),
.A2(n_529),
.B(n_211),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1085),
.B(n_73),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1092),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1043),
.B(n_73),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1092),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1096),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1019),
.B(n_74),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1096),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1068),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1122),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_1018),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1091),
.B(n_209),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1068),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_1035),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1019),
.B(n_74),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1054),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1008),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1056),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1057),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1008),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_983),
.B(n_75),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1010),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_997),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1123),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1010),
.Y(n_1274)
);

XOR2xp5_ASAP7_75t_L g1275 ( 
.A(n_980),
.B(n_987),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1062),
.B(n_213),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_983),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1070),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1101),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1122),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1090),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1111),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1141),
.Y(n_1283)
);

XNOR2x2_ASAP7_75t_L g1284 ( 
.A(n_1147),
.B(n_75),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1098),
.Y(n_1285)
);

NAND2xp33_ASAP7_75t_R g1286 ( 
.A(n_989),
.B(n_76),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1108),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1106),
.B(n_76),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1063),
.B(n_1076),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1146),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1064),
.A2(n_526),
.B(n_218),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1065),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1001),
.Y(n_1293)
);

XOR2xp5_ASAP7_75t_L g1294 ( 
.A(n_992),
.B(n_78),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1005),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1119),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1119),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1186),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1187),
.Y(n_1299)
);

XOR2xp5_ASAP7_75t_L g1300 ( 
.A(n_1012),
.B(n_79),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1121),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1151),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1153),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1168),
.Y(n_1304)
);

AND2x6_ASAP7_75t_L g1305 ( 
.A(n_1117),
.B(n_217),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1020),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1170),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1174),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1078),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1114),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1024),
.B(n_219),
.Y(n_1311)
);

INVxp67_ASAP7_75t_SL g1312 ( 
.A(n_1110),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1110),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1042),
.B(n_79),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1167),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1055),
.B(n_1058),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1167),
.Y(n_1317)
);

INVxp33_ASAP7_75t_L g1318 ( 
.A(n_1036),
.Y(n_1318)
);

NOR2xp67_ASAP7_75t_L g1319 ( 
.A(n_1034),
.B(n_80),
.Y(n_1319)
);

NAND2xp33_ASAP7_75t_SL g1320 ( 
.A(n_1069),
.B(n_81),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1180),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1023),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1066),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1099),
.B(n_81),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1067),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1077),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1099),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1132),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1084),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1112),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1184),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1127),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1127),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1045),
.B(n_82),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1102),
.B(n_1031),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1176),
.B(n_223),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1109),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_981),
.Y(n_1338)
);

NAND2xp33_ASAP7_75t_R g1339 ( 
.A(n_1022),
.B(n_83),
.Y(n_1339)
);

INVxp33_ASAP7_75t_L g1340 ( 
.A(n_981),
.Y(n_1340)
);

INVxp33_ASAP7_75t_L g1341 ( 
.A(n_995),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1083),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1025),
.B(n_84),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1095),
.Y(n_1344)
);

INVx3_ASAP7_75t_L g1345 ( 
.A(n_1171),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1131),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1040),
.B(n_1017),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1072),
.B(n_224),
.Y(n_1348)
);

XOR2xp5_ASAP7_75t_L g1349 ( 
.A(n_1032),
.B(n_85),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1131),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1103),
.B(n_85),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1118),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_988),
.B(n_86),
.Y(n_1353)
);

INVxp33_ASAP7_75t_L g1354 ( 
.A(n_1016),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1144),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1113),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1113),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_1026),
.Y(n_1358)
);

XNOR2xp5_ASAP7_75t_L g1359 ( 
.A(n_993),
.B(n_86),
.Y(n_1359)
);

NAND2xp33_ASAP7_75t_R g1360 ( 
.A(n_1107),
.B(n_88),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1115),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1181),
.Y(n_1362)
);

XNOR2xp5_ASAP7_75t_L g1363 ( 
.A(n_1051),
.B(n_88),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1181),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1182),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1182),
.Y(n_1366)
);

BUFx5_ASAP7_75t_L g1367 ( 
.A(n_1137),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1188),
.Y(n_1368)
);

XOR2x2_ASAP7_75t_L g1369 ( 
.A(n_1100),
.B(n_89),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1188),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1071),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1073),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1156),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1139),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1164),
.Y(n_1375)
);

INVxp67_ASAP7_75t_L g1376 ( 
.A(n_1124),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1185),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1094),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1134),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1002),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1123),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1029),
.B(n_89),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1147),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1060),
.B(n_227),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1129),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1136),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1161),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1140),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1178),
.B(n_229),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1135),
.B(n_90),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1136),
.B(n_90),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1142),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1142),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1145),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1145),
.B(n_91),
.Y(n_1395)
);

NAND2xp33_ASAP7_75t_R g1396 ( 
.A(n_1003),
.B(n_91),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_1148),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1052),
.A2(n_238),
.B(n_231),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1155),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1161),
.Y(n_1400)
);

INVxp67_ASAP7_75t_SL g1401 ( 
.A(n_1130),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1183),
.B(n_242),
.Y(n_1402)
);

NAND2xp33_ASAP7_75t_R g1403 ( 
.A(n_1143),
.B(n_93),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1125),
.B(n_244),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1159),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1128),
.B(n_247),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1160),
.Y(n_1407)
);

INVxp67_ASAP7_75t_SL g1408 ( 
.A(n_1138),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1169),
.B(n_94),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1173),
.Y(n_1410)
);

XOR2x2_ASAP7_75t_L g1411 ( 
.A(n_1175),
.B(n_95),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1116),
.Y(n_1412)
);

XOR2xp5_ASAP7_75t_L g1413 ( 
.A(n_1158),
.B(n_95),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1149),
.B(n_253),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1165),
.B(n_254),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1152),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1133),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1162),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1166),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1154),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1157),
.B(n_96),
.Y(n_1421)
);

INVx4_ASAP7_75t_SL g1422 ( 
.A(n_1074),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1074),
.B(n_255),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1163),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1172),
.B(n_256),
.Y(n_1425)
);

INVxp33_ASAP7_75t_L g1426 ( 
.A(n_1179),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_985),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1086),
.Y(n_1428)
);

INVxp33_ASAP7_75t_L g1429 ( 
.A(n_1179),
.Y(n_1429)
);

XOR2xp5_ASAP7_75t_L g1430 ( 
.A(n_1059),
.B(n_98),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_985),
.B(n_99),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1086),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1086),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1086),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1086),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1086),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1093),
.B(n_259),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1150),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_985),
.B(n_99),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_SL g1440 ( 
.A(n_993),
.B(n_260),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1086),
.Y(n_1441)
);

INVxp33_ASAP7_75t_L g1442 ( 
.A(n_1179),
.Y(n_1442)
);

XOR2xp5_ASAP7_75t_L g1443 ( 
.A(n_1059),
.B(n_100),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1086),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1086),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1086),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1080),
.B(n_100),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1086),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1086),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1086),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1150),
.Y(n_1451)
);

OR2x6_ASAP7_75t_L g1452 ( 
.A(n_1047),
.B(n_101),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_985),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1150),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1086),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1086),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1150),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1093),
.B(n_261),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1093),
.B(n_263),
.Y(n_1459)
);

XOR2xp5_ASAP7_75t_L g1460 ( 
.A(n_1059),
.B(n_102),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1093),
.B(n_264),
.Y(n_1461)
);

XNOR2xp5_ASAP7_75t_L g1462 ( 
.A(n_997),
.B(n_104),
.Y(n_1462)
);

XOR2xp5_ASAP7_75t_L g1463 ( 
.A(n_1059),
.B(n_105),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1086),
.Y(n_1464)
);

INVxp33_ASAP7_75t_L g1465 ( 
.A(n_1179),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1150),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1126),
.A2(n_523),
.B(n_267),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1093),
.B(n_265),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1093),
.B(n_268),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_985),
.B(n_106),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1086),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_985),
.Y(n_1472)
);

NAND2xp33_ASAP7_75t_R g1473 ( 
.A(n_1080),
.B(n_106),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1093),
.B(n_269),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1080),
.B(n_107),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_985),
.Y(n_1476)
);

XNOR2xp5_ASAP7_75t_L g1477 ( 
.A(n_997),
.B(n_107),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1086),
.Y(n_1478)
);

XOR2xp5_ASAP7_75t_L g1479 ( 
.A(n_1059),
.B(n_109),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_985),
.B(n_109),
.Y(n_1480)
);

CKINVDCx20_ASAP7_75t_R g1481 ( 
.A(n_985),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1093),
.B(n_271),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1196),
.B(n_110),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1196),
.B(n_110),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1472),
.B(n_111),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_SL g1486 ( 
.A(n_1440),
.B(n_1472),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1427),
.B(n_1199),
.Y(n_1487)
);

OAI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1309),
.A2(n_1194),
.B(n_1191),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1273),
.Y(n_1489)
);

INVx2_ASAP7_75t_SL g1490 ( 
.A(n_1453),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1371),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1190),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1192),
.B(n_111),
.Y(n_1493)
);

AND2x2_ASAP7_75t_SL g1494 ( 
.A(n_1259),
.B(n_112),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1426),
.B(n_112),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1377),
.B(n_114),
.Y(n_1496)
);

INVxp33_ASAP7_75t_L g1497 ( 
.A(n_1429),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1428),
.B(n_115),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1432),
.B(n_115),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1372),
.Y(n_1500)
);

BUFx6f_ASAP7_75t_L g1501 ( 
.A(n_1273),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1433),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1434),
.B(n_116),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1435),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1442),
.B(n_117),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1436),
.B(n_1441),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1444),
.B(n_117),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1445),
.B(n_119),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1476),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1446),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1448),
.B(n_120),
.Y(n_1511)
);

BUFx12f_ASAP7_75t_SL g1512 ( 
.A(n_1452),
.Y(n_1512)
);

INVxp67_ASAP7_75t_L g1513 ( 
.A(n_1237),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1449),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1450),
.B(n_120),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1273),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1381),
.Y(n_1517)
);

INVx4_ASAP7_75t_L g1518 ( 
.A(n_1452),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1328),
.Y(n_1519)
);

INVxp67_ASAP7_75t_SL g1520 ( 
.A(n_1481),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1455),
.Y(n_1521)
);

OR2x6_ASAP7_75t_L g1522 ( 
.A(n_1452),
.B(n_121),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1456),
.Y(n_1523)
);

OR2x2_ASAP7_75t_SL g1524 ( 
.A(n_1347),
.B(n_121),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1464),
.B(n_123),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1471),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1478),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1197),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1465),
.B(n_124),
.Y(n_1529)
);

INVxp67_ASAP7_75t_L g1530 ( 
.A(n_1324),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1312),
.Y(n_1531)
);

INVx4_ASAP7_75t_L g1532 ( 
.A(n_1195),
.Y(n_1532)
);

INVxp67_ASAP7_75t_SL g1533 ( 
.A(n_1312),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1224),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1387),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1390),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1324),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1217),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1214),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1292),
.B(n_124),
.Y(n_1540)
);

BUFx4f_ASAP7_75t_SL g1541 ( 
.A(n_1232),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1209),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1390),
.Y(n_1543)
);

AND2x2_ASAP7_75t_SL g1544 ( 
.A(n_1440),
.B(n_126),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1203),
.B(n_127),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1246),
.B(n_127),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1212),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1200),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1201),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1202),
.B(n_128),
.Y(n_1550)
);

OAI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1191),
.A2(n_274),
.B(n_272),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1215),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1194),
.A2(n_284),
.B(n_276),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1206),
.B(n_1242),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1391),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1313),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1431),
.B(n_128),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1289),
.B(n_129),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1283),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1216),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1218),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1219),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1298),
.B(n_129),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1289),
.B(n_1327),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1221),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1290),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1247),
.B(n_130),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1299),
.B(n_130),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1470),
.B(n_131),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1480),
.B(n_131),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1439),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1437),
.A2(n_290),
.B(n_287),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1205),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1223),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1340),
.B(n_132),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1342),
.B(n_133),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1302),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1344),
.B(n_133),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1282),
.B(n_134),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1400),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1303),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1316),
.B(n_134),
.Y(n_1582)
);

OAI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1437),
.A2(n_292),
.B(n_291),
.Y(n_1583)
);

OAI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1474),
.A2(n_295),
.B(n_294),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1395),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1318),
.B(n_135),
.Y(n_1586)
);

OAI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1474),
.A2(n_300),
.B(n_296),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1304),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1267),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1351),
.B(n_135),
.Y(n_1590)
);

OAI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1482),
.A2(n_307),
.B(n_303),
.Y(n_1591)
);

OR2x6_ASAP7_75t_L g1592 ( 
.A(n_1447),
.B(n_136),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1447),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1352),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1330),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1268),
.Y(n_1596)
);

INVxp33_ASAP7_75t_L g1597 ( 
.A(n_1335),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1337),
.Y(n_1598)
);

OR2x6_ASAP7_75t_L g1599 ( 
.A(n_1475),
.B(n_137),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1307),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1308),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1351),
.B(n_138),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1323),
.B(n_139),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1325),
.B(n_1326),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1405),
.B(n_1245),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1482),
.B(n_520),
.Y(n_1606)
);

BUFx6f_ASAP7_75t_L g1607 ( 
.A(n_1278),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1249),
.B(n_139),
.Y(n_1608)
);

OAI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1458),
.A2(n_312),
.B(n_311),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1334),
.B(n_140),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1277),
.B(n_140),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1475),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1220),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1281),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1285),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1220),
.Y(n_1616)
);

INVx4_ASAP7_75t_L g1617 ( 
.A(n_1243),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1314),
.B(n_142),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1288),
.B(n_143),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1233),
.B(n_144),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1248),
.B(n_1322),
.Y(n_1621)
);

OAI21xp33_ASAP7_75t_L g1622 ( 
.A1(n_1253),
.A2(n_145),
.B(n_146),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1287),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1238),
.B(n_148),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1288),
.B(n_148),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1343),
.B(n_149),
.Y(n_1626)
);

AND2x2_ASAP7_75t_SL g1627 ( 
.A(n_1383),
.B(n_150),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1417),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1348),
.B(n_1258),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1279),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1220),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1256),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1388),
.B(n_151),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1361),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1388),
.B(n_153),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1382),
.B(n_153),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1379),
.B(n_154),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1263),
.B(n_154),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1418),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1419),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1220),
.B(n_155),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1286),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1239),
.Y(n_1643)
);

BUFx6f_ASAP7_75t_L g1644 ( 
.A(n_1345),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1301),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1348),
.B(n_1262),
.Y(n_1646)
);

BUFx5_ASAP7_75t_L g1647 ( 
.A(n_1305),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1276),
.B(n_313),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1355),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1213),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1373),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1421),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1420),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1424),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1264),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1204),
.B(n_1438),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1360),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1378),
.B(n_1275),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1265),
.Y(n_1659)
);

CKINVDCx20_ASAP7_75t_R g1660 ( 
.A(n_1397),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1263),
.B(n_155),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1276),
.B(n_314),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1265),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1459),
.A2(n_411),
.B(n_517),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1193),
.Y(n_1665)
);

INVxp67_ASAP7_75t_SL g1666 ( 
.A(n_1386),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1251),
.B(n_156),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1422),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1252),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1473),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1422),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1380),
.B(n_157),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1240),
.B(n_159),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1270),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1254),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1451),
.B(n_161),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_1345),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1422),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1454),
.Y(n_1679)
);

INVxp67_ASAP7_75t_SL g1680 ( 
.A(n_1392),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1255),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1457),
.B(n_161),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1466),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1412),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1257),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1362),
.B(n_162),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1226),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1416),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1227),
.Y(n_1689)
);

INVxp67_ASAP7_75t_SL g1690 ( 
.A(n_1393),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1261),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1394),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1230),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1261),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1461),
.A2(n_416),
.B(n_516),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1231),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1364),
.B(n_162),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1235),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1346),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1365),
.B(n_163),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1410),
.B(n_164),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1350),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1401),
.B(n_165),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1366),
.B(n_165),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1208),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1320),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1368),
.B(n_166),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1236),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1401),
.B(n_166),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1284),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1208),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1370),
.B(n_167),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1305),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1332),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1339),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1331),
.B(n_167),
.Y(n_1716)
);

BUFx3_ASAP7_75t_L g1717 ( 
.A(n_1333),
.Y(n_1717)
);

AND2x2_ASAP7_75t_SL g1718 ( 
.A(n_1280),
.B(n_168),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1293),
.B(n_168),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1266),
.B(n_169),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1269),
.Y(n_1721)
);

INVx2_ASAP7_75t_SL g1722 ( 
.A(n_1315),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1271),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1274),
.B(n_170),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1356),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1296),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1374),
.B(n_170),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1408),
.B(n_171),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1375),
.B(n_171),
.Y(n_1729)
);

AND2x2_ASAP7_75t_SL g1730 ( 
.A(n_1297),
.B(n_172),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1357),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1306),
.B(n_172),
.Y(n_1732)
);

NAND2x1p5_ASAP7_75t_L g1733 ( 
.A(n_1317),
.B(n_173),
.Y(n_1733)
);

OAI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1468),
.A2(n_426),
.B(n_514),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1338),
.B(n_174),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1305),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_1305),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1225),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1198),
.B(n_175),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1225),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1409),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1310),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1462),
.B(n_178),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1198),
.B(n_318),
.Y(n_1744)
);

NAND2x1p5_ASAP7_75t_L g1745 ( 
.A(n_1402),
.B(n_179),
.Y(n_1745)
);

NAND2x1p5_ASAP7_75t_L g1746 ( 
.A(n_1319),
.B(n_179),
.Y(n_1746)
);

AND2x2_ASAP7_75t_SL g1747 ( 
.A(n_1228),
.B(n_180),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1477),
.B(n_181),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1367),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1384),
.B(n_181),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1469),
.B(n_322),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1341),
.B(n_519),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1354),
.B(n_1329),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1228),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1398),
.B(n_323),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_SL g1756 ( 
.A(n_1398),
.B(n_1250),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1244),
.A2(n_324),
.B(n_327),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1367),
.B(n_511),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1359),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_1413),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1234),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1363),
.B(n_328),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1300),
.B(n_329),
.Y(n_1763)
);

BUFx3_ASAP7_75t_L g1764 ( 
.A(n_1321),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1353),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1353),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1423),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1369),
.B(n_333),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1358),
.B(n_507),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1385),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1425),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1367),
.B(n_338),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1294),
.B(n_501),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1367),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1376),
.B(n_340),
.Y(n_1775)
);

INVx4_ASAP7_75t_L g1776 ( 
.A(n_1367),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1207),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1403),
.Y(n_1778)
);

BUFx3_ASAP7_75t_L g1779 ( 
.A(n_1407),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1389),
.B(n_495),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1250),
.Y(n_1781)
);

INVxp67_ASAP7_75t_L g1782 ( 
.A(n_1241),
.Y(n_1782)
);

BUFx5_ASAP7_75t_L g1783 ( 
.A(n_1467),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1404),
.B(n_348),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1406),
.B(n_494),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1467),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1272),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1376),
.B(n_355),
.Y(n_1788)
);

INVx3_ASAP7_75t_SL g1789 ( 
.A(n_1411),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1430),
.B(n_356),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1349),
.Y(n_1791)
);

AND2x6_ASAP7_75t_L g1792 ( 
.A(n_1210),
.B(n_358),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1222),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_SL g1794 ( 
.A(n_1291),
.B(n_1311),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1229),
.B(n_490),
.Y(n_1795)
);

AND2x2_ASAP7_75t_SL g1796 ( 
.A(n_1414),
.B(n_1336),
.Y(n_1796)
);

INVxp67_ASAP7_75t_L g1797 ( 
.A(n_1443),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_1396),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1291),
.B(n_361),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1295),
.B(n_489),
.Y(n_1800)
);

HB1xp67_ASAP7_75t_L g1801 ( 
.A(n_1479),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1415),
.Y(n_1802)
);

NAND2x1p5_ASAP7_75t_L g1803 ( 
.A(n_1399),
.B(n_363),
.Y(n_1803)
);

INVx3_ASAP7_75t_L g1804 ( 
.A(n_1260),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1211),
.B(n_365),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1460),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1463),
.B(n_367),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1523),
.Y(n_1808)
);

OR2x6_ASAP7_75t_L g1809 ( 
.A(n_1522),
.B(n_372),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1597),
.B(n_373),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1509),
.B(n_374),
.Y(n_1811)
);

AND2x6_ASAP7_75t_L g1812 ( 
.A(n_1484),
.B(n_378),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_SL g1813 ( 
.A(n_1512),
.B(n_379),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1518),
.B(n_386),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_SL g1815 ( 
.A(n_1512),
.B(n_387),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1538),
.Y(n_1816)
);

OR2x6_ASAP7_75t_L g1817 ( 
.A(n_1522),
.B(n_388),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1523),
.B(n_389),
.Y(n_1818)
);

OR2x6_ASAP7_75t_L g1819 ( 
.A(n_1522),
.B(n_391),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1506),
.B(n_487),
.Y(n_1820)
);

CKINVDCx8_ASAP7_75t_R g1821 ( 
.A(n_1592),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1527),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1490),
.B(n_392),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1506),
.B(n_485),
.Y(n_1824)
);

AND2x2_ASAP7_75t_SL g1825 ( 
.A(n_1544),
.B(n_396),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_L g1826 ( 
.A(n_1597),
.B(n_398),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1506),
.Y(n_1827)
);

BUFx6f_ASAP7_75t_L g1828 ( 
.A(n_1501),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1621),
.B(n_399),
.Y(n_1829)
);

BUFx2_ASAP7_75t_L g1830 ( 
.A(n_1520),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1649),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_SL g1832 ( 
.A(n_1518),
.B(n_404),
.Y(n_1832)
);

OR2x6_ASAP7_75t_L g1833 ( 
.A(n_1592),
.B(n_405),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1492),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1502),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1487),
.B(n_410),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1504),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1527),
.B(n_412),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1542),
.Y(n_1839)
);

OR2x6_ASAP7_75t_L g1840 ( 
.A(n_1592),
.B(n_417),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1510),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1564),
.B(n_419),
.Y(n_1842)
);

AND2x4_ASAP7_75t_L g1843 ( 
.A(n_1651),
.B(n_484),
.Y(n_1843)
);

NAND2x1p5_ASAP7_75t_L g1844 ( 
.A(n_1501),
.B(n_421),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1543),
.B(n_483),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1632),
.B(n_424),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1514),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1787),
.B(n_425),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1564),
.B(n_428),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1501),
.Y(n_1850)
);

CKINVDCx16_ASAP7_75t_R g1851 ( 
.A(n_1599),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1658),
.B(n_429),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1558),
.B(n_430),
.Y(n_1853)
);

OR2x6_ASAP7_75t_L g1854 ( 
.A(n_1599),
.B(n_431),
.Y(n_1854)
);

INVx4_ASAP7_75t_L g1855 ( 
.A(n_1501),
.Y(n_1855)
);

OR2x6_ASAP7_75t_L g1856 ( 
.A(n_1599),
.B(n_433),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_SL g1857 ( 
.A(n_1544),
.B(n_434),
.Y(n_1857)
);

BUFx2_ASAP7_75t_L g1858 ( 
.A(n_1513),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_L g1859 ( 
.A(n_1497),
.B(n_436),
.Y(n_1859)
);

NAND2x1p5_ASAP7_75t_L g1860 ( 
.A(n_1516),
.B(n_438),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1543),
.B(n_442),
.Y(n_1861)
);

AND2x2_ASAP7_75t_SL g1862 ( 
.A(n_1494),
.B(n_444),
.Y(n_1862)
);

BUFx6f_ASAP7_75t_L g1863 ( 
.A(n_1516),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1558),
.B(n_445),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1760),
.B(n_446),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1521),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1526),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1484),
.B(n_1741),
.Y(n_1868)
);

CKINVDCx16_ASAP7_75t_R g1869 ( 
.A(n_1660),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1656),
.Y(n_1870)
);

INVx1_ASAP7_75t_SL g1871 ( 
.A(n_1541),
.Y(n_1871)
);

AND2x4_ASAP7_75t_L g1872 ( 
.A(n_1613),
.B(n_450),
.Y(n_1872)
);

BUFx12f_ASAP7_75t_L g1873 ( 
.A(n_1617),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1632),
.B(n_451),
.Y(n_1874)
);

BUFx2_ASAP7_75t_L g1875 ( 
.A(n_1484),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1679),
.B(n_453),
.Y(n_1876)
);

INVx5_ASAP7_75t_L g1877 ( 
.A(n_1516),
.Y(n_1877)
);

AND2x4_ASAP7_75t_L g1878 ( 
.A(n_1613),
.B(n_482),
.Y(n_1878)
);

INVx4_ASAP7_75t_L g1879 ( 
.A(n_1516),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1655),
.B(n_1674),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1655),
.B(n_455),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1594),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1594),
.Y(n_1883)
);

BUFx4f_ASAP7_75t_L g1884 ( 
.A(n_1803),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1497),
.B(n_456),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1674),
.B(n_457),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1547),
.Y(n_1887)
);

INVx2_ASAP7_75t_SL g1888 ( 
.A(n_1541),
.Y(n_1888)
);

BUFx24_ASAP7_75t_SL g1889 ( 
.A(n_1798),
.Y(n_1889)
);

NOR2xp67_ASAP7_75t_L g1890 ( 
.A(n_1617),
.B(n_459),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1537),
.Y(n_1891)
);

BUFx3_ASAP7_75t_L g1892 ( 
.A(n_1598),
.Y(n_1892)
);

INVx5_ASAP7_75t_L g1893 ( 
.A(n_1536),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1685),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1679),
.B(n_460),
.Y(n_1895)
);

HB1xp67_ASAP7_75t_L g1896 ( 
.A(n_1537),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1491),
.Y(n_1897)
);

BUFx2_ASAP7_75t_L g1898 ( 
.A(n_1660),
.Y(n_1898)
);

OR2x6_ASAP7_75t_L g1899 ( 
.A(n_1803),
.B(n_462),
.Y(n_1899)
);

BUFx2_ASAP7_75t_L g1900 ( 
.A(n_1498),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1685),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1616),
.B(n_463),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1491),
.Y(n_1903)
);

BUFx6f_ASAP7_75t_L g1904 ( 
.A(n_1489),
.Y(n_1904)
);

BUFx8_ASAP7_75t_L g1905 ( 
.A(n_1590),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1683),
.B(n_464),
.Y(n_1906)
);

INVx5_ASAP7_75t_L g1907 ( 
.A(n_1536),
.Y(n_1907)
);

INVx4_ASAP7_75t_L g1908 ( 
.A(n_1489),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1683),
.B(n_465),
.Y(n_1909)
);

NAND2x1p5_ASAP7_75t_L g1910 ( 
.A(n_1532),
.B(n_466),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1500),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1555),
.B(n_468),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1582),
.B(n_469),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1604),
.B(n_470),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1549),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1493),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1499),
.Y(n_1917)
);

BUFx6f_ASAP7_75t_L g1918 ( 
.A(n_1536),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1500),
.Y(n_1919)
);

AND2x6_ASAP7_75t_L g1920 ( 
.A(n_1713),
.B(n_1624),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1555),
.B(n_471),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1633),
.B(n_473),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1633),
.B(n_474),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1539),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1511),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1635),
.B(n_475),
.Y(n_1926)
);

AND2x2_ASAP7_75t_SL g1927 ( 
.A(n_1494),
.B(n_476),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1635),
.B(n_1534),
.Y(n_1928)
);

NAND2x1p5_ASAP7_75t_L g1929 ( 
.A(n_1532),
.B(n_1616),
.Y(n_1929)
);

INVx4_ASAP7_75t_L g1930 ( 
.A(n_1536),
.Y(n_1930)
);

BUFx6f_ASAP7_75t_L g1931 ( 
.A(n_1631),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1554),
.B(n_1576),
.Y(n_1932)
);

BUFx10_ASAP7_75t_L g1933 ( 
.A(n_1498),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1515),
.Y(n_1934)
);

BUFx3_ASAP7_75t_L g1935 ( 
.A(n_1598),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1578),
.B(n_1634),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1539),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1559),
.B(n_1566),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1552),
.Y(n_1939)
);

BUFx4f_ASAP7_75t_L g1940 ( 
.A(n_1746),
.Y(n_1940)
);

NAND2x1p5_ASAP7_75t_L g1941 ( 
.A(n_1631),
.B(n_1498),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1585),
.B(n_1602),
.Y(n_1942)
);

BUFx2_ASAP7_75t_L g1943 ( 
.A(n_1508),
.Y(n_1943)
);

CKINVDCx6p67_ASAP7_75t_R g1944 ( 
.A(n_1764),
.Y(n_1944)
);

INVx5_ASAP7_75t_L g1945 ( 
.A(n_1644),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1585),
.B(n_1719),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1612),
.B(n_1677),
.Y(n_1947)
);

INVx3_ASAP7_75t_L g1948 ( 
.A(n_1644),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1525),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1801),
.Y(n_1950)
);

INVx3_ASAP7_75t_L g1951 ( 
.A(n_1644),
.Y(n_1951)
);

NAND2xp33_ASAP7_75t_L g1952 ( 
.A(n_1647),
.B(n_1713),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1612),
.B(n_1677),
.Y(n_1953)
);

INVx2_ASAP7_75t_SL g1954 ( 
.A(n_1508),
.Y(n_1954)
);

BUFx2_ASAP7_75t_L g1955 ( 
.A(n_1508),
.Y(n_1955)
);

INVx4_ASAP7_75t_L g1956 ( 
.A(n_1644),
.Y(n_1956)
);

AND2x4_ASAP7_75t_L g1957 ( 
.A(n_1548),
.B(n_1530),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1715),
.B(n_1657),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1577),
.B(n_1581),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1687),
.Y(n_1960)
);

BUFx3_ASAP7_75t_L g1961 ( 
.A(n_1580),
.Y(n_1961)
);

AND2x4_ASAP7_75t_L g1962 ( 
.A(n_1689),
.B(n_1693),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1804),
.B(n_1571),
.Y(n_1963)
);

AND2x4_ASAP7_75t_L g1964 ( 
.A(n_1696),
.B(n_1698),
.Y(n_1964)
);

BUFx6f_ASAP7_75t_L g1965 ( 
.A(n_1668),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1708),
.B(n_1721),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1801),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1588),
.B(n_1600),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1601),
.B(n_1496),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1496),
.B(n_1620),
.Y(n_1970)
);

BUFx6f_ASAP7_75t_L g1971 ( 
.A(n_1668),
.Y(n_1971)
);

CKINVDCx8_ASAP7_75t_R g1972 ( 
.A(n_1713),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1586),
.B(n_1626),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1779),
.Y(n_1974)
);

INVxp67_ASAP7_75t_L g1975 ( 
.A(n_1593),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1804),
.B(n_1765),
.Y(n_1976)
);

AND2x2_ASAP7_75t_SL g1977 ( 
.A(n_1718),
.B(n_1747),
.Y(n_1977)
);

AOI21x1_ASAP7_75t_L g1978 ( 
.A1(n_1756),
.A2(n_1755),
.B(n_1794),
.Y(n_1978)
);

BUFx6f_ASAP7_75t_L g1979 ( 
.A(n_1671),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1723),
.B(n_1764),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1743),
.B(n_1748),
.Y(n_1981)
);

AND2x4_ASAP7_75t_L g1982 ( 
.A(n_1650),
.B(n_1722),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1732),
.B(n_1773),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1699),
.Y(n_1984)
);

NAND2x1p5_ASAP7_75t_L g1985 ( 
.A(n_1624),
.B(n_1673),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1766),
.B(n_1670),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1806),
.B(n_1779),
.Y(n_1987)
);

AND2x4_ASAP7_75t_L g1988 ( 
.A(n_1650),
.B(n_1645),
.Y(n_1988)
);

INVx4_ASAP7_75t_L g1989 ( 
.A(n_1624),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1586),
.B(n_1636),
.Y(n_1990)
);

INVx3_ASAP7_75t_L g1991 ( 
.A(n_1671),
.Y(n_1991)
);

NAND2xp33_ASAP7_75t_L g1992 ( 
.A(n_1647),
.B(n_1713),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1768),
.B(n_1618),
.Y(n_1993)
);

BUFx6f_ASAP7_75t_L g1994 ( 
.A(n_1678),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1495),
.B(n_1505),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1678),
.Y(n_1996)
);

INVx4_ASAP7_75t_L g1997 ( 
.A(n_1673),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1610),
.B(n_1563),
.Y(n_1998)
);

BUFx8_ASAP7_75t_L g1999 ( 
.A(n_1753),
.Y(n_1999)
);

OR2x2_ASAP7_75t_L g2000 ( 
.A(n_1806),
.B(n_1759),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1568),
.B(n_1605),
.Y(n_2001)
);

NAND2x1p5_ASAP7_75t_L g2002 ( 
.A(n_1673),
.B(n_1567),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1529),
.B(n_1670),
.Y(n_2003)
);

INVxp67_ASAP7_75t_L g2004 ( 
.A(n_1485),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1699),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1702),
.Y(n_2006)
);

AND2x4_ASAP7_75t_L g2007 ( 
.A(n_1528),
.B(n_1736),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1503),
.B(n_1507),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1800),
.B(n_1769),
.Y(n_2009)
);

INVx5_ASAP7_75t_L g2010 ( 
.A(n_1567),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1702),
.Y(n_2011)
);

INVx5_ASAP7_75t_L g2012 ( 
.A(n_1567),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1789),
.B(n_1762),
.Y(n_2013)
);

INVx4_ASAP7_75t_L g2014 ( 
.A(n_1580),
.Y(n_2014)
);

NOR2x1_ASAP7_75t_L g2015 ( 
.A(n_1736),
.B(n_1737),
.Y(n_2015)
);

INVx5_ASAP7_75t_L g2016 ( 
.A(n_1737),
.Y(n_2016)
);

INVxp67_ASAP7_75t_SL g2017 ( 
.A(n_1531),
.Y(n_2017)
);

INVxp67_ASAP7_75t_SL g2018 ( 
.A(n_1531),
.Y(n_2018)
);

INVx6_ASAP7_75t_SL g2019 ( 
.A(n_1524),
.Y(n_2019)
);

CKINVDCx20_ASAP7_75t_R g2020 ( 
.A(n_1573),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1503),
.B(n_1507),
.Y(n_2021)
);

BUFx12f_ASAP7_75t_L g2022 ( 
.A(n_1746),
.Y(n_2022)
);

AND2x4_ASAP7_75t_L g2023 ( 
.A(n_1706),
.B(n_1517),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_L g2024 ( 
.A(n_1778),
.B(n_1642),
.Y(n_2024)
);

OR2x6_ASAP7_75t_SL g2025 ( 
.A(n_1763),
.B(n_1790),
.Y(n_2025)
);

BUFx2_ASAP7_75t_L g2026 ( 
.A(n_1778),
.Y(n_2026)
);

INVx2_ASAP7_75t_SL g2027 ( 
.A(n_1733),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1552),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1560),
.Y(n_2029)
);

BUFx4f_ASAP7_75t_L g2030 ( 
.A(n_1733),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1560),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1561),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1561),
.Y(n_2033)
);

NOR2xp33_ASAP7_75t_L g2034 ( 
.A(n_1517),
.B(n_1770),
.Y(n_2034)
);

INVx4_ASAP7_75t_L g2035 ( 
.A(n_1718),
.Y(n_2035)
);

INVx4_ASAP7_75t_L g2036 ( 
.A(n_1627),
.Y(n_2036)
);

BUFx2_ASAP7_75t_L g2037 ( 
.A(n_1533),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1562),
.Y(n_2038)
);

NAND2x1_ASAP7_75t_SL g2039 ( 
.A(n_1710),
.B(n_1775),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_1726),
.B(n_1714),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1789),
.B(n_1730),
.Y(n_2041)
);

AND2x6_ASAP7_75t_L g2042 ( 
.A(n_1714),
.B(n_1717),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1562),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1747),
.B(n_1705),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1728),
.B(n_1652),
.Y(n_2045)
);

NOR2xp33_ASAP7_75t_L g2046 ( 
.A(n_1535),
.B(n_1665),
.Y(n_2046)
);

OR2x6_ASAP7_75t_L g2047 ( 
.A(n_1710),
.B(n_1782),
.Y(n_2047)
);

AND2x6_ASAP7_75t_L g2048 ( 
.A(n_1717),
.B(n_1556),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1565),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1565),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1574),
.Y(n_2051)
);

AND2x2_ASAP7_75t_SL g2052 ( 
.A(n_1730),
.B(n_1627),
.Y(n_2052)
);

HB1xp67_ASAP7_75t_L g2053 ( 
.A(n_1574),
.Y(n_2053)
);

INVx1_ASAP7_75t_SL g2054 ( 
.A(n_1575),
.Y(n_2054)
);

OR2x2_ASAP7_75t_L g2055 ( 
.A(n_1791),
.B(n_1797),
.Y(n_2055)
);

BUFx2_ASAP7_75t_L g2056 ( 
.A(n_1483),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1692),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_1791),
.Y(n_2058)
);

INVxp67_ASAP7_75t_L g2059 ( 
.A(n_1667),
.Y(n_2059)
);

AND2x4_ASAP7_75t_L g2060 ( 
.A(n_1669),
.B(n_1675),
.Y(n_2060)
);

INVx1_ASAP7_75t_SL g2061 ( 
.A(n_1686),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1637),
.B(n_1603),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1637),
.B(n_1652),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1628),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1807),
.B(n_1545),
.Y(n_2065)
);

INVx2_ASAP7_75t_SL g2066 ( 
.A(n_1697),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1728),
.B(n_1672),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1628),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1672),
.B(n_1738),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1807),
.B(n_1557),
.Y(n_2070)
);

OR2x6_ASAP7_75t_L g2071 ( 
.A(n_1805),
.B(n_1619),
.Y(n_2071)
);

AND2x4_ASAP7_75t_L g2072 ( 
.A(n_1681),
.B(n_1608),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1738),
.B(n_1740),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1692),
.Y(n_2074)
);

OR2x6_ASAP7_75t_L g2075 ( 
.A(n_1625),
.B(n_1752),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1639),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1569),
.B(n_1570),
.Y(n_2077)
);

INVx1_ASAP7_75t_SL g2078 ( 
.A(n_1700),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1639),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_1540),
.B(n_1546),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1704),
.B(n_1707),
.Y(n_2081)
);

AND2x4_ASAP7_75t_L g2082 ( 
.A(n_1712),
.B(n_1611),
.Y(n_2082)
);

NAND2x1p5_ASAP7_75t_L g2083 ( 
.A(n_1535),
.B(n_1776),
.Y(n_2083)
);

BUFx12f_ASAP7_75t_L g2084 ( 
.A(n_1735),
.Y(n_2084)
);

OR2x6_ASAP7_75t_L g2085 ( 
.A(n_1788),
.B(n_1745),
.Y(n_2085)
);

BUFx2_ASAP7_75t_L g2086 ( 
.A(n_1703),
.Y(n_2086)
);

AND2x4_ASAP7_75t_L g2087 ( 
.A(n_1688),
.B(n_1776),
.Y(n_2087)
);

HB1xp67_ASAP7_75t_L g2088 ( 
.A(n_1709),
.Y(n_2088)
);

BUFx3_ASAP7_75t_L g2089 ( 
.A(n_1742),
.Y(n_2089)
);

NOR2x1_ASAP7_75t_L g2090 ( 
.A(n_1641),
.B(n_1720),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1638),
.B(n_1661),
.Y(n_2091)
);

INVx5_ASAP7_75t_L g2092 ( 
.A(n_1589),
.Y(n_2092)
);

BUFx3_ASAP7_75t_L g2093 ( 
.A(n_1643),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1740),
.B(n_1754),
.Y(n_2094)
);

BUFx8_ASAP7_75t_L g2095 ( 
.A(n_1647),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1640),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1754),
.B(n_1727),
.Y(n_2097)
);

INVx4_ASAP7_75t_L g2098 ( 
.A(n_1589),
.Y(n_2098)
);

OR2x6_ASAP7_75t_L g2099 ( 
.A(n_1745),
.B(n_1724),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_1595),
.B(n_1729),
.Y(n_2100)
);

INVx1_ASAP7_75t_SL g2101 ( 
.A(n_1676),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1640),
.Y(n_2102)
);

BUFx4f_ASAP7_75t_L g2103 ( 
.A(n_1684),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1750),
.B(n_1682),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_SL g2105 ( 
.A(n_1647),
.B(n_1622),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1666),
.B(n_1680),
.Y(n_2106)
);

INVx5_ASAP7_75t_L g2107 ( 
.A(n_1589),
.Y(n_2107)
);

NOR2xp67_ASAP7_75t_L g2108 ( 
.A(n_1716),
.B(n_1579),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1690),
.B(n_1629),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1725),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1550),
.Y(n_2111)
);

NOR2xp33_ASAP7_75t_L g2112 ( 
.A(n_1629),
.B(n_1646),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_1595),
.B(n_1643),
.Y(n_2113)
);

HB1xp67_ASAP7_75t_L g2114 ( 
.A(n_1596),
.Y(n_2114)
);

INVxp67_ASAP7_75t_SL g2115 ( 
.A(n_1705),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_1688),
.B(n_1725),
.Y(n_2116)
);

AND2x4_ASAP7_75t_L g2117 ( 
.A(n_1731),
.B(n_1684),
.Y(n_2117)
);

NAND2x1p5_ASAP7_75t_L g2118 ( 
.A(n_1659),
.B(n_1663),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1731),
.Y(n_2119)
);

BUFx2_ASAP7_75t_L g2120 ( 
.A(n_1647),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1556),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1646),
.B(n_1711),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1701),
.Y(n_2123)
);

AND2x4_ASAP7_75t_L g2124 ( 
.A(n_1749),
.B(n_1659),
.Y(n_2124)
);

BUFx3_ASAP7_75t_L g2125 ( 
.A(n_1663),
.Y(n_2125)
);

HB1xp67_ASAP7_75t_L g2126 ( 
.A(n_1614),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_1615),
.B(n_1623),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1615),
.Y(n_2128)
);

NAND2x1p5_ASAP7_75t_L g2129 ( 
.A(n_1623),
.B(n_1589),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1630),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_1774),
.B(n_1711),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1653),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2133)
);

OR2x2_ASAP7_75t_L g2134 ( 
.A(n_1739),
.B(n_1654),
.Y(n_2134)
);

BUFx12f_ASAP7_75t_L g2135 ( 
.A(n_1607),
.Y(n_2135)
);

OR2x6_ASAP7_75t_L g2136 ( 
.A(n_1486),
.B(n_1757),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_SL g2137 ( 
.A(n_1647),
.B(n_1691),
.Y(n_2137)
);

AND2x4_ASAP7_75t_L g2138 ( 
.A(n_1694),
.B(n_1486),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1781),
.B(n_1786),
.Y(n_2139)
);

NOR2xp33_ASAP7_75t_L g2140 ( 
.A(n_1796),
.B(n_1777),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1781),
.B(n_1786),
.Y(n_2141)
);

NOR2xp33_ASAP7_75t_L g2142 ( 
.A(n_1796),
.B(n_1780),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_SL g2143 ( 
.A(n_1607),
.B(n_1519),
.Y(n_2143)
);

INVx4_ASAP7_75t_L g2144 ( 
.A(n_1519),
.Y(n_2144)
);

AND2x6_ASAP7_75t_L g2145 ( 
.A(n_1761),
.B(n_1784),
.Y(n_2145)
);

BUFx8_ASAP7_75t_SL g2146 ( 
.A(n_1653),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_SL g2147 ( 
.A(n_1802),
.B(n_1793),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_1654),
.B(n_1785),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1756),
.B(n_1783),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1783),
.B(n_1802),
.Y(n_2150)
);

INVx1_ASAP7_75t_SL g2151 ( 
.A(n_1648),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1648),
.Y(n_2152)
);

CKINVDCx8_ASAP7_75t_R g2153 ( 
.A(n_1851),
.Y(n_2153)
);

NOR2x1_ASAP7_75t_SL g2154 ( 
.A(n_1833),
.B(n_1840),
.Y(n_2154)
);

INVx5_ASAP7_75t_L g2155 ( 
.A(n_1809),
.Y(n_2155)
);

INVx3_ASAP7_75t_L g2156 ( 
.A(n_2135),
.Y(n_2156)
);

INVx3_ASAP7_75t_L g2157 ( 
.A(n_1893),
.Y(n_2157)
);

INVx2_ASAP7_75t_SL g2158 ( 
.A(n_1884),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1839),
.B(n_1783),
.Y(n_2159)
);

BUFx3_ASAP7_75t_L g2160 ( 
.A(n_2146),
.Y(n_2160)
);

CKINVDCx11_ASAP7_75t_R g2161 ( 
.A(n_1821),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1839),
.B(n_1783),
.Y(n_2162)
);

NAND2x1p5_ASAP7_75t_L g2163 ( 
.A(n_2010),
.B(n_1755),
.Y(n_2163)
);

BUFx3_ASAP7_75t_L g2164 ( 
.A(n_1873),
.Y(n_2164)
);

BUFx4_ASAP7_75t_SL g2165 ( 
.A(n_1809),
.Y(n_2165)
);

BUFx6f_ASAP7_75t_L g2166 ( 
.A(n_1828),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1938),
.Y(n_2167)
);

BUFx8_ASAP7_75t_L g2168 ( 
.A(n_1898),
.Y(n_2168)
);

BUFx4_ASAP7_75t_SL g2169 ( 
.A(n_1817),
.Y(n_2169)
);

INVx4_ASAP7_75t_L g2170 ( 
.A(n_1817),
.Y(n_2170)
);

BUFx3_ASAP7_75t_L g2171 ( 
.A(n_1892),
.Y(n_2171)
);

BUFx12f_ASAP7_75t_L g2172 ( 
.A(n_1888),
.Y(n_2172)
);

INVx1_ASAP7_75t_SL g2173 ( 
.A(n_2037),
.Y(n_2173)
);

NAND2x1p5_ASAP7_75t_L g2174 ( 
.A(n_2010),
.B(n_1662),
.Y(n_2174)
);

BUFx6f_ASAP7_75t_L g2175 ( 
.A(n_1828),
.Y(n_2175)
);

BUFx2_ASAP7_75t_L g2176 ( 
.A(n_1819),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1870),
.B(n_1783),
.Y(n_2177)
);

BUFx3_ASAP7_75t_L g2178 ( 
.A(n_1935),
.Y(n_2178)
);

INVx3_ASAP7_75t_L g2179 ( 
.A(n_1893),
.Y(n_2179)
);

INVx2_ASAP7_75t_SL g2180 ( 
.A(n_2030),
.Y(n_2180)
);

BUFx12f_ASAP7_75t_L g2181 ( 
.A(n_1816),
.Y(n_2181)
);

BUFx8_ASAP7_75t_L g2182 ( 
.A(n_2022),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1993),
.B(n_1662),
.Y(n_2183)
);

INVx5_ASAP7_75t_L g2184 ( 
.A(n_1819),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1959),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_1981),
.B(n_1783),
.Y(n_2186)
);

BUFx4_ASAP7_75t_SL g2187 ( 
.A(n_1833),
.Y(n_2187)
);

BUFx8_ASAP7_75t_L g2188 ( 
.A(n_1830),
.Y(n_2188)
);

BUFx24_ASAP7_75t_L g2189 ( 
.A(n_1845),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2052),
.B(n_1793),
.Y(n_2190)
);

BUFx2_ASAP7_75t_L g2191 ( 
.A(n_1840),
.Y(n_2191)
);

INVx1_ASAP7_75t_SL g2192 ( 
.A(n_1985),
.Y(n_2192)
);

NOR2xp33_ASAP7_75t_L g2193 ( 
.A(n_2130),
.B(n_1794),
.Y(n_2193)
);

BUFx2_ASAP7_75t_L g2194 ( 
.A(n_1854),
.Y(n_2194)
);

CKINVDCx14_ASAP7_75t_R g2195 ( 
.A(n_1854),
.Y(n_2195)
);

HB1xp67_ASAP7_75t_L g2196 ( 
.A(n_2002),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1968),
.Y(n_2197)
);

INVx3_ASAP7_75t_L g2198 ( 
.A(n_1893),
.Y(n_2198)
);

INVx3_ASAP7_75t_L g2199 ( 
.A(n_1907),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2028),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1831),
.Y(n_2201)
);

INVxp67_ASAP7_75t_SL g2202 ( 
.A(n_1941),
.Y(n_2202)
);

BUFx6f_ASAP7_75t_L g2203 ( 
.A(n_1828),
.Y(n_2203)
);

INVx2_ASAP7_75t_SL g2204 ( 
.A(n_2103),
.Y(n_2204)
);

INVx1_ASAP7_75t_SL g2205 ( 
.A(n_1933),
.Y(n_2205)
);

INVx1_ASAP7_75t_SL g2206 ( 
.A(n_1933),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_1946),
.B(n_1584),
.Y(n_2207)
);

INVx4_ASAP7_75t_L g2208 ( 
.A(n_1856),
.Y(n_2208)
);

BUFx3_ASAP7_75t_L g2209 ( 
.A(n_1944),
.Y(n_2209)
);

BUFx3_ASAP7_75t_L g2210 ( 
.A(n_1871),
.Y(n_2210)
);

INVx5_ASAP7_75t_L g2211 ( 
.A(n_1856),
.Y(n_2211)
);

INVx6_ASAP7_75t_SL g2212 ( 
.A(n_1899),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1834),
.Y(n_2213)
);

BUFx3_ASAP7_75t_L g2214 ( 
.A(n_1858),
.Y(n_2214)
);

BUFx2_ASAP7_75t_SL g2215 ( 
.A(n_1907),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1835),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1837),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2028),
.Y(n_2218)
);

INVx5_ASAP7_75t_L g2219 ( 
.A(n_1812),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1841),
.Y(n_2220)
);

INVx4_ASAP7_75t_L g2221 ( 
.A(n_1907),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_1942),
.B(n_1983),
.Y(n_2222)
);

INVx1_ASAP7_75t_SL g2223 ( 
.A(n_2087),
.Y(n_2223)
);

INVx5_ASAP7_75t_SL g2224 ( 
.A(n_1899),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1847),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1866),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1867),
.Y(n_2227)
);

BUFx12f_ASAP7_75t_L g2228 ( 
.A(n_1974),
.Y(n_2228)
);

CKINVDCx20_ASAP7_75t_R g2229 ( 
.A(n_1869),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1977),
.B(n_1587),
.Y(n_2230)
);

NAND2x1p5_ASAP7_75t_L g2231 ( 
.A(n_2010),
.B(n_1744),
.Y(n_2231)
);

BUFx3_ASAP7_75t_L g2232 ( 
.A(n_1999),
.Y(n_2232)
);

BUFx10_ASAP7_75t_L g2233 ( 
.A(n_1845),
.Y(n_2233)
);

BUFx2_ASAP7_75t_L g2234 ( 
.A(n_1861),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_2029),
.Y(n_2235)
);

INVx1_ASAP7_75t_SL g2236 ( 
.A(n_2087),
.Y(n_2236)
);

INVx3_ASAP7_75t_L g2237 ( 
.A(n_1972),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_2029),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1887),
.Y(n_2239)
);

INVxp67_ASAP7_75t_SL g2240 ( 
.A(n_1875),
.Y(n_2240)
);

INVxp67_ASAP7_75t_SL g2241 ( 
.A(n_2053),
.Y(n_2241)
);

INVx1_ASAP7_75t_SL g2242 ( 
.A(n_1820),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1915),
.Y(n_2243)
);

NAND2x1p5_ASAP7_75t_L g2244 ( 
.A(n_2012),
.B(n_1744),
.Y(n_2244)
);

BUFx6f_ASAP7_75t_L g2245 ( 
.A(n_1850),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_2043),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2009),
.B(n_1583),
.Y(n_2247)
);

INVx1_ASAP7_75t_SL g2248 ( 
.A(n_1820),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2043),
.Y(n_2249)
);

BUFx2_ASAP7_75t_SL g2250 ( 
.A(n_1861),
.Y(n_2250)
);

OR2x2_ASAP7_75t_L g2251 ( 
.A(n_2000),
.B(n_1799),
.Y(n_2251)
);

BUFx3_ASAP7_75t_L g2252 ( 
.A(n_1999),
.Y(n_2252)
);

BUFx3_ASAP7_75t_L g2253 ( 
.A(n_1961),
.Y(n_2253)
);

INVx3_ASAP7_75t_L g2254 ( 
.A(n_1930),
.Y(n_2254)
);

AND2x4_ASAP7_75t_L g2255 ( 
.A(n_1824),
.B(n_1591),
.Y(n_2255)
);

CKINVDCx8_ASAP7_75t_R g2256 ( 
.A(n_1950),
.Y(n_2256)
);

BUFx3_ASAP7_75t_L g2257 ( 
.A(n_1940),
.Y(n_2257)
);

CKINVDCx11_ASAP7_75t_R g2258 ( 
.A(n_2025),
.Y(n_2258)
);

BUFx6f_ASAP7_75t_L g2259 ( 
.A(n_1863),
.Y(n_2259)
);

BUFx2_ASAP7_75t_L g2260 ( 
.A(n_1812),
.Y(n_2260)
);

BUFx6f_ASAP7_75t_L g2261 ( 
.A(n_1863),
.Y(n_2261)
);

NAND2x1p5_ASAP7_75t_L g2262 ( 
.A(n_2012),
.B(n_1606),
.Y(n_2262)
);

INVx1_ASAP7_75t_SL g2263 ( 
.A(n_1824),
.Y(n_2263)
);

INVx1_ASAP7_75t_SL g2264 ( 
.A(n_1900),
.Y(n_2264)
);

CKINVDCx16_ASAP7_75t_R g2265 ( 
.A(n_1813),
.Y(n_2265)
);

AOI22xp5_ASAP7_75t_L g2266 ( 
.A1(n_1862),
.A2(n_1792),
.B1(n_1771),
.B2(n_1606),
.Y(n_2266)
);

BUFx3_ASAP7_75t_L g2267 ( 
.A(n_1905),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1960),
.Y(n_2268)
);

INVx3_ASAP7_75t_SL g2269 ( 
.A(n_1927),
.Y(n_2269)
);

BUFx2_ASAP7_75t_L g2270 ( 
.A(n_1812),
.Y(n_2270)
);

BUFx2_ASAP7_75t_L g2271 ( 
.A(n_1812),
.Y(n_2271)
);

BUFx3_ASAP7_75t_L g2272 ( 
.A(n_1905),
.Y(n_2272)
);

INVx5_ASAP7_75t_L g2273 ( 
.A(n_2042),
.Y(n_2273)
);

INVx1_ASAP7_75t_SL g2274 ( 
.A(n_1943),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_1808),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1960),
.Y(n_2276)
);

NAND2x1p5_ASAP7_75t_L g2277 ( 
.A(n_2012),
.B(n_1761),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_1808),
.Y(n_2278)
);

NAND2x1p5_ASAP7_75t_L g2279 ( 
.A(n_1989),
.B(n_1761),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1822),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1894),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1894),
.Y(n_2282)
);

INVx4_ASAP7_75t_L g2283 ( 
.A(n_1877),
.Y(n_2283)
);

CKINVDCx16_ASAP7_75t_R g2284 ( 
.A(n_1815),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2133),
.B(n_1488),
.Y(n_2285)
);

BUFx6f_ASAP7_75t_L g2286 ( 
.A(n_1863),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1901),
.Y(n_2287)
);

BUFx6f_ASAP7_75t_L g2288 ( 
.A(n_1877),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_1822),
.Y(n_2289)
);

BUFx3_ASAP7_75t_L g2290 ( 
.A(n_1918),
.Y(n_2290)
);

INVx5_ASAP7_75t_L g2291 ( 
.A(n_2042),
.Y(n_2291)
);

INVx3_ASAP7_75t_SL g2292 ( 
.A(n_1825),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1901),
.Y(n_2293)
);

NAND2x1p5_ASAP7_75t_L g2294 ( 
.A(n_1989),
.B(n_1761),
.Y(n_2294)
);

BUFx3_ASAP7_75t_L g2295 ( 
.A(n_1918),
.Y(n_2295)
);

INVx1_ASAP7_75t_SL g2296 ( 
.A(n_1955),
.Y(n_2296)
);

CKINVDCx20_ASAP7_75t_R g2297 ( 
.A(n_2020),
.Y(n_2297)
);

BUFx3_ASAP7_75t_L g2298 ( 
.A(n_1918),
.Y(n_2298)
);

INVx4_ASAP7_75t_L g2299 ( 
.A(n_1877),
.Y(n_2299)
);

BUFx12f_ASAP7_75t_L g2300 ( 
.A(n_1967),
.Y(n_2300)
);

BUFx3_ASAP7_75t_L g2301 ( 
.A(n_1988),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_1882),
.Y(n_2302)
);

AOI22xp33_ASAP7_75t_L g2303 ( 
.A1(n_2019),
.A2(n_1792),
.B1(n_1771),
.B2(n_1767),
.Y(n_2303)
);

NAND2x1p5_ASAP7_75t_L g2304 ( 
.A(n_1997),
.B(n_1945),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1984),
.Y(n_2305)
);

BUFx4f_ASAP7_75t_SL g2306 ( 
.A(n_2019),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_1883),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2064),
.Y(n_2308)
);

AOI22xp33_ASAP7_75t_L g2309 ( 
.A1(n_2035),
.A2(n_1792),
.B1(n_1767),
.B2(n_1734),
.Y(n_2309)
);

BUFx3_ASAP7_75t_L g2310 ( 
.A(n_1988),
.Y(n_2310)
);

BUFx12f_ASAP7_75t_L g2311 ( 
.A(n_2058),
.Y(n_2311)
);

BUFx2_ASAP7_75t_L g2312 ( 
.A(n_1920),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2068),
.Y(n_2313)
);

INVx3_ASAP7_75t_L g2314 ( 
.A(n_1930),
.Y(n_2314)
);

HB1xp67_ASAP7_75t_L g2315 ( 
.A(n_2114),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2076),
.Y(n_2316)
);

HB1xp67_ASAP7_75t_L g2317 ( 
.A(n_2126),
.Y(n_2317)
);

NAND2x1p5_ASAP7_75t_L g2318 ( 
.A(n_1997),
.B(n_1772),
.Y(n_2318)
);

BUFx2_ASAP7_75t_L g2319 ( 
.A(n_1920),
.Y(n_2319)
);

CKINVDCx20_ASAP7_75t_R g2320 ( 
.A(n_2095),
.Y(n_2320)
);

INVx3_ASAP7_75t_SL g2321 ( 
.A(n_2047),
.Y(n_2321)
);

INVx6_ASAP7_75t_SL g2322 ( 
.A(n_2047),
.Y(n_2322)
);

INVx5_ASAP7_75t_L g2323 ( 
.A(n_2042),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2079),
.Y(n_2324)
);

INVx1_ASAP7_75t_SL g2325 ( 
.A(n_2113),
.Y(n_2325)
);

INVxp67_ASAP7_75t_SL g2326 ( 
.A(n_2115),
.Y(n_2326)
);

INVx1_ASAP7_75t_SL g2327 ( 
.A(n_2093),
.Y(n_2327)
);

INVx2_ASAP7_75t_SL g2328 ( 
.A(n_1982),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2065),
.B(n_1551),
.Y(n_2329)
);

BUFx3_ASAP7_75t_L g2330 ( 
.A(n_1929),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2070),
.B(n_1553),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2067),
.B(n_1792),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1984),
.Y(n_2333)
);

BUFx12f_ASAP7_75t_L g2334 ( 
.A(n_1987),
.Y(n_2334)
);

BUFx3_ASAP7_75t_L g2335 ( 
.A(n_1982),
.Y(n_2335)
);

CKINVDCx16_ASAP7_75t_R g2336 ( 
.A(n_1832),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2005),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2005),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2096),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2006),
.Y(n_2340)
);

INVx6_ASAP7_75t_L g2341 ( 
.A(n_2084),
.Y(n_2341)
);

INVx3_ASAP7_75t_L g2342 ( 
.A(n_2042),
.Y(n_2342)
);

BUFx3_ASAP7_75t_L g2343 ( 
.A(n_1904),
.Y(n_2343)
);

BUFx12f_ASAP7_75t_L g2344 ( 
.A(n_2055),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2140),
.B(n_1792),
.Y(n_2345)
);

INVx4_ASAP7_75t_L g2346 ( 
.A(n_1945),
.Y(n_2346)
);

BUFx2_ASAP7_75t_L g2347 ( 
.A(n_1920),
.Y(n_2347)
);

BUFx5_ASAP7_75t_L g2348 ( 
.A(n_2048),
.Y(n_2348)
);

INVx4_ASAP7_75t_L g2349 ( 
.A(n_1945),
.Y(n_2349)
);

BUFx10_ASAP7_75t_L g2350 ( 
.A(n_2027),
.Y(n_2350)
);

INVx4_ASAP7_75t_L g2351 ( 
.A(n_1920),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2102),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_1897),
.Y(n_2353)
);

BUFx3_ASAP7_75t_L g2354 ( 
.A(n_1904),
.Y(n_2354)
);

INVx3_ASAP7_75t_L g2355 ( 
.A(n_1931),
.Y(n_2355)
);

BUFx3_ASAP7_75t_L g2356 ( 
.A(n_1904),
.Y(n_2356)
);

BUFx8_ASAP7_75t_L g2357 ( 
.A(n_2026),
.Y(n_2357)
);

CKINVDCx8_ASAP7_75t_R g2358 ( 
.A(n_1980),
.Y(n_2358)
);

INVx4_ASAP7_75t_L g2359 ( 
.A(n_2092),
.Y(n_2359)
);

BUFx2_ASAP7_75t_L g2360 ( 
.A(n_2035),
.Y(n_2360)
);

BUFx3_ASAP7_75t_L g2361 ( 
.A(n_2089),
.Y(n_2361)
);

OR2x6_ASAP7_75t_L g2362 ( 
.A(n_2036),
.B(n_1572),
.Y(n_2362)
);

BUFx3_ASAP7_75t_L g2363 ( 
.A(n_1980),
.Y(n_2363)
);

NOR2xp33_ASAP7_75t_L g2364 ( 
.A(n_1970),
.B(n_1758),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_1880),
.B(n_1609),
.Y(n_2365)
);

CKINVDCx11_ASAP7_75t_R g2366 ( 
.A(n_1889),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_1903),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_1911),
.Y(n_2368)
);

BUFx5_ASAP7_75t_L g2369 ( 
.A(n_2048),
.Y(n_2369)
);

BUFx3_ASAP7_75t_L g2370 ( 
.A(n_2083),
.Y(n_2370)
);

NAND2x1p5_ASAP7_75t_L g2371 ( 
.A(n_2092),
.B(n_1751),
.Y(n_2371)
);

BUFx3_ASAP7_75t_L g2372 ( 
.A(n_1931),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2041),
.B(n_1664),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_1919),
.Y(n_2374)
);

AOI22xp33_ASAP7_75t_L g2375 ( 
.A1(n_2036),
.A2(n_1695),
.B1(n_1795),
.B2(n_2062),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2006),
.Y(n_2376)
);

INVx4_ASAP7_75t_SL g2377 ( 
.A(n_2048),
.Y(n_2377)
);

BUFx3_ASAP7_75t_L g2378 ( 
.A(n_1931),
.Y(n_2378)
);

BUFx12f_ASAP7_75t_L g2379 ( 
.A(n_2095),
.Y(n_2379)
);

INVx6_ASAP7_75t_L g2380 ( 
.A(n_2014),
.Y(n_2380)
);

INVx4_ASAP7_75t_L g2381 ( 
.A(n_2092),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_1924),
.Y(n_2382)
);

BUFx3_ASAP7_75t_L g2383 ( 
.A(n_2034),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_1937),
.Y(n_2384)
);

BUFx24_ASAP7_75t_L g2385 ( 
.A(n_1872),
.Y(n_2385)
);

INVx1_ASAP7_75t_SL g2386 ( 
.A(n_2127),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2011),
.Y(n_2387)
);

BUFx2_ASAP7_75t_SL g2388 ( 
.A(n_1890),
.Y(n_2388)
);

INVx5_ASAP7_75t_L g2389 ( 
.A(n_2048),
.Y(n_2389)
);

BUFx24_ASAP7_75t_L g2390 ( 
.A(n_1872),
.Y(n_2390)
);

BUFx3_ASAP7_75t_L g2391 ( 
.A(n_2014),
.Y(n_2391)
);

CKINVDCx5p33_ASAP7_75t_R g2392 ( 
.A(n_1963),
.Y(n_2392)
);

INVx1_ASAP7_75t_SL g2393 ( 
.A(n_1891),
.Y(n_2393)
);

BUFx2_ASAP7_75t_SL g2394 ( 
.A(n_1878),
.Y(n_2394)
);

BUFx3_ASAP7_75t_L g2395 ( 
.A(n_1908),
.Y(n_2395)
);

INVx5_ASAP7_75t_L g2396 ( 
.A(n_1855),
.Y(n_2396)
);

BUFx6f_ASAP7_75t_L g2397 ( 
.A(n_2107),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_1939),
.Y(n_2398)
);

INVx2_ASAP7_75t_SL g2399 ( 
.A(n_1957),
.Y(n_2399)
);

INVx4_ASAP7_75t_L g2400 ( 
.A(n_2107),
.Y(n_2400)
);

BUFx4f_ASAP7_75t_SL g2401 ( 
.A(n_1908),
.Y(n_2401)
);

BUFx6f_ASAP7_75t_L g2402 ( 
.A(n_2107),
.Y(n_2402)
);

OAI22xp5_ASAP7_75t_SL g2403 ( 
.A1(n_1969),
.A2(n_1928),
.B1(n_1868),
.B2(n_1976),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2011),
.Y(n_2404)
);

BUFx8_ASAP7_75t_L g2405 ( 
.A(n_2013),
.Y(n_2405)
);

BUFx3_ASAP7_75t_L g2406 ( 
.A(n_2023),
.Y(n_2406)
);

INVx4_ASAP7_75t_L g2407 ( 
.A(n_1855),
.Y(n_2407)
);

INVx3_ASAP7_75t_L g2408 ( 
.A(n_1956),
.Y(n_2408)
);

INVx3_ASAP7_75t_L g2409 ( 
.A(n_1956),
.Y(n_2409)
);

INVx2_ASAP7_75t_SL g2410 ( 
.A(n_1957),
.Y(n_2410)
);

OR2x6_ASAP7_75t_SL g2411 ( 
.A(n_1852),
.B(n_1865),
.Y(n_2411)
);

BUFx3_ASAP7_75t_L g2412 ( 
.A(n_2023),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2057),
.Y(n_2413)
);

INVx4_ASAP7_75t_L g2414 ( 
.A(n_1879),
.Y(n_2414)
);

AOI22xp33_ASAP7_75t_L g2415 ( 
.A1(n_2269),
.A2(n_2142),
.B1(n_2044),
.B2(n_2086),
.Y(n_2415)
);

AOI22xp5_ASAP7_75t_L g2416 ( 
.A1(n_2269),
.A2(n_2054),
.B1(n_1990),
.B2(n_1973),
.Y(n_2416)
);

INVx3_ASAP7_75t_L g2417 ( 
.A(n_2273),
.Y(n_2417)
);

AOI22xp33_ASAP7_75t_SL g2418 ( 
.A1(n_2154),
.A2(n_1857),
.B1(n_1843),
.B2(n_2105),
.Y(n_2418)
);

BUFx6f_ASAP7_75t_L g2419 ( 
.A(n_2397),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2200),
.Y(n_2420)
);

CKINVDCx20_ASAP7_75t_R g2421 ( 
.A(n_2182),
.Y(n_2421)
);

INVx2_ASAP7_75t_SL g2422 ( 
.A(n_2182),
.Y(n_2422)
);

OAI22xp33_ASAP7_75t_L g2423 ( 
.A1(n_2292),
.A2(n_1954),
.B1(n_1932),
.B2(n_2045),
.Y(n_2423)
);

BUFx4_ASAP7_75t_SL g2424 ( 
.A(n_2320),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2201),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2243),
.Y(n_2426)
);

AOI22xp33_ASAP7_75t_L g2427 ( 
.A1(n_2292),
.A2(n_2056),
.B1(n_2088),
.B2(n_2008),
.Y(n_2427)
);

CKINVDCx5p33_ASAP7_75t_R g2428 ( 
.A(n_2165),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2413),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2218),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2213),
.Y(n_2431)
);

CKINVDCx11_ASAP7_75t_R g2432 ( 
.A(n_2181),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2235),
.Y(n_2433)
);

INVxp67_ASAP7_75t_SL g2434 ( 
.A(n_2326),
.Y(n_2434)
);

CKINVDCx6p67_ASAP7_75t_R g2435 ( 
.A(n_2160),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2216),
.Y(n_2436)
);

INVx1_ASAP7_75t_SL g2437 ( 
.A(n_2165),
.Y(n_2437)
);

CKINVDCx11_ASAP7_75t_R g2438 ( 
.A(n_2256),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2238),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2217),
.Y(n_2440)
);

AOI22xp33_ASAP7_75t_SL g2441 ( 
.A1(n_2224),
.A2(n_1843),
.B1(n_1829),
.B2(n_2018),
.Y(n_2441)
);

BUFx12f_ASAP7_75t_L g2442 ( 
.A(n_2161),
.Y(n_2442)
);

BUFx6f_ASAP7_75t_L g2443 ( 
.A(n_2397),
.Y(n_2443)
);

BUFx10_ASAP7_75t_L g2444 ( 
.A(n_2341),
.Y(n_2444)
);

AOI22xp33_ASAP7_75t_SL g2445 ( 
.A1(n_2224),
.A2(n_2017),
.B1(n_2085),
.B2(n_1878),
.Y(n_2445)
);

OAI22xp5_ASAP7_75t_SL g2446 ( 
.A1(n_2195),
.A2(n_1910),
.B1(n_2085),
.B2(n_1848),
.Y(n_2446)
);

AOI22xp33_ASAP7_75t_L g2447 ( 
.A1(n_2403),
.A2(n_2021),
.B1(n_2082),
.B2(n_2063),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2220),
.Y(n_2448)
);

OAI22xp5_ASAP7_75t_L g2449 ( 
.A1(n_2195),
.A2(n_2078),
.B1(n_2061),
.B2(n_2077),
.Y(n_2449)
);

BUFx6f_ASAP7_75t_L g2450 ( 
.A(n_2397),
.Y(n_2450)
);

BUFx2_ASAP7_75t_L g2451 ( 
.A(n_2212),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2225),
.Y(n_2452)
);

OAI21xp33_ASAP7_75t_L g2453 ( 
.A1(n_2173),
.A2(n_1998),
.B(n_1995),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2246),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2249),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2226),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2275),
.Y(n_2457)
);

BUFx12f_ASAP7_75t_L g2458 ( 
.A(n_2161),
.Y(n_2458)
);

AOI22xp33_ASAP7_75t_L g2459 ( 
.A1(n_2403),
.A2(n_2082),
.B1(n_2123),
.B2(n_1925),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2167),
.B(n_2001),
.Y(n_2460)
);

AOI22xp33_ASAP7_75t_L g2461 ( 
.A1(n_2258),
.A2(n_1916),
.B1(n_1949),
.B2(n_1934),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_SL g2462 ( 
.A(n_2257),
.Y(n_2462)
);

BUFx4f_ASAP7_75t_SL g2463 ( 
.A(n_2379),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2268),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2276),
.Y(n_2465)
);

BUFx3_ASAP7_75t_L g2466 ( 
.A(n_2164),
.Y(n_2466)
);

AOI22xp33_ASAP7_75t_SL g2467 ( 
.A1(n_2224),
.A2(n_1902),
.B1(n_2099),
.B2(n_1921),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2159),
.Y(n_2468)
);

CKINVDCx20_ASAP7_75t_R g2469 ( 
.A(n_2320),
.Y(n_2469)
);

BUFx12f_ASAP7_75t_L g2470 ( 
.A(n_2168),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2227),
.Y(n_2471)
);

INVx1_ASAP7_75t_SL g2472 ( 
.A(n_2169),
.Y(n_2472)
);

AOI22xp33_ASAP7_75t_L g2473 ( 
.A1(n_2258),
.A2(n_2111),
.B1(n_1917),
.B2(n_2080),
.Y(n_2473)
);

AOI22xp33_ASAP7_75t_L g2474 ( 
.A1(n_2208),
.A2(n_2069),
.B1(n_2003),
.B2(n_2075),
.Y(n_2474)
);

AOI22xp33_ASAP7_75t_L g2475 ( 
.A1(n_2208),
.A2(n_2075),
.B1(n_2108),
.B2(n_2104),
.Y(n_2475)
);

OAI21xp5_ASAP7_75t_SL g2476 ( 
.A1(n_2176),
.A2(n_1902),
.B(n_1874),
.Y(n_2476)
);

BUFx3_ASAP7_75t_L g2477 ( 
.A(n_2232),
.Y(n_2477)
);

OAI22xp5_ASAP7_75t_L g2478 ( 
.A1(n_2250),
.A2(n_2059),
.B1(n_1827),
.B2(n_2099),
.Y(n_2478)
);

BUFx6f_ASAP7_75t_L g2479 ( 
.A(n_2402),
.Y(n_2479)
);

BUFx2_ASAP7_75t_L g2480 ( 
.A(n_2212),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2239),
.Y(n_2481)
);

NAND2x1p5_ASAP7_75t_L g2482 ( 
.A(n_2155),
.B(n_1879),
.Y(n_2482)
);

OAI22xp5_ASAP7_75t_L g2483 ( 
.A1(n_2242),
.A2(n_2073),
.B1(n_2094),
.B2(n_2134),
.Y(n_2483)
);

OAI22xp33_ASAP7_75t_L g2484 ( 
.A1(n_2211),
.A2(n_2101),
.B1(n_2106),
.B2(n_2004),
.Y(n_2484)
);

BUFx3_ASAP7_75t_L g2485 ( 
.A(n_2252),
.Y(n_2485)
);

BUFx12f_ASAP7_75t_L g2486 ( 
.A(n_2168),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2281),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2282),
.Y(n_2488)
);

AOI22xp33_ASAP7_75t_SL g2489 ( 
.A1(n_2155),
.A2(n_1846),
.B1(n_1881),
.B2(n_1886),
.Y(n_2489)
);

BUFx3_ASAP7_75t_L g2490 ( 
.A(n_2209),
.Y(n_2490)
);

INVx6_ASAP7_75t_L g2491 ( 
.A(n_2188),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2278),
.Y(n_2492)
);

BUFx8_ASAP7_75t_L g2493 ( 
.A(n_2267),
.Y(n_2493)
);

BUFx6f_ASAP7_75t_L g2494 ( 
.A(n_2402),
.Y(n_2494)
);

AOI22xp33_ASAP7_75t_L g2495 ( 
.A1(n_2170),
.A2(n_2024),
.B1(n_2091),
.B2(n_2066),
.Y(n_2495)
);

AOI21xp33_ASAP7_75t_L g2496 ( 
.A1(n_2364),
.A2(n_1810),
.B(n_1826),
.Y(n_2496)
);

AOI22xp33_ASAP7_75t_L g2497 ( 
.A1(n_2170),
.A2(n_2090),
.B1(n_2071),
.B2(n_2081),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2287),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2280),
.Y(n_2499)
);

INVx6_ASAP7_75t_L g2500 ( 
.A(n_2188),
.Y(n_2500)
);

AOI22xp33_ASAP7_75t_SL g2501 ( 
.A1(n_2155),
.A2(n_1912),
.B1(n_2137),
.B2(n_1836),
.Y(n_2501)
);

AOI22xp33_ASAP7_75t_SL g2502 ( 
.A1(n_2184),
.A2(n_2007),
.B1(n_2120),
.B2(n_2112),
.Y(n_2502)
);

BUFx3_ASAP7_75t_L g2503 ( 
.A(n_2361),
.Y(n_2503)
);

AOI22xp5_ASAP7_75t_L g2504 ( 
.A1(n_2190),
.A2(n_1986),
.B1(n_1958),
.B2(n_1936),
.Y(n_2504)
);

INVx6_ASAP7_75t_L g2505 ( 
.A(n_2172),
.Y(n_2505)
);

AOI22xp33_ASAP7_75t_SL g2506 ( 
.A1(n_2184),
.A2(n_2007),
.B1(n_2016),
.B2(n_2040),
.Y(n_2506)
);

INVx2_ASAP7_75t_SL g2507 ( 
.A(n_2169),
.Y(n_2507)
);

OAI22xp5_ASAP7_75t_L g2508 ( 
.A1(n_2242),
.A2(n_2097),
.B1(n_2071),
.B2(n_1913),
.Y(n_2508)
);

BUFx6f_ASAP7_75t_L g2509 ( 
.A(n_2402),
.Y(n_2509)
);

INVx4_ASAP7_75t_L g2510 ( 
.A(n_2273),
.Y(n_2510)
);

BUFx4f_ASAP7_75t_SL g2511 ( 
.A(n_2272),
.Y(n_2511)
);

AOI22xp33_ASAP7_75t_L g2512 ( 
.A1(n_2211),
.A2(n_2072),
.B1(n_2100),
.B2(n_2040),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2293),
.Y(n_2513)
);

BUFx12f_ASAP7_75t_L g2514 ( 
.A(n_2228),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2305),
.Y(n_2515)
);

NAND2x1p5_ASAP7_75t_L g2516 ( 
.A(n_2184),
.B(n_2016),
.Y(n_2516)
);

HB1xp67_ASAP7_75t_L g2517 ( 
.A(n_2173),
.Y(n_2517)
);

BUFx3_ASAP7_75t_L g2518 ( 
.A(n_2334),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2185),
.B(n_1962),
.Y(n_2519)
);

BUFx2_ASAP7_75t_L g2520 ( 
.A(n_2401),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2289),
.Y(n_2521)
);

AOI22xp33_ASAP7_75t_L g2522 ( 
.A1(n_2211),
.A2(n_2373),
.B1(n_2194),
.B2(n_2191),
.Y(n_2522)
);

AOI22xp33_ASAP7_75t_SL g2523 ( 
.A1(n_2394),
.A2(n_2016),
.B1(n_1953),
.B2(n_1947),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2333),
.Y(n_2524)
);

AOI22xp33_ASAP7_75t_SL g2525 ( 
.A1(n_2234),
.A2(n_1947),
.B1(n_1953),
.B2(n_1859),
.Y(n_2525)
);

BUFx3_ASAP7_75t_L g2526 ( 
.A(n_2171),
.Y(n_2526)
);

AOI22xp5_ASAP7_75t_L g2527 ( 
.A1(n_2248),
.A2(n_2072),
.B1(n_2046),
.B2(n_1975),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2197),
.B(n_1962),
.Y(n_2528)
);

OAI22xp33_ASAP7_75t_L g2529 ( 
.A1(n_2265),
.A2(n_1823),
.B1(n_1811),
.B2(n_1896),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2337),
.Y(n_2530)
);

INVx4_ASAP7_75t_L g2531 ( 
.A(n_2273),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2338),
.Y(n_2532)
);

CKINVDCx5p33_ASAP7_75t_R g2533 ( 
.A(n_2187),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2302),
.Y(n_2534)
);

INVx8_ASAP7_75t_L g2535 ( 
.A(n_2156),
.Y(n_2535)
);

AOI22xp33_ASAP7_75t_L g2536 ( 
.A1(n_2230),
.A2(n_2138),
.B1(n_2147),
.B2(n_1885),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2307),
.Y(n_2537)
);

CKINVDCx5p33_ASAP7_75t_R g2538 ( 
.A(n_2187),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2340),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2308),
.Y(n_2540)
);

CKINVDCx20_ASAP7_75t_R g2541 ( 
.A(n_2229),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2376),
.Y(n_2542)
);

OAI22xp5_ASAP7_75t_L g2543 ( 
.A1(n_2248),
.A2(n_2051),
.B1(n_2031),
.B2(n_2033),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2313),
.Y(n_2544)
);

CKINVDCx20_ASAP7_75t_R g2545 ( 
.A(n_2229),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2387),
.Y(n_2546)
);

AOI22xp33_ASAP7_75t_L g2547 ( 
.A1(n_2186),
.A2(n_2138),
.B1(n_1964),
.B2(n_2060),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2404),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2316),
.Y(n_2549)
);

OAI22xp33_ASAP7_75t_L g2550 ( 
.A1(n_2284),
.A2(n_2074),
.B1(n_2109),
.B2(n_1926),
.Y(n_2550)
);

INVx6_ASAP7_75t_L g2551 ( 
.A(n_2350),
.Y(n_2551)
);

AOI22xp33_ASAP7_75t_L g2552 ( 
.A1(n_2366),
.A2(n_2060),
.B1(n_1966),
.B2(n_1964),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2324),
.Y(n_2553)
);

BUFx6f_ASAP7_75t_L g2554 ( 
.A(n_2288),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2159),
.Y(n_2555)
);

BUFx12f_ASAP7_75t_L g2556 ( 
.A(n_2341),
.Y(n_2556)
);

AOI21xp5_ASAP7_75t_L g2557 ( 
.A1(n_2255),
.A2(n_2326),
.B(n_2263),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2162),
.Y(n_2558)
);

AOI22xp33_ASAP7_75t_SL g2559 ( 
.A1(n_2189),
.A2(n_2145),
.B1(n_1923),
.B2(n_1922),
.Y(n_2559)
);

OAI22xp5_ASAP7_75t_L g2560 ( 
.A1(n_2263),
.A2(n_2049),
.B1(n_2032),
.B2(n_2050),
.Y(n_2560)
);

CKINVDCx6p67_ASAP7_75t_R g2561 ( 
.A(n_2189),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2222),
.B(n_1966),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2162),
.Y(n_2563)
);

CKINVDCx5p33_ASAP7_75t_R g2564 ( 
.A(n_2300),
.Y(n_2564)
);

AOI22xp33_ASAP7_75t_SL g2565 ( 
.A1(n_2360),
.A2(n_2336),
.B1(n_2233),
.B2(n_2385),
.Y(n_2565)
);

BUFx6f_ASAP7_75t_L g2566 ( 
.A(n_2288),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2177),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2339),
.Y(n_2568)
);

AOI22xp33_ASAP7_75t_L g2569 ( 
.A1(n_2366),
.A2(n_2116),
.B1(n_2117),
.B2(n_1914),
.Y(n_2569)
);

AOI22xp33_ASAP7_75t_L g2570 ( 
.A1(n_2193),
.A2(n_2183),
.B1(n_2255),
.B2(n_2344),
.Y(n_2570)
);

BUFx6f_ASAP7_75t_L g2571 ( 
.A(n_2288),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2352),
.Y(n_2572)
);

OAI22xp5_ASAP7_75t_L g2573 ( 
.A1(n_2385),
.A2(n_2038),
.B1(n_1818),
.B2(n_1838),
.Y(n_2573)
);

AOI22xp33_ASAP7_75t_L g2574 ( 
.A1(n_2193),
.A2(n_2364),
.B1(n_2331),
.B2(n_2329),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2241),
.B(n_2116),
.Y(n_2575)
);

BUFx2_ASAP7_75t_L g2576 ( 
.A(n_2401),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2177),
.Y(n_2577)
);

AOI22xp33_ASAP7_75t_SL g2578 ( 
.A1(n_2446),
.A2(n_2260),
.B1(n_2271),
.B2(n_2270),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2429),
.Y(n_2579)
);

CKINVDCx20_ASAP7_75t_R g2580 ( 
.A(n_2421),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2420),
.Y(n_2581)
);

NOR2xp33_ASAP7_75t_L g2582 ( 
.A(n_2449),
.B(n_2392),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2430),
.Y(n_2583)
);

BUFx3_ASAP7_75t_L g2584 ( 
.A(n_2466),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2425),
.Y(n_2585)
);

BUFx6f_ASAP7_75t_L g2586 ( 
.A(n_2520),
.Y(n_2586)
);

AND2x2_ASAP7_75t_L g2587 ( 
.A(n_2562),
.B(n_2241),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2433),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2426),
.Y(n_2589)
);

CKINVDCx20_ASAP7_75t_R g2590 ( 
.A(n_2469),
.Y(n_2590)
);

AOI22xp33_ASAP7_75t_L g2591 ( 
.A1(n_2447),
.A2(n_2247),
.B1(n_2362),
.B2(n_2207),
.Y(n_2591)
);

HB1xp67_ASAP7_75t_L g2592 ( 
.A(n_2517),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2431),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_L g2594 ( 
.A(n_2576),
.B(n_2321),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2439),
.Y(n_2595)
);

OAI22xp5_ASAP7_75t_L g2596 ( 
.A1(n_2561),
.A2(n_2390),
.B1(n_2219),
.B2(n_2303),
.Y(n_2596)
);

BUFx6f_ASAP7_75t_L g2597 ( 
.A(n_2419),
.Y(n_2597)
);

OAI22xp5_ASAP7_75t_L g2598 ( 
.A1(n_2476),
.A2(n_2219),
.B1(n_2390),
.B2(n_2266),
.Y(n_2598)
);

INVx3_ASAP7_75t_L g2599 ( 
.A(n_2510),
.Y(n_2599)
);

OAI22xp5_ASAP7_75t_L g2600 ( 
.A1(n_2459),
.A2(n_2219),
.B1(n_2303),
.B2(n_2266),
.Y(n_2600)
);

AOI222xp33_ASAP7_75t_L g2601 ( 
.A1(n_2437),
.A2(n_2306),
.B1(n_2321),
.B2(n_2405),
.C1(n_2357),
.C2(n_2233),
.Y(n_2601)
);

OAI21xp5_ASAP7_75t_SL g2602 ( 
.A1(n_2445),
.A2(n_2309),
.B(n_2342),
.Y(n_2602)
);

AOI22xp33_ASAP7_75t_L g2603 ( 
.A1(n_2423),
.A2(n_2362),
.B1(n_2365),
.B2(n_2345),
.Y(n_2603)
);

AOI22xp33_ASAP7_75t_L g2604 ( 
.A1(n_2574),
.A2(n_2362),
.B1(n_2345),
.B2(n_2322),
.Y(n_2604)
);

BUFx3_ASAP7_75t_L g2605 ( 
.A(n_2535),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2436),
.Y(n_2606)
);

OAI22xp5_ASAP7_75t_L g2607 ( 
.A1(n_2441),
.A2(n_2411),
.B1(n_2358),
.B2(n_2309),
.Y(n_2607)
);

BUFx3_ASAP7_75t_L g2608 ( 
.A(n_2535),
.Y(n_2608)
);

OAI22xp5_ASAP7_75t_L g2609 ( 
.A1(n_2467),
.A2(n_2323),
.B1(n_2386),
.B2(n_2325),
.Y(n_2609)
);

INVx4_ASAP7_75t_L g2610 ( 
.A(n_2551),
.Y(n_2610)
);

HB1xp67_ASAP7_75t_L g2611 ( 
.A(n_2575),
.Y(n_2611)
);

AOI22xp33_ASAP7_75t_L g2612 ( 
.A1(n_2453),
.A2(n_2322),
.B1(n_2332),
.B2(n_2375),
.Y(n_2612)
);

OAI22xp5_ASAP7_75t_L g2613 ( 
.A1(n_2565),
.A2(n_2323),
.B1(n_2386),
.B2(n_2325),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2440),
.Y(n_2614)
);

CKINVDCx8_ASAP7_75t_R g2615 ( 
.A(n_2428),
.Y(n_2615)
);

OAI22xp33_ASAP7_75t_L g2616 ( 
.A1(n_2472),
.A2(n_2323),
.B1(n_2291),
.B2(n_2153),
.Y(n_2616)
);

BUFx4f_ASAP7_75t_L g2617 ( 
.A(n_2470),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2448),
.Y(n_2618)
);

AOI222xp33_ASAP7_75t_L g2619 ( 
.A1(n_2507),
.A2(n_2306),
.B1(n_2405),
.B2(n_2357),
.C1(n_2214),
.C2(n_2393),
.Y(n_2619)
);

BUFx12f_ASAP7_75t_L g2620 ( 
.A(n_2432),
.Y(n_2620)
);

BUFx4f_ASAP7_75t_SL g2621 ( 
.A(n_2486),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2452),
.Y(n_2622)
);

AOI22xp33_ASAP7_75t_L g2623 ( 
.A1(n_2496),
.A2(n_2332),
.B1(n_2375),
.B2(n_2410),
.Y(n_2623)
);

OAI22xp5_ASAP7_75t_L g2624 ( 
.A1(n_2434),
.A2(n_2291),
.B1(n_2317),
.B2(n_2315),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2456),
.Y(n_2625)
);

OAI21xp33_ASAP7_75t_L g2626 ( 
.A1(n_2416),
.A2(n_2039),
.B(n_2383),
.Y(n_2626)
);

INVxp67_ASAP7_75t_SL g2627 ( 
.A(n_2483),
.Y(n_2627)
);

INVx4_ASAP7_75t_L g2628 ( 
.A(n_2551),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2454),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2471),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2481),
.Y(n_2631)
);

AOI22xp5_ASAP7_75t_L g2632 ( 
.A1(n_2473),
.A2(n_2399),
.B1(n_2240),
.B2(n_2274),
.Y(n_2632)
);

AOI222xp33_ASAP7_75t_L g2633 ( 
.A1(n_2552),
.A2(n_2393),
.B1(n_2240),
.B2(n_2315),
.C1(n_2317),
.C2(n_2296),
.Y(n_2633)
);

AOI22xp33_ASAP7_75t_L g2634 ( 
.A1(n_2570),
.A2(n_2569),
.B1(n_2418),
.B2(n_2508),
.Y(n_2634)
);

OAI21xp33_ASAP7_75t_L g2635 ( 
.A1(n_2461),
.A2(n_2039),
.B(n_2210),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2460),
.B(n_2264),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2519),
.B(n_2264),
.Y(n_2637)
);

INVx3_ASAP7_75t_L g2638 ( 
.A(n_2510),
.Y(n_2638)
);

INVxp67_ASAP7_75t_L g2639 ( 
.A(n_2503),
.Y(n_2639)
);

AOI22xp33_ASAP7_75t_L g2640 ( 
.A1(n_2547),
.A2(n_2301),
.B1(n_2310),
.B2(n_2251),
.Y(n_2640)
);

AOI22xp33_ASAP7_75t_L g2641 ( 
.A1(n_2489),
.A2(n_2406),
.B1(n_2412),
.B2(n_2274),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2487),
.Y(n_2642)
);

AOI22xp33_ASAP7_75t_SL g2643 ( 
.A1(n_2478),
.A2(n_2291),
.B1(n_2342),
.B2(n_2202),
.Y(n_2643)
);

AND2x4_ASAP7_75t_L g2644 ( 
.A(n_2419),
.B(n_2377),
.Y(n_2644)
);

OAI22xp5_ASAP7_75t_L g2645 ( 
.A1(n_2559),
.A2(n_2291),
.B1(n_2223),
.B2(n_2236),
.Y(n_2645)
);

OAI21xp5_ASAP7_75t_SL g2646 ( 
.A1(n_2501),
.A2(n_2304),
.B(n_2312),
.Y(n_2646)
);

OAI22xp5_ASAP7_75t_L g2647 ( 
.A1(n_2427),
.A2(n_2192),
.B1(n_2236),
.B2(n_2223),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2488),
.Y(n_2648)
);

OAI21xp5_ASAP7_75t_SL g2649 ( 
.A1(n_2523),
.A2(n_2502),
.B(n_2506),
.Y(n_2649)
);

AOI22xp33_ASAP7_75t_L g2650 ( 
.A1(n_2525),
.A2(n_2296),
.B1(n_2328),
.B2(n_2335),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_2541),
.B(n_2297),
.Y(n_2651)
);

AND2x2_ASAP7_75t_L g2652 ( 
.A(n_2528),
.B(n_2327),
.Y(n_2652)
);

BUFx6f_ASAP7_75t_L g2653 ( 
.A(n_2419),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2457),
.B(n_2327),
.Y(n_2654)
);

AOI22xp33_ASAP7_75t_L g2655 ( 
.A1(n_2550),
.A2(n_2363),
.B1(n_2196),
.B2(n_2388),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2498),
.Y(n_2656)
);

HB1xp67_ASAP7_75t_L g2657 ( 
.A(n_2492),
.Y(n_2657)
);

OAI22xp5_ASAP7_75t_L g2658 ( 
.A1(n_2475),
.A2(n_2192),
.B1(n_2202),
.B2(n_2351),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2513),
.B(n_2285),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2455),
.Y(n_2660)
);

BUFx4f_ASAP7_75t_SL g2661 ( 
.A(n_2556),
.Y(n_2661)
);

BUFx4f_ASAP7_75t_SL g2662 ( 
.A(n_2514),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2499),
.B(n_2521),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2515),
.B(n_2285),
.Y(n_2664)
);

INVx3_ASAP7_75t_L g2665 ( 
.A(n_2531),
.Y(n_2665)
);

OAI22xp5_ASAP7_75t_L g2666 ( 
.A1(n_2415),
.A2(n_2351),
.B1(n_2196),
.B2(n_2389),
.Y(n_2666)
);

AOI22xp33_ASAP7_75t_SL g2667 ( 
.A1(n_2573),
.A2(n_2347),
.B1(n_2319),
.B2(n_2389),
.Y(n_2667)
);

AOI22xp33_ASAP7_75t_SL g2668 ( 
.A1(n_2491),
.A2(n_2500),
.B1(n_2538),
.B2(n_2533),
.Y(n_2668)
);

AOI22xp33_ASAP7_75t_L g2669 ( 
.A1(n_2536),
.A2(n_2015),
.B1(n_2391),
.B2(n_2237),
.Y(n_2669)
);

AOI22xp33_ASAP7_75t_L g2670 ( 
.A1(n_2474),
.A2(n_2237),
.B1(n_2380),
.B2(n_2117),
.Y(n_2670)
);

AOI22xp33_ASAP7_75t_L g2671 ( 
.A1(n_2484),
.A2(n_2380),
.B1(n_2395),
.B2(n_2148),
.Y(n_2671)
);

NAND2xp33_ASAP7_75t_SL g2672 ( 
.A(n_2531),
.B(n_2297),
.Y(n_2672)
);

BUFx2_ASAP7_75t_L g2673 ( 
.A(n_2443),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2524),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2530),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2532),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2539),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2542),
.B(n_2215),
.Y(n_2678)
);

HB1xp67_ASAP7_75t_L g2679 ( 
.A(n_2443),
.Y(n_2679)
);

OAI22xp5_ASAP7_75t_L g2680 ( 
.A1(n_2512),
.A2(n_2389),
.B1(n_2205),
.B2(n_2206),
.Y(n_2680)
);

NAND2x1p5_ASAP7_75t_L g2681 ( 
.A(n_2526),
.B(n_2396),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2546),
.Y(n_2682)
);

AOI22xp33_ASAP7_75t_L g2683 ( 
.A1(n_2495),
.A2(n_1842),
.B1(n_1849),
.B2(n_2206),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2534),
.Y(n_2684)
);

AND2x2_ASAP7_75t_SL g2685 ( 
.A(n_2451),
.B(n_2221),
.Y(n_2685)
);

OAI22xp5_ASAP7_75t_SL g2686 ( 
.A1(n_2491),
.A2(n_2180),
.B1(n_2158),
.B2(n_2311),
.Y(n_2686)
);

OAI22xp5_ASAP7_75t_L g2687 ( 
.A1(n_2497),
.A2(n_2205),
.B1(n_2304),
.B2(n_2179),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2548),
.B(n_2110),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2464),
.B(n_2110),
.Y(n_2689)
);

OAI22xp33_ASAP7_75t_L g2690 ( 
.A1(n_2500),
.A2(n_2221),
.B1(n_2283),
.B2(n_2299),
.Y(n_2690)
);

AOI22xp33_ASAP7_75t_L g2691 ( 
.A1(n_2522),
.A2(n_2253),
.B1(n_2145),
.B2(n_2179),
.Y(n_2691)
);

INVxp67_ASAP7_75t_L g2692 ( 
.A(n_2657),
.Y(n_2692)
);

OAI22xp5_ASAP7_75t_L g2693 ( 
.A1(n_2607),
.A2(n_2527),
.B1(n_2529),
.B2(n_2516),
.Y(n_2693)
);

AOI22xp33_ASAP7_75t_SL g2694 ( 
.A1(n_2598),
.A2(n_2480),
.B1(n_2417),
.B2(n_2463),
.Y(n_2694)
);

AOI22xp33_ASAP7_75t_L g2695 ( 
.A1(n_2598),
.A2(n_2504),
.B1(n_2464),
.B2(n_2465),
.Y(n_2695)
);

AOI22xp33_ASAP7_75t_L g2696 ( 
.A1(n_2591),
.A2(n_2465),
.B1(n_2468),
.B2(n_2555),
.Y(n_2696)
);

NAND3xp33_ASAP7_75t_L g2697 ( 
.A(n_2619),
.B(n_2557),
.C(n_2493),
.Y(n_2697)
);

OAI22xp5_ASAP7_75t_L g2698 ( 
.A1(n_2634),
.A2(n_2482),
.B1(n_2545),
.B2(n_2417),
.Y(n_2698)
);

OAI22xp5_ASAP7_75t_L g2699 ( 
.A1(n_2603),
.A2(n_2468),
.B1(n_2555),
.B2(n_2558),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2579),
.Y(n_2700)
);

AOI22xp33_ASAP7_75t_L g2701 ( 
.A1(n_2604),
.A2(n_2558),
.B1(n_2563),
.B2(n_2577),
.Y(n_2701)
);

NAND3xp33_ASAP7_75t_L g2702 ( 
.A(n_2619),
.B(n_2493),
.C(n_2543),
.Y(n_2702)
);

OAI22xp5_ASAP7_75t_L g2703 ( 
.A1(n_2655),
.A2(n_2563),
.B1(n_2567),
.B2(n_2577),
.Y(n_2703)
);

AOI22xp33_ASAP7_75t_L g2704 ( 
.A1(n_2612),
.A2(n_2567),
.B1(n_2136),
.B2(n_2442),
.Y(n_2704)
);

AOI22xp33_ASAP7_75t_L g2705 ( 
.A1(n_2600),
.A2(n_2136),
.B1(n_2458),
.B2(n_2145),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2611),
.B(n_2537),
.Y(n_2706)
);

OAI22xp5_ASAP7_75t_L g2707 ( 
.A1(n_2641),
.A2(n_2422),
.B1(n_2414),
.B2(n_2407),
.Y(n_2707)
);

AOI22xp33_ASAP7_75t_L g2708 ( 
.A1(n_2627),
.A2(n_2145),
.B1(n_2560),
.B2(n_2346),
.Y(n_2708)
);

AOI22xp33_ASAP7_75t_L g2709 ( 
.A1(n_2635),
.A2(n_2346),
.B1(n_2349),
.B2(n_2518),
.Y(n_2709)
);

NOR3xp33_ASAP7_75t_L g2710 ( 
.A(n_2610),
.B(n_2156),
.C(n_2204),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2652),
.B(n_2572),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2587),
.B(n_2540),
.Y(n_2712)
);

AOI22xp33_ASAP7_75t_L g2713 ( 
.A1(n_2623),
.A2(n_2349),
.B1(n_2314),
.B2(n_2254),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2581),
.Y(n_2714)
);

AOI22xp33_ASAP7_75t_L g2715 ( 
.A1(n_2633),
.A2(n_2254),
.B1(n_2314),
.B2(n_2299),
.Y(n_2715)
);

AOI22xp33_ASAP7_75t_L g2716 ( 
.A1(n_2633),
.A2(n_2283),
.B1(n_2407),
.B2(n_2414),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2663),
.B(n_2544),
.Y(n_2717)
);

AOI22xp33_ASAP7_75t_SL g2718 ( 
.A1(n_2596),
.A2(n_2511),
.B1(n_2505),
.B2(n_2369),
.Y(n_2718)
);

AOI22xp33_ASAP7_75t_L g2719 ( 
.A1(n_2582),
.A2(n_2672),
.B1(n_2683),
.B2(n_2626),
.Y(n_2719)
);

AOI22xp33_ASAP7_75t_L g2720 ( 
.A1(n_2609),
.A2(n_2359),
.B1(n_2381),
.B2(n_2400),
.Y(n_2720)
);

AOI22xp5_ASAP7_75t_L g2721 ( 
.A1(n_2649),
.A2(n_2505),
.B1(n_2462),
.B2(n_2477),
.Y(n_2721)
);

INVx4_ASAP7_75t_R g2722 ( 
.A(n_2605),
.Y(n_2722)
);

OA21x2_ASAP7_75t_L g2723 ( 
.A1(n_2602),
.A2(n_2149),
.B(n_1978),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2593),
.B(n_2606),
.Y(n_2724)
);

AOI22xp33_ASAP7_75t_L g2725 ( 
.A1(n_2613),
.A2(n_2650),
.B1(n_2640),
.B2(n_2645),
.Y(n_2725)
);

AOI22xp33_ASAP7_75t_L g2726 ( 
.A1(n_2601),
.A2(n_2553),
.B1(n_2568),
.B2(n_2549),
.Y(n_2726)
);

AOI22xp33_ASAP7_75t_L g2727 ( 
.A1(n_2601),
.A2(n_2119),
.B1(n_2485),
.B2(n_2131),
.Y(n_2727)
);

NOR2xp33_ASAP7_75t_L g2728 ( 
.A(n_2639),
.B(n_2590),
.Y(n_2728)
);

AOI22xp33_ASAP7_75t_L g2729 ( 
.A1(n_2645),
.A2(n_2359),
.B1(n_2381),
.B2(n_2400),
.Y(n_2729)
);

AOI22xp33_ASAP7_75t_L g2730 ( 
.A1(n_2592),
.A2(n_2119),
.B1(n_2131),
.B2(n_2435),
.Y(n_2730)
);

AOI22xp33_ASAP7_75t_L g2731 ( 
.A1(n_2647),
.A2(n_2408),
.B1(n_2409),
.B2(n_2198),
.Y(n_2731)
);

AOI22xp33_ASAP7_75t_L g2732 ( 
.A1(n_2624),
.A2(n_2408),
.B1(n_2409),
.B2(n_2198),
.Y(n_2732)
);

AOI22xp33_ASAP7_75t_SL g2733 ( 
.A1(n_2624),
.A2(n_2369),
.B1(n_2348),
.B2(n_2199),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2614),
.B(n_2443),
.Y(n_2734)
);

AOI22xp33_ASAP7_75t_L g2735 ( 
.A1(n_2678),
.A2(n_2157),
.B1(n_2199),
.B2(n_2152),
.Y(n_2735)
);

AOI222xp33_ASAP7_75t_L g2736 ( 
.A1(n_2617),
.A2(n_2462),
.B1(n_2438),
.B2(n_2490),
.C1(n_2330),
.C2(n_2444),
.Y(n_2736)
);

OAI22xp5_ASAP7_75t_L g2737 ( 
.A1(n_2649),
.A2(n_2578),
.B1(n_2643),
.B2(n_2671),
.Y(n_2737)
);

OAI22xp5_ASAP7_75t_L g2738 ( 
.A1(n_2646),
.A2(n_2157),
.B1(n_2396),
.B2(n_2371),
.Y(n_2738)
);

OAI22xp5_ASAP7_75t_L g2739 ( 
.A1(n_2646),
.A2(n_2396),
.B1(n_2371),
.B2(n_2294),
.Y(n_2739)
);

AOI22xp33_ASAP7_75t_L g2740 ( 
.A1(n_2654),
.A2(n_2152),
.B1(n_1853),
.B2(n_1864),
.Y(n_2740)
);

AOI22xp33_ASAP7_75t_L g2741 ( 
.A1(n_2669),
.A2(n_2369),
.B1(n_2348),
.B2(n_2125),
.Y(n_2741)
);

AOI22xp33_ASAP7_75t_SL g2742 ( 
.A1(n_2685),
.A2(n_2369),
.B1(n_2348),
.B2(n_2571),
.Y(n_2742)
);

OA21x2_ASAP7_75t_L g2743 ( 
.A1(n_2602),
.A2(n_1978),
.B(n_2139),
.Y(n_2743)
);

OAI22xp5_ASAP7_75t_L g2744 ( 
.A1(n_2632),
.A2(n_2279),
.B1(n_2294),
.B2(n_2277),
.Y(n_2744)
);

AND2x2_ASAP7_75t_L g2745 ( 
.A(n_2585),
.B(n_2450),
.Y(n_2745)
);

OAI22xp5_ASAP7_75t_L g2746 ( 
.A1(n_2667),
.A2(n_2279),
.B1(n_2277),
.B2(n_2244),
.Y(n_2746)
);

AOI22xp33_ASAP7_75t_L g2747 ( 
.A1(n_2586),
.A2(n_2369),
.B1(n_2348),
.B2(n_1814),
.Y(n_2747)
);

OA21x2_ASAP7_75t_L g2748 ( 
.A1(n_2659),
.A2(n_2141),
.B(n_2150),
.Y(n_2748)
);

INVx2_ASAP7_75t_SL g2749 ( 
.A(n_2584),
.Y(n_2749)
);

AOI221xp5_ASAP7_75t_L g2750 ( 
.A1(n_2636),
.A2(n_2178),
.B1(n_2370),
.B2(n_2564),
.C(n_2122),
.Y(n_2750)
);

AOI22xp33_ASAP7_75t_L g2751 ( 
.A1(n_2586),
.A2(n_2348),
.B1(n_2151),
.B2(n_2124),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2618),
.B(n_2450),
.Y(n_2752)
);

AOI22xp33_ASAP7_75t_L g2753 ( 
.A1(n_2586),
.A2(n_2124),
.B1(n_2566),
.B2(n_2494),
.Y(n_2753)
);

AOI22xp33_ASAP7_75t_L g2754 ( 
.A1(n_2637),
.A2(n_2368),
.B1(n_2367),
.B2(n_2353),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2589),
.Y(n_2755)
);

INVxp67_ASAP7_75t_SL g2756 ( 
.A(n_2679),
.Y(n_2756)
);

OAI222xp33_ASAP7_75t_L g2757 ( 
.A1(n_2690),
.A2(n_2424),
.B1(n_2163),
.B2(n_2231),
.C1(n_2244),
.C2(n_2174),
.Y(n_2757)
);

OAI221xp5_ASAP7_75t_SL g2758 ( 
.A1(n_2670),
.A2(n_2374),
.B1(n_2382),
.B2(n_2384),
.C(n_2398),
.Y(n_2758)
);

OAI22xp5_ASAP7_75t_L g2759 ( 
.A1(n_2681),
.A2(n_2231),
.B1(n_2318),
.B2(n_2174),
.Y(n_2759)
);

OAI221xp5_ASAP7_75t_SL g2760 ( 
.A1(n_2695),
.A2(n_2691),
.B1(n_2664),
.B2(n_2616),
.C(n_2668),
.Y(n_2760)
);

OAI21xp33_ASAP7_75t_L g2761 ( 
.A1(n_2695),
.A2(n_2681),
.B(n_2631),
.Y(n_2761)
);

OA21x2_ASAP7_75t_L g2762 ( 
.A1(n_2708),
.A2(n_2696),
.B(n_2705),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2692),
.B(n_2642),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2711),
.B(n_2706),
.Y(n_2764)
);

AND2x2_ASAP7_75t_L g2765 ( 
.A(n_2700),
.B(n_2648),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2712),
.B(n_2755),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2714),
.B(n_2656),
.Y(n_2767)
);

OA21x2_ASAP7_75t_L g2768 ( 
.A1(n_2696),
.A2(n_2689),
.B(n_2674),
.Y(n_2768)
);

NAND3xp33_ASAP7_75t_L g2769 ( 
.A(n_2697),
.B(n_2628),
.C(n_2610),
.Y(n_2769)
);

OAI221xp5_ASAP7_75t_L g2770 ( 
.A1(n_2727),
.A2(n_2617),
.B1(n_2594),
.B2(n_2651),
.C(n_2628),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2717),
.B(n_2675),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2723),
.B(n_2676),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2724),
.B(n_2677),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2745),
.B(n_2682),
.Y(n_2774)
);

AND2x2_ASAP7_75t_L g2775 ( 
.A(n_2723),
.B(n_2622),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2723),
.B(n_2625),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2756),
.B(n_2630),
.Y(n_2777)
);

AOI22xp33_ASAP7_75t_SL g2778 ( 
.A1(n_2737),
.A2(n_2702),
.B1(n_2698),
.B2(n_2693),
.Y(n_2778)
);

AOI21xp33_ASAP7_75t_L g2779 ( 
.A1(n_2719),
.A2(n_2687),
.B(n_2680),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2699),
.B(n_2583),
.Y(n_2780)
);

AND2x2_ASAP7_75t_L g2781 ( 
.A(n_2748),
.B(n_2588),
.Y(n_2781)
);

OAI21xp5_ASAP7_75t_L g2782 ( 
.A1(n_2694),
.A2(n_2638),
.B(n_2599),
.Y(n_2782)
);

AND2x2_ASAP7_75t_L g2783 ( 
.A(n_2748),
.B(n_2595),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2701),
.B(n_2629),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2748),
.B(n_2660),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2734),
.B(n_2684),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_SL g2787 ( 
.A(n_2718),
.B(n_2599),
.Y(n_2787)
);

OAI21xp5_ASAP7_75t_L g2788 ( 
.A1(n_2721),
.A2(n_2638),
.B(n_2665),
.Y(n_2788)
);

OAI22xp5_ASAP7_75t_L g2789 ( 
.A1(n_2727),
.A2(n_2665),
.B1(n_2658),
.B2(n_2580),
.Y(n_2789)
);

OAI221xp5_ASAP7_75t_SL g2790 ( 
.A1(n_2726),
.A2(n_2608),
.B1(n_2688),
.B2(n_2673),
.C(n_2372),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_SL g2791 ( 
.A(n_2742),
.B(n_2661),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2752),
.B(n_2666),
.Y(n_2792)
);

AND2x2_ASAP7_75t_L g2793 ( 
.A(n_2743),
.B(n_2597),
.Y(n_2793)
);

AOI221xp5_ASAP7_75t_L g2794 ( 
.A1(n_2726),
.A2(n_2686),
.B1(n_2644),
.B2(n_2554),
.C(n_2566),
.Y(n_2794)
);

AND2x2_ASAP7_75t_SL g2795 ( 
.A(n_2743),
.B(n_2644),
.Y(n_2795)
);

AND2x2_ASAP7_75t_L g2796 ( 
.A(n_2743),
.B(n_2597),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2703),
.B(n_2597),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2754),
.B(n_2653),
.Y(n_2798)
);

AOI22xp33_ASAP7_75t_L g2799 ( 
.A1(n_2778),
.A2(n_2725),
.B1(n_2750),
.B2(n_2704),
.Y(n_2799)
);

NOR3xp33_ASAP7_75t_L g2800 ( 
.A(n_2760),
.B(n_2769),
.C(n_2770),
.Y(n_2800)
);

NAND3xp33_ASAP7_75t_L g2801 ( 
.A(n_2779),
.B(n_2730),
.C(n_2709),
.Y(n_2801)
);

NAND3xp33_ASAP7_75t_L g2802 ( 
.A(n_2761),
.B(n_2730),
.C(n_2715),
.Y(n_2802)
);

AND2x2_ASAP7_75t_L g2803 ( 
.A(n_2772),
.B(n_2733),
.Y(n_2803)
);

OR2x2_ASAP7_75t_L g2804 ( 
.A(n_2764),
.B(n_2766),
.Y(n_2804)
);

INVx2_ASAP7_75t_SL g2805 ( 
.A(n_2781),
.Y(n_2805)
);

AND2x4_ASAP7_75t_L g2806 ( 
.A(n_2772),
.B(n_2749),
.Y(n_2806)
);

NAND4xp75_ASAP7_75t_L g2807 ( 
.A(n_2791),
.B(n_2728),
.C(n_2722),
.D(n_2736),
.Y(n_2807)
);

BUFx3_ASAP7_75t_L g2808 ( 
.A(n_2769),
.Y(n_2808)
);

OR2x2_ASAP7_75t_L g2809 ( 
.A(n_2777),
.B(n_2754),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2767),
.B(n_2740),
.Y(n_2810)
);

OR2x2_ASAP7_75t_L g2811 ( 
.A(n_2763),
.B(n_2774),
.Y(n_2811)
);

AND2x2_ASAP7_75t_L g2812 ( 
.A(n_2775),
.B(n_2735),
.Y(n_2812)
);

NOR3xp33_ASAP7_75t_L g2813 ( 
.A(n_2761),
.B(n_2789),
.C(n_2794),
.Y(n_2813)
);

OAI21xp5_ASAP7_75t_L g2814 ( 
.A1(n_2787),
.A2(n_2738),
.B(n_2739),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2781),
.Y(n_2815)
);

NAND4xp75_ASAP7_75t_L g2816 ( 
.A(n_2782),
.B(n_2620),
.C(n_2621),
.D(n_2662),
.Y(n_2816)
);

AND2x2_ASAP7_75t_L g2817 ( 
.A(n_2775),
.B(n_2732),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2783),
.Y(n_2818)
);

NAND3xp33_ASAP7_75t_L g2819 ( 
.A(n_2776),
.B(n_2731),
.C(n_2758),
.Y(n_2819)
);

AND2x4_ASAP7_75t_L g2820 ( 
.A(n_2776),
.B(n_2653),
.Y(n_2820)
);

NAND3xp33_ASAP7_75t_L g2821 ( 
.A(n_2797),
.B(n_2716),
.C(n_2710),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_2783),
.B(n_2741),
.Y(n_2822)
);

AO21x2_ASAP7_75t_L g2823 ( 
.A1(n_2788),
.A2(n_2757),
.B(n_2744),
.Y(n_2823)
);

AOI22xp33_ASAP7_75t_SL g2824 ( 
.A1(n_2762),
.A2(n_2707),
.B1(n_2746),
.B2(n_2759),
.Y(n_2824)
);

OR2x2_ASAP7_75t_L g2825 ( 
.A(n_2771),
.B(n_2753),
.Y(n_2825)
);

AO21x2_ASAP7_75t_L g2826 ( 
.A1(n_2798),
.A2(n_2143),
.B(n_1909),
.Y(n_2826)
);

AND2x2_ASAP7_75t_L g2827 ( 
.A(n_2785),
.B(n_2765),
.Y(n_2827)
);

NOR2xp33_ASAP7_75t_L g2828 ( 
.A(n_2773),
.B(n_2713),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2765),
.Y(n_2829)
);

AOI221xp5_ASAP7_75t_L g2830 ( 
.A1(n_2784),
.A2(n_2729),
.B1(n_2720),
.B2(n_2751),
.C(n_2747),
.Y(n_2830)
);

INVx5_ASAP7_75t_L g2831 ( 
.A(n_2808),
.Y(n_2831)
);

OR2x2_ASAP7_75t_L g2832 ( 
.A(n_2804),
.B(n_2786),
.Y(n_2832)
);

NOR4xp25_ASAP7_75t_L g2833 ( 
.A(n_2799),
.B(n_2790),
.C(n_2780),
.D(n_2767),
.Y(n_2833)
);

INVx5_ASAP7_75t_L g2834 ( 
.A(n_2808),
.Y(n_2834)
);

NOR4xp25_ASAP7_75t_L g2835 ( 
.A(n_2799),
.B(n_2792),
.C(n_2796),
.D(n_2793),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2815),
.Y(n_2836)
);

XOR2x2_ASAP7_75t_L g2837 ( 
.A(n_2816),
.B(n_2762),
.Y(n_2837)
);

AOI22xp5_ASAP7_75t_L g2838 ( 
.A1(n_2800),
.A2(n_2762),
.B1(n_2768),
.B2(n_2795),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2827),
.B(n_2805),
.Y(n_2839)
);

NAND4xp75_ASAP7_75t_L g2840 ( 
.A(n_2814),
.B(n_2762),
.C(n_2795),
.D(n_2768),
.Y(n_2840)
);

OAI31xp33_ASAP7_75t_L g2841 ( 
.A1(n_2813),
.A2(n_2801),
.A3(n_2821),
.B(n_2802),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2812),
.B(n_2817),
.Y(n_2842)
);

NAND4xp75_ASAP7_75t_L g2843 ( 
.A(n_2807),
.B(n_2795),
.C(n_2768),
.D(n_2796),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2815),
.Y(n_2844)
);

HB1xp67_ASAP7_75t_L g2845 ( 
.A(n_2805),
.Y(n_2845)
);

HB1xp67_ASAP7_75t_L g2846 ( 
.A(n_2818),
.Y(n_2846)
);

BUFx2_ASAP7_75t_L g2847 ( 
.A(n_2806),
.Y(n_2847)
);

NAND4xp75_ASAP7_75t_L g2848 ( 
.A(n_2803),
.B(n_2768),
.C(n_2793),
.D(n_2785),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2827),
.B(n_2653),
.Y(n_2849)
);

XNOR2xp5_ASAP7_75t_L g2850 ( 
.A(n_2824),
.B(n_2615),
.Y(n_2850)
);

XOR2x2_ASAP7_75t_L g2851 ( 
.A(n_2828),
.B(n_2444),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2829),
.Y(n_2852)
);

NAND4xp75_ASAP7_75t_SL g2853 ( 
.A(n_2803),
.B(n_2377),
.C(n_2163),
.D(n_2350),
.Y(n_2853)
);

BUFx3_ASAP7_75t_L g2854 ( 
.A(n_2806),
.Y(n_2854)
);

BUFx2_ASAP7_75t_L g2855 ( 
.A(n_2806),
.Y(n_2855)
);

XNOR2x2_ASAP7_75t_L g2856 ( 
.A(n_2819),
.B(n_2377),
.Y(n_2856)
);

OR2x2_ASAP7_75t_L g2857 ( 
.A(n_2818),
.B(n_2811),
.Y(n_2857)
);

AND2x2_ASAP7_75t_L g2858 ( 
.A(n_2817),
.B(n_2450),
.Y(n_2858)
);

HB1xp67_ASAP7_75t_L g2859 ( 
.A(n_2831),
.Y(n_2859)
);

OAI22xp5_ASAP7_75t_L g2860 ( 
.A1(n_2840),
.A2(n_2828),
.B1(n_2809),
.B2(n_2825),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2857),
.Y(n_2861)
);

NOR2xp33_ASAP7_75t_L g2862 ( 
.A(n_2850),
.B(n_2810),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2839),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2857),
.Y(n_2864)
);

INVx2_ASAP7_75t_SL g2865 ( 
.A(n_2847),
.Y(n_2865)
);

XOR2x2_ASAP7_75t_L g2866 ( 
.A(n_2851),
.B(n_2823),
.Y(n_2866)
);

XOR2x2_ASAP7_75t_L g2867 ( 
.A(n_2851),
.B(n_2823),
.Y(n_2867)
);

OAI22xp5_ASAP7_75t_SL g2868 ( 
.A1(n_2835),
.A2(n_2833),
.B1(n_2831),
.B2(n_2834),
.Y(n_2868)
);

XNOR2xp5_ASAP7_75t_L g2869 ( 
.A(n_2837),
.B(n_2812),
.Y(n_2869)
);

AO22x2_ASAP7_75t_L g2870 ( 
.A1(n_2848),
.A2(n_2822),
.B1(n_2820),
.B2(n_2830),
.Y(n_2870)
);

XNOR2x1_ASAP7_75t_L g2871 ( 
.A(n_2837),
.B(n_2822),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2832),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2832),
.Y(n_2873)
);

AND2x2_ASAP7_75t_L g2874 ( 
.A(n_2855),
.B(n_2820),
.Y(n_2874)
);

AOI22x1_ASAP7_75t_L g2875 ( 
.A1(n_2870),
.A2(n_2856),
.B1(n_2845),
.B2(n_2841),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2872),
.Y(n_2876)
);

XNOR2xp5_ASAP7_75t_L g2877 ( 
.A(n_2866),
.B(n_2867),
.Y(n_2877)
);

BUFx3_ASAP7_75t_L g2878 ( 
.A(n_2865),
.Y(n_2878)
);

INVx1_ASAP7_75t_SL g2879 ( 
.A(n_2859),
.Y(n_2879)
);

XNOR2x1_ASAP7_75t_L g2880 ( 
.A(n_2871),
.B(n_2856),
.Y(n_2880)
);

HB1xp67_ASAP7_75t_L g2881 ( 
.A(n_2873),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2861),
.Y(n_2882)
);

XOR2x2_ASAP7_75t_L g2883 ( 
.A(n_2862),
.B(n_2843),
.Y(n_2883)
);

INVx4_ASAP7_75t_L g2884 ( 
.A(n_2859),
.Y(n_2884)
);

XNOR2x2_ASAP7_75t_L g2885 ( 
.A(n_2870),
.B(n_2838),
.Y(n_2885)
);

AOI22x1_ASAP7_75t_L g2886 ( 
.A1(n_2870),
.A2(n_2839),
.B1(n_2846),
.B2(n_2831),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2864),
.Y(n_2887)
);

AOI22xp5_ASAP7_75t_SL g2888 ( 
.A1(n_2860),
.A2(n_2854),
.B1(n_2842),
.B2(n_2849),
.Y(n_2888)
);

NOR2x1_ASAP7_75t_L g2889 ( 
.A(n_2860),
.B(n_2854),
.Y(n_2889)
);

OA22x2_ASAP7_75t_L g2890 ( 
.A1(n_2868),
.A2(n_2849),
.B1(n_2852),
.B2(n_2858),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2863),
.Y(n_2891)
);

AO22x2_ASAP7_75t_L g2892 ( 
.A1(n_2868),
.A2(n_2853),
.B1(n_2834),
.B2(n_2831),
.Y(n_2892)
);

AOI22x1_ASAP7_75t_L g2893 ( 
.A1(n_2869),
.A2(n_2834),
.B1(n_2831),
.B2(n_2836),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2881),
.Y(n_2894)
);

NOR2x1_ASAP7_75t_L g2895 ( 
.A(n_2884),
.B(n_2874),
.Y(n_2895)
);

CKINVDCx20_ASAP7_75t_R g2896 ( 
.A(n_2878),
.Y(n_2896)
);

OAI322xp33_ASAP7_75t_L g2897 ( 
.A1(n_2885),
.A2(n_2844),
.A3(n_2836),
.B1(n_2858),
.B2(n_2834),
.C1(n_2262),
.C2(n_2318),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2884),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2876),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2876),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2887),
.Y(n_2901)
);

INVx1_ASAP7_75t_SL g2902 ( 
.A(n_2879),
.Y(n_2902)
);

INVx2_ASAP7_75t_SL g2903 ( 
.A(n_2889),
.Y(n_2903)
);

BUFx2_ASAP7_75t_L g2904 ( 
.A(n_2892),
.Y(n_2904)
);

OAI322xp33_ASAP7_75t_L g2905 ( 
.A1(n_2877),
.A2(n_2844),
.A3(n_2834),
.B1(n_2262),
.B2(n_1895),
.C1(n_1906),
.C2(n_1876),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2891),
.Y(n_2906)
);

OAI322xp33_ASAP7_75t_L g2907 ( 
.A1(n_2875),
.A2(n_1844),
.A3(n_1860),
.B1(n_2509),
.B2(n_2571),
.C1(n_2566),
.C2(n_2554),
.Y(n_2907)
);

XOR2xp5_ASAP7_75t_L g2908 ( 
.A(n_2883),
.B(n_2820),
.Y(n_2908)
);

OA22x2_ASAP7_75t_L g2909 ( 
.A1(n_2903),
.A2(n_2880),
.B1(n_2886),
.B2(n_2890),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2898),
.Y(n_2910)
);

NOR4xp25_ASAP7_75t_L g2911 ( 
.A(n_2902),
.B(n_2882),
.C(n_2891),
.D(n_2888),
.Y(n_2911)
);

AND4x1_ASAP7_75t_L g2912 ( 
.A(n_2895),
.B(n_2882),
.C(n_2893),
.D(n_2892),
.Y(n_2912)
);

AOI22xp33_ASAP7_75t_SL g2913 ( 
.A1(n_2904),
.A2(n_2826),
.B1(n_2571),
.B2(n_2479),
.Y(n_2913)
);

NOR4xp25_ASAP7_75t_L g2914 ( 
.A(n_2902),
.B(n_1991),
.C(n_2355),
.D(n_1952),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2894),
.Y(n_2915)
);

NAND4xp75_ASAP7_75t_L g2916 ( 
.A(n_2899),
.B(n_2132),
.C(n_2128),
.D(n_2121),
.Y(n_2916)
);

AOI31xp33_ASAP7_75t_L g2917 ( 
.A1(n_2908),
.A2(n_2118),
.A3(n_2129),
.B(n_2121),
.Y(n_2917)
);

NOR4xp25_ASAP7_75t_L g2918 ( 
.A(n_2897),
.B(n_1991),
.C(n_1951),
.D(n_1948),
.Y(n_2918)
);

OAI322xp33_ASAP7_75t_L g2919 ( 
.A1(n_2896),
.A2(n_2479),
.A3(n_2554),
.B1(n_2509),
.B2(n_2494),
.C1(n_2826),
.C2(n_2355),
.Y(n_2919)
);

OAI22xp5_ASAP7_75t_L g2920 ( 
.A1(n_2896),
.A2(n_2901),
.B1(n_2900),
.B2(n_2906),
.Y(n_2920)
);

A2O1A1Ixp33_ASAP7_75t_L g2921 ( 
.A1(n_2907),
.A2(n_2356),
.B(n_2343),
.C(n_2354),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2910),
.Y(n_2922)
);

AOI22xp5_ASAP7_75t_L g2923 ( 
.A1(n_2909),
.A2(n_2905),
.B1(n_2509),
.B2(n_2494),
.Y(n_2923)
);

HB1xp67_ASAP7_75t_L g2924 ( 
.A(n_2915),
.Y(n_2924)
);

OA22x2_ASAP7_75t_L g2925 ( 
.A1(n_2920),
.A2(n_1948),
.B1(n_1951),
.B2(n_2144),
.Y(n_2925)
);

OAI22xp5_ASAP7_75t_L g2926 ( 
.A1(n_2917),
.A2(n_2479),
.B1(n_2378),
.B2(n_2298),
.Y(n_2926)
);

AOI22xp5_ASAP7_75t_L g2927 ( 
.A1(n_2911),
.A2(n_1992),
.B1(n_2290),
.B2(n_2295),
.Y(n_2927)
);

AOI22xp33_ASAP7_75t_SL g2928 ( 
.A1(n_2912),
.A2(n_2261),
.B1(n_2175),
.B2(n_2203),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2916),
.Y(n_2929)
);

OAI22xp5_ASAP7_75t_L g2930 ( 
.A1(n_2913),
.A2(n_1965),
.B1(n_1971),
.B2(n_1979),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2919),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2924),
.Y(n_2932)
);

AOI22xp5_ASAP7_75t_L g2933 ( 
.A1(n_2931),
.A2(n_2929),
.B1(n_2923),
.B2(n_2928),
.Y(n_2933)
);

AOI221xp5_ASAP7_75t_L g2934 ( 
.A1(n_2922),
.A2(n_2918),
.B1(n_2914),
.B2(n_2921),
.C(n_1994),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2925),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2927),
.B(n_2918),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_SL g2937 ( 
.A(n_2930),
.B(n_2261),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2926),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2924),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2932),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2939),
.Y(n_2941)
);

AOI22xp5_ASAP7_75t_L g2942 ( 
.A1(n_2933),
.A2(n_1965),
.B1(n_1971),
.B2(n_1979),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2938),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2935),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2944),
.B(n_2936),
.Y(n_2945)
);

OA22x2_ASAP7_75t_L g2946 ( 
.A1(n_2943),
.A2(n_2937),
.B1(n_2934),
.B2(n_2144),
.Y(n_2946)
);

AOI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2940),
.A2(n_2941),
.B1(n_2942),
.B2(n_2286),
.Y(n_2947)
);

NAND3xp33_ASAP7_75t_L g2948 ( 
.A(n_2944),
.B(n_2098),
.C(n_1971),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2945),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2948),
.Y(n_2950)
);

AOI22xp5_ASAP7_75t_L g2951 ( 
.A1(n_2949),
.A2(n_2946),
.B1(n_2947),
.B2(n_2261),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2950),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2952),
.Y(n_2953)
);

INVx3_ASAP7_75t_L g2954 ( 
.A(n_2951),
.Y(n_2954)
);

AOI22xp5_ASAP7_75t_L g2955 ( 
.A1(n_2953),
.A2(n_2259),
.B1(n_2166),
.B2(n_2175),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2955),
.Y(n_2956)
);

OAI22xp33_ASAP7_75t_L g2957 ( 
.A1(n_2956),
.A2(n_2954),
.B1(n_2259),
.B2(n_2245),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2957),
.Y(n_2958)
);

AOI221xp5_ASAP7_75t_L g2959 ( 
.A1(n_2958),
.A2(n_2954),
.B1(n_1979),
.B2(n_1994),
.C(n_1996),
.Y(n_2959)
);

AOI211xp5_ASAP7_75t_L g2960 ( 
.A1(n_2959),
.A2(n_2954),
.B(n_2286),
.C(n_2259),
.Y(n_2960)
);


endmodule