module fake_jpeg_2130_n_580 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_580);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_580;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_57),
.Y(n_134)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_63),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_64),
.Y(n_170)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_65),
.Y(n_213)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_18),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_68),
.B(n_84),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_69),
.B(n_89),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_70),
.Y(n_174)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_71),
.Y(n_162)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_72),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_73),
.Y(n_177)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_74),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_75),
.Y(n_209)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_77),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_35),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_78),
.A2(n_56),
.B1(n_55),
.B2(n_44),
.Y(n_136)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_81),
.Y(n_150)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_83),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_36),
.B(n_0),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx5_ASAP7_75t_SL g217 ( 
.A(n_85),
.Y(n_217)
);

BUFx4f_ASAP7_75t_SL g86 ( 
.A(n_37),
.Y(n_86)
);

BUFx4f_ASAP7_75t_SL g163 ( 
.A(n_86),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_35),
.B(n_0),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_5),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_90),
.Y(n_173)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_91),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_92),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_93),
.Y(n_190)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_95),
.Y(n_175)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_96),
.Y(n_179)
);

BUFx24_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

BUFx10_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_98),
.Y(n_207)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_100),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_35),
.B(n_3),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_102),
.B(n_5),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_105),
.Y(n_188)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_47),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_125),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_42),
.Y(n_113)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_20),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_116),
.Y(n_208)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_20),
.Y(n_118)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_118),
.Y(n_215)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_20),
.Y(n_119)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_47),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_120),
.B(n_121),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_22),
.Y(n_122)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_22),
.Y(n_123)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_47),
.Y(n_124)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_22),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_23),
.B(n_4),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_55),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_61),
.A2(n_56),
.B1(n_55),
.B2(n_50),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_127),
.A2(n_139),
.B1(n_143),
.B2(n_178),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_136),
.A2(n_160),
.B1(n_31),
.B2(n_6),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_23),
.B1(n_26),
.B2(n_52),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_141),
.B(n_144),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_26),
.B1(n_43),
.B2(n_52),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_84),
.B(n_45),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_146),
.A2(n_191),
.B(n_34),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_68),
.B(n_45),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_148),
.B(n_155),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_92),
.A2(n_51),
.B1(n_50),
.B2(n_49),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_154),
.A2(n_181),
.B1(n_189),
.B2(n_39),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_86),
.B(n_43),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_89),
.B(n_56),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_156),
.B(n_166),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_90),
.A2(n_50),
.B1(n_49),
.B2(n_44),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_49),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_63),
.A2(n_44),
.B1(n_54),
.B2(n_29),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_79),
.A2(n_51),
.B1(n_54),
.B2(n_29),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_108),
.B(n_34),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_183),
.B(n_192),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_64),
.A2(n_54),
.B1(n_53),
.B2(n_28),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_185),
.A2(n_194),
.B1(n_8),
.B2(n_9),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_85),
.A2(n_53),
.B1(n_28),
.B2(n_39),
.Y(n_189)
);

HAxp5_ASAP7_75t_SL g191 ( 
.A(n_97),
.B(n_47),
.CON(n_191),
.SN(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_109),
.B(n_33),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_70),
.A2(n_101),
.B1(n_75),
.B2(n_80),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_110),
.B(n_33),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_199),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_113),
.B(n_33),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_122),
.Y(n_203)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_73),
.B(n_53),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_206),
.B(n_212),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_120),
.B(n_38),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_216),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_124),
.B(n_38),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_153),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_218),
.Y(n_333)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_153),
.Y(n_219)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_219),
.Y(n_336)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_158),
.Y(n_220)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_220),
.Y(n_296)
);

NAND2xp33_ASAP7_75t_SL g222 ( 
.A(n_191),
.B(n_28),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_222),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_225),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_226),
.A2(n_244),
.B1(n_277),
.B2(n_279),
.Y(n_317)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_228),
.Y(n_348)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_157),
.Y(n_229)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_229),
.Y(n_303)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_131),
.Y(n_230)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_230),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

INVx6_ASAP7_75t_L g319 ( 
.A(n_231),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_217),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_232),
.B(n_256),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_233),
.Y(n_297)
);

A2O1A1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_149),
.A2(n_39),
.B(n_38),
.C(n_34),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_234),
.B(n_239),
.Y(n_312)
);

BUFx6f_ASAP7_75t_SL g237 ( 
.A(n_217),
.Y(n_237)
);

INVx13_ASAP7_75t_L g329 ( 
.A(n_237),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_127),
.A2(n_107),
.B1(n_103),
.B2(n_93),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_238),
.A2(n_255),
.B1(n_263),
.B2(n_275),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_168),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_240),
.B(n_249),
.Y(n_324)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_140),
.Y(n_241)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_159),
.Y(n_242)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_242),
.Y(n_313)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_243),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_134),
.A2(n_31),
.B1(n_29),
.B2(n_83),
.Y(n_244)
);

O2A1O1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_168),
.A2(n_189),
.B(n_154),
.C(n_215),
.Y(n_245)
);

O2A1O1Ixp33_ASAP7_75t_L g346 ( 
.A1(n_245),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_346)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_247),
.Y(n_335)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_248),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_128),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_137),
.Y(n_250)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_250),
.Y(n_316)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_251),
.Y(n_328)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_133),
.Y(n_252)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_252),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_200),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_253),
.B(n_257),
.Y(n_301)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_169),
.Y(n_254)
);

INVx8_ASAP7_75t_L g314 ( 
.A(n_254),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_178),
.A2(n_81),
.B1(n_31),
.B2(n_7),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_173),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_145),
.Y(n_258)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_258),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_162),
.B(n_5),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_259),
.B(n_264),
.Y(n_305)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_167),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_260),
.B(n_265),
.Y(n_347)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_175),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_261),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_185),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_204),
.B(n_6),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_137),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_193),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_266),
.B(n_267),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_135),
.B(n_6),
.Y(n_267)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_175),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_268),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_161),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_269),
.Y(n_326)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_151),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_270),
.B(n_271),
.Y(n_318)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_164),
.Y(n_271)
);

AND2x2_ASAP7_75t_SL g272 ( 
.A(n_129),
.B(n_138),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_208),
.C(n_211),
.Y(n_307)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_130),
.Y(n_273)
);

INVx8_ASAP7_75t_L g325 ( 
.A(n_273),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_207),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_274),
.B(n_276),
.Y(n_321)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_152),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_171),
.Y(n_277)
);

BUFx4f_ASAP7_75t_SL g278 ( 
.A(n_165),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_280),
.Y(n_299)
);

INVx11_ASAP7_75t_L g279 ( 
.A(n_165),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_172),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_201),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_281),
.A2(n_282),
.B1(n_284),
.B2(n_286),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_213),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_173),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_291),
.Y(n_295)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_210),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_202),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_179),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_147),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_187),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_213),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_187),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_161),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_293),
.B(n_182),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_236),
.A2(n_181),
.B1(n_198),
.B2(n_176),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_300),
.A2(n_337),
.B1(n_343),
.B2(n_346),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_226),
.A2(n_198),
.B1(n_142),
.B2(n_190),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_302),
.A2(n_323),
.B1(n_341),
.B2(n_331),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_307),
.B(n_291),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_163),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_340),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_L g323 ( 
.A1(n_245),
.A2(n_150),
.B1(n_190),
.B2(n_184),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_222),
.A2(n_165),
.B(n_163),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_331),
.Y(n_389)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_332),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_246),
.B(n_142),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_344),
.Y(n_350)
);

OAI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_225),
.A2(n_182),
.B1(n_176),
.B2(n_177),
.Y(n_337)
);

FAx1_ASAP7_75t_L g338 ( 
.A(n_292),
.B(n_130),
.CI(n_184),
.CON(n_338),
.SN(n_338)
);

A2O1A1Ixp33_ASAP7_75t_L g357 ( 
.A1(n_338),
.A2(n_244),
.B(n_232),
.C(n_237),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_262),
.B(n_209),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_227),
.A2(n_150),
.B1(n_177),
.B2(n_174),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_234),
.A2(n_209),
.B1(n_174),
.B2(n_170),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_235),
.B(n_170),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_333),
.Y(n_349)
);

INVx6_ASAP7_75t_L g401 ( 
.A(n_349),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_324),
.B(n_223),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_351),
.B(n_378),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_272),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_352),
.B(n_355),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_354),
.B(n_368),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_344),
.B(n_272),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_303),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_356),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_357),
.A2(n_332),
.B(n_327),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_221),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_358),
.B(n_372),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_338),
.A2(n_289),
.B1(n_260),
.B2(n_266),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_359),
.A2(n_365),
.B1(n_370),
.B2(n_323),
.Y(n_395)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_303),
.Y(n_361)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_361),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_336),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_362),
.Y(n_424)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_306),
.Y(n_364)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_364),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_338),
.A2(n_252),
.B1(n_230),
.B2(n_254),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_298),
.A2(n_261),
.B1(n_268),
.B2(n_273),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_366),
.A2(n_326),
.B(n_304),
.Y(n_408)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_306),
.Y(n_367)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_367),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_311),
.B(n_224),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_308),
.B(n_305),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_369),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_312),
.B(n_293),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_371),
.B(n_386),
.C(n_310),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_309),
.B(n_281),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_319),
.Y(n_373)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_373),
.Y(n_418)
);

AOI32xp33_ASAP7_75t_L g374 ( 
.A1(n_295),
.A2(n_276),
.A3(n_243),
.B1(n_290),
.B2(n_265),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_374),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_295),
.B(n_269),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_375),
.B(n_376),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_307),
.B(n_231),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_301),
.Y(n_377)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_377),
.Y(n_422)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_313),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_313),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_379),
.B(n_380),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_299),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_341),
.A2(n_219),
.B1(n_218),
.B2(n_287),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_381),
.A2(n_390),
.B1(n_326),
.B2(n_310),
.Y(n_396)
);

BUFx5_ASAP7_75t_L g382 ( 
.A(n_348),
.Y(n_382)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_294),
.B(n_250),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_383),
.B(n_384),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_294),
.B(n_278),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_385),
.A2(n_388),
.B1(n_336),
.B2(n_347),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_298),
.B(n_288),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_294),
.B(n_278),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_387),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_345),
.A2(n_279),
.B1(n_11),
.B2(n_12),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_345),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_328),
.B(n_13),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_391),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_389),
.A2(n_357),
.B(n_387),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_392),
.A2(n_414),
.B(n_425),
.Y(n_456)
);

A2O1A1Ixp33_ASAP7_75t_L g393 ( 
.A1(n_389),
.A2(n_346),
.B(n_302),
.C(n_318),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_393),
.B(n_366),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_395),
.A2(n_423),
.B1(n_426),
.B2(n_360),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_396),
.A2(n_398),
.B1(n_371),
.B2(n_390),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_370),
.A2(n_317),
.B1(n_342),
.B2(n_299),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_362),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_400),
.B(n_413),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_404),
.A2(n_392),
.B1(n_414),
.B2(n_409),
.Y(n_448)
);

INVxp33_ASAP7_75t_SL g436 ( 
.A(n_408),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_409),
.B(n_363),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_372),
.Y(n_413)
);

FAx1_ASAP7_75t_L g414 ( 
.A(n_359),
.B(n_304),
.CI(n_321),
.CON(n_414),
.SN(n_414)
);

OAI32xp33_ASAP7_75t_L g421 ( 
.A1(n_350),
.A2(n_339),
.A3(n_328),
.B1(n_330),
.B2(n_315),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_421),
.B(n_350),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_365),
.A2(n_384),
.B1(n_353),
.B2(n_383),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_353),
.A2(n_339),
.B(n_347),
.Y(n_425)
);

BUFx5_ASAP7_75t_L g427 ( 
.A(n_414),
.Y(n_427)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_427),
.Y(n_464)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_399),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_428),
.Y(n_481)
);

NAND3xp33_ASAP7_75t_L g429 ( 
.A(n_394),
.B(n_354),
.C(n_358),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_429),
.B(n_444),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_424),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_430),
.B(n_432),
.Y(n_484)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_410),
.Y(n_433)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_433),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_425),
.Y(n_434)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_434),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_413),
.B(n_355),
.Y(n_435)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_435),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_437),
.A2(n_447),
.B1(n_412),
.B2(n_396),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_421),
.B(n_376),
.Y(n_438)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_438),
.Y(n_483)
);

AO22x1_ASAP7_75t_SL g439 ( 
.A1(n_414),
.A2(n_360),
.B1(n_354),
.B2(n_386),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_443),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_397),
.B(n_363),
.C(n_368),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_440),
.B(n_422),
.C(n_394),
.Y(n_469)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_410),
.Y(n_441)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_441),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_451),
.Y(n_466)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_411),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_405),
.B(n_352),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_445),
.A2(n_446),
.B1(n_448),
.B2(n_458),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_417),
.A2(n_381),
.B1(n_361),
.B2(n_356),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_416),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_449),
.A2(n_450),
.B(n_403),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_422),
.B(n_297),
.Y(n_450)
);

OAI32xp33_ASAP7_75t_L g451 ( 
.A1(n_420),
.A2(n_416),
.A3(n_423),
.B1(n_419),
.B2(n_393),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_395),
.A2(n_373),
.B1(n_319),
.B2(n_314),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_452),
.A2(n_453),
.B1(n_454),
.B2(n_455),
.Y(n_467)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_411),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_404),
.A2(n_314),
.B1(n_349),
.B2(n_325),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_399),
.Y(n_455)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_418),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_457),
.A2(n_406),
.B1(n_418),
.B2(n_400),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_398),
.A2(n_325),
.B1(n_385),
.B2(n_333),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_459),
.A2(n_460),
.B1(n_465),
.B2(n_479),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_445),
.A2(n_407),
.B1(n_405),
.B2(n_420),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_440),
.B(n_397),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_463),
.B(n_469),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_438),
.A2(n_407),
.B1(n_412),
.B2(n_402),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_468),
.B(n_487),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_442),
.B(n_444),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_472),
.B(n_473),
.C(n_474),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_434),
.B(n_315),
.C(n_330),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_432),
.B(n_408),
.Y(n_474)
);

FAx1_ASAP7_75t_SL g475 ( 
.A(n_435),
.B(n_402),
.CI(n_406),
.CON(n_475),
.SN(n_475)
);

FAx1_ASAP7_75t_SL g506 ( 
.A(n_475),
.B(n_453),
.CI(n_441),
.CON(n_506),
.SN(n_506)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_476),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_439),
.B(n_347),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_477),
.B(n_482),
.C(n_485),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_436),
.A2(n_415),
.B1(n_333),
.B2(n_401),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_439),
.B(n_297),
.C(n_316),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_449),
.B(n_316),
.C(n_348),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_456),
.B(n_296),
.C(n_320),
.Y(n_487)
);

AOI21x1_ASAP7_75t_L g488 ( 
.A1(n_464),
.A2(n_431),
.B(n_456),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_488),
.A2(n_499),
.B(n_504),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_SL g489 ( 
.A(n_466),
.B(n_451),
.Y(n_489)
);

MAJx2_ASAP7_75t_L g521 ( 
.A(n_489),
.B(n_498),
.C(n_462),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_431),
.Y(n_492)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_492),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_459),
.A2(n_483),
.B1(n_465),
.B2(n_460),
.Y(n_494)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_494),
.Y(n_511)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_471),
.Y(n_495)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_495),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_481),
.B(n_428),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_496),
.B(n_502),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_466),
.B(n_427),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_461),
.A2(n_454),
.B(n_458),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_486),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_500),
.A2(n_503),
.B1(n_505),
.B2(n_506),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_455),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_484),
.A2(n_446),
.B1(n_430),
.B2(n_443),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_462),
.A2(n_452),
.B(n_457),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_473),
.Y(n_505)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_479),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_510),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_485),
.B(n_433),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_509),
.B(n_475),
.Y(n_527)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_467),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_510),
.A2(n_493),
.B1(n_478),
.B2(n_499),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_514),
.A2(n_490),
.B1(n_494),
.B2(n_503),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_472),
.C(n_463),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_520),
.C(n_526),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_491),
.B(n_482),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_518),
.B(n_521),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_505),
.B(n_469),
.Y(n_519)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_519),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_507),
.B(n_487),
.C(n_470),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_491),
.B(n_474),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_523),
.B(n_525),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_501),
.B(n_477),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_501),
.B(n_475),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_527),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_512),
.A2(n_497),
.B(n_488),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_529),
.B(n_536),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_520),
.B(n_509),
.C(n_493),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_530),
.B(n_535),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_531),
.A2(n_532),
.B1(n_335),
.B2(n_382),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_522),
.A2(n_490),
.B1(n_508),
.B2(n_492),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_514),
.A2(n_502),
.B1(n_504),
.B2(n_500),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_533),
.A2(n_542),
.B1(n_517),
.B2(n_511),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_518),
.B(n_498),
.C(n_489),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_523),
.B(n_496),
.C(n_495),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_516),
.B(n_415),
.C(n_506),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_537),
.B(n_521),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_512),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_SL g548 ( 
.A1(n_539),
.A2(n_515),
.B1(n_322),
.B2(n_335),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_526),
.A2(n_527),
.B(n_525),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_543),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_532),
.A2(n_513),
.B(n_511),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g562 ( 
.A1(n_544),
.A2(n_537),
.B(n_535),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_545),
.B(n_552),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_540),
.A2(n_515),
.B1(n_506),
.B2(n_524),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_547),
.B(n_548),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_536),
.B(n_401),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_549),
.B(n_551),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_541),
.A2(n_401),
.B1(n_322),
.B2(n_296),
.Y(n_551)
);

CKINVDCx16_ASAP7_75t_R g552 ( 
.A(n_530),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_553),
.B(n_554),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_541),
.A2(n_329),
.B1(n_14),
.B2(n_16),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_550),
.B(n_538),
.C(n_528),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_556),
.B(n_561),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_545),
.B(n_528),
.C(n_538),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_562),
.B(n_546),
.Y(n_564)
);

NOR2x1_ASAP7_75t_L g563 ( 
.A(n_547),
.B(n_534),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_563),
.A2(n_534),
.B(n_544),
.Y(n_565)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_564),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g572 ( 
.A1(n_565),
.A2(n_566),
.B(n_567),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_556),
.B(n_549),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_555),
.A2(n_560),
.B(n_563),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_560),
.B(n_559),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_569),
.A2(n_558),
.B(n_557),
.Y(n_570)
);

AOI21xp33_ASAP7_75t_L g574 ( 
.A1(n_570),
.A2(n_564),
.B(n_551),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_568),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_571),
.B(n_553),
.Y(n_575)
);

AOI21x1_ASAP7_75t_L g576 ( 
.A1(n_574),
.A2(n_575),
.B(n_572),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_576),
.B(n_573),
.Y(n_577)
);

O2A1O1Ixp33_ASAP7_75t_SL g578 ( 
.A1(n_577),
.A2(n_554),
.B(n_329),
.C(n_14),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_14),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_579),
.Y(n_580)
);


endmodule