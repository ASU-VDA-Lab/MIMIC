module fake_netlist_5_1793_n_1861 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1861);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1861;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_15),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_121),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_107),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_113),
.Y(n_188)
);

CKINVDCx11_ASAP7_75t_R g189 ( 
.A(n_111),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_118),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_183),
.Y(n_191)
);

BUFx2_ASAP7_75t_R g192 ( 
.A(n_34),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_77),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_132),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_136),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_25),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_79),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_102),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_109),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_39),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_70),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_58),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_96),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_43),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_74),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_6),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_27),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_141),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_42),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_40),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_29),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_150),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_112),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_68),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_9),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_127),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_184),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_148),
.Y(n_224)
);

BUFx8_ASAP7_75t_SL g225 ( 
.A(n_126),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_133),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_147),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_43),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_23),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_8),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_91),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_20),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_83),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_163),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_116),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_23),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_122),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_168),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_39),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g240 ( 
.A(n_87),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_138),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_28),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_101),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_120),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_50),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_8),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_30),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_131),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_181),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_90),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_62),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_178),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_26),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_128),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_78),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_86),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_12),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_33),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_28),
.Y(n_259)
);

BUFx8_ASAP7_75t_SL g260 ( 
.A(n_6),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_169),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_19),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_58),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_125),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_40),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_24),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_93),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_81),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_57),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_21),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_100),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_129),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_73),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_171),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_26),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_153),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_10),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_47),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_108),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_155),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_145),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_173),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_95),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_63),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_104),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_166),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_1),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_46),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_18),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_160),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_165),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_106),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_5),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_162),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_51),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_142),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_179),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_16),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_82),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_34),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_22),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_156),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_59),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_66),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_72),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_16),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_161),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_27),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_22),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_174),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_146),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_33),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_167),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_17),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_19),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_59),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_50),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_180),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_44),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_119),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_17),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_85),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_80),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_56),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_44),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_61),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_3),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_177),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_14),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_31),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_105),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_10),
.Y(n_332)
);

BUFx10_ASAP7_75t_L g333 ( 
.A(n_2),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_18),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_139),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_31),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_158),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_36),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_71),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_60),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_149),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_24),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_92),
.Y(n_343)
);

BUFx5_ASAP7_75t_L g344 ( 
.A(n_41),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_25),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_130),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_144),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_94),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_14),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_3),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_76),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_38),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_2),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_115),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_20),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_97),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_46),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_21),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_124),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_15),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_57),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_37),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_53),
.Y(n_363)
);

BUFx10_ASAP7_75t_L g364 ( 
.A(n_123),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_65),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_29),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_344),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_187),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_344),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_312),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_344),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_344),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_239),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_344),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_225),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_344),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_247),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_344),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_260),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_344),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_212),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_201),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_189),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_212),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_212),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_222),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_212),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_295),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_200),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_223),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_212),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_270),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_200),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_270),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_284),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_300),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_226),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_300),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_358),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_358),
.Y(n_400)
);

INVxp33_ASAP7_75t_L g401 ( 
.A(n_210),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_215),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_227),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_233),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_221),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_230),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_259),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_333),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_234),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_235),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_243),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_262),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_241),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_265),
.Y(n_414)
);

INVxp33_ASAP7_75t_SL g415 ( 
.A(n_204),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_229),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_197),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_266),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_275),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_209),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_249),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_278),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_289),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_293),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_333),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_339),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_301),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_197),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_306),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_308),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_251),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_316),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_244),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_185),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_333),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_324),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_213),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_330),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_342),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_349),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_224),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_273),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_362),
.Y(n_443)
);

INVxp33_ASAP7_75t_SL g444 ( 
.A(n_204),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_294),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_318),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_224),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_196),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_272),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_272),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_196),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_252),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_194),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_232),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_351),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_351),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_198),
.Y(n_457)
);

INVxp33_ASAP7_75t_SL g458 ( 
.A(n_207),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_369),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_453),
.B(n_268),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_369),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_381),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_370),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_386),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_381),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_384),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_397),
.B(n_268),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_368),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_384),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_373),
.A2(n_363),
.B1(n_236),
.B2(n_298),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_385),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_385),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_387),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_L g474 ( 
.A(n_404),
.B(n_207),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_387),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_428),
.B(n_218),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_391),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_434),
.B(n_218),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_382),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_367),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_391),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_367),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_371),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_409),
.B(n_328),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_371),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_457),
.B(n_328),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_372),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_372),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_374),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_388),
.A2(n_361),
.B1(n_360),
.B2(n_357),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_374),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_410),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_376),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_376),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_389),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_378),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_417),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_408),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_457),
.B(n_202),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_378),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_R g501 ( 
.A(n_375),
.B(n_331),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_413),
.B(n_205),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_437),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_441),
.B(n_218),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_380),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_380),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_395),
.B(n_383),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_412),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_390),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_412),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_447),
.B(n_250),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_421),
.B(n_206),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_423),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_425),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_423),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_393),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_448),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_448),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_451),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_431),
.B(n_208),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_451),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_455),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_449),
.B(n_450),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_L g524 ( 
.A(n_452),
.B(n_216),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_455),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_417),
.B(n_231),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_392),
.B(n_250),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_392),
.B(n_250),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_394),
.B(n_274),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_456),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_420),
.B(n_238),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_456),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_402),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_426),
.B(n_248),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_377),
.A2(n_288),
.B1(n_314),
.B2(n_216),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_402),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_405),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_468),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_501),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_459),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_497),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_482),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_523),
.B(n_305),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_461),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_467),
.B(n_415),
.Y(n_545)
);

BUFx4f_ASAP7_75t_L g546 ( 
.A(n_485),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_461),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_485),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_459),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_523),
.B(n_458),
.Y(n_550)
);

OR2x6_ASAP7_75t_L g551 ( 
.A(n_497),
.B(n_440),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_523),
.B(n_460),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_482),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_461),
.Y(n_554)
);

NOR2x1p5_ASAP7_75t_L g555 ( 
.A(n_464),
.B(n_379),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_498),
.B(n_416),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_459),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_503),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_470),
.A2(n_355),
.B1(n_357),
.B2(n_353),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_461),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_484),
.B(n_444),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_480),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_460),
.A2(n_401),
.B1(n_320),
.B2(n_237),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_488),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_480),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_480),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_523),
.B(n_255),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_483),
.Y(n_568)
);

NAND3xp33_ASAP7_75t_L g569 ( 
.A(n_460),
.B(n_406),
.C(n_405),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_502),
.B(n_454),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_483),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_497),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_476),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_459),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_492),
.B(n_435),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_483),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_487),
.Y(n_577)
);

INVx5_ASAP7_75t_L g578 ( 
.A(n_485),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_498),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_487),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_459),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_488),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_459),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_485),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_512),
.B(n_394),
.Y(n_585)
);

NAND3xp33_ASAP7_75t_L g586 ( 
.A(n_474),
.B(n_398),
.C(n_396),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_485),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_487),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_494),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_489),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_520),
.B(n_396),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_494),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_494),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_476),
.B(n_274),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_489),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_460),
.B(n_261),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_485),
.Y(n_597)
);

AND2x6_ASAP7_75t_L g598 ( 
.A(n_491),
.B(n_237),
.Y(n_598)
);

INVxp33_ASAP7_75t_SL g599 ( 
.A(n_463),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_491),
.B(n_264),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_L g601 ( 
.A(n_531),
.B(n_237),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_500),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_496),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_500),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_496),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_505),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_499),
.A2(n_237),
.B1(n_320),
.B2(n_398),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_505),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_506),
.B(n_271),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_493),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_514),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_500),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_506),
.Y(n_613)
);

AO21x2_ASAP7_75t_L g614 ( 
.A1(n_534),
.A2(n_256),
.B(n_254),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_462),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_504),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_462),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_493),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_479),
.Y(n_619)
);

BUFx4f_ASAP7_75t_L g620 ( 
.A(n_493),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_504),
.B(n_279),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_511),
.B(n_280),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_511),
.B(n_486),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_527),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_495),
.B(n_399),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_537),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_493),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_493),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_499),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_499),
.A2(n_237),
.B1(n_320),
.B2(n_399),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_507),
.B(n_400),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_537),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_470),
.A2(n_338),
.B1(n_217),
.B2(n_345),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_516),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_465),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_493),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_537),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_499),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_465),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_466),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_537),
.Y(n_641)
);

BUFx2_ASAP7_75t_L g642 ( 
.A(n_527),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_537),
.Y(n_643)
);

CKINVDCx14_ASAP7_75t_R g644 ( 
.A(n_509),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_537),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_486),
.B(n_281),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_466),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_472),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_472),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_469),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_475),
.Y(n_651)
);

INVxp67_ASAP7_75t_SL g652 ( 
.A(n_526),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_475),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_535),
.A2(n_338),
.B1(n_217),
.B2(n_345),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_535),
.A2(n_350),
.B1(n_352),
.B2(n_353),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_477),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_477),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_481),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_481),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_528),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_469),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_517),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_486),
.B(n_282),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_469),
.Y(n_664)
);

BUFx10_ASAP7_75t_L g665 ( 
.A(n_486),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_533),
.Y(n_666)
);

INVx5_ASAP7_75t_L g667 ( 
.A(n_469),
.Y(n_667)
);

INVxp67_ASAP7_75t_SL g668 ( 
.A(n_469),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_529),
.B(n_286),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_533),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_529),
.B(n_291),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_524),
.B(n_400),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_517),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_521),
.B(n_292),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_517),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_533),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_478),
.B(n_490),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_503),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_536),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_518),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_519),
.B(n_406),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_518),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_490),
.B(n_446),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_519),
.B(n_407),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_518),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_522),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_536),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_530),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_677),
.A2(n_321),
.B1(n_320),
.B2(n_322),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_552),
.A2(n_442),
.B1(n_403),
.B2(n_411),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_573),
.B(n_186),
.Y(n_691)
);

NOR3xp33_ASAP7_75t_L g692 ( 
.A(n_683),
.B(n_240),
.C(n_191),
.Y(n_692)
);

NOR2xp67_ASAP7_75t_L g693 ( 
.A(n_539),
.B(n_530),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_652),
.B(n_521),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_687),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_585),
.B(n_521),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_615),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_573),
.B(n_186),
.Y(n_698)
);

INVxp67_ASAP7_75t_SL g699 ( 
.A(n_597),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_617),
.Y(n_700)
);

O2A1O1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_616),
.A2(n_532),
.B(n_436),
.C(n_432),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_616),
.B(n_188),
.Y(n_702)
);

NOR2x1p5_ASAP7_75t_L g703 ( 
.A(n_539),
.B(n_350),
.Y(n_703)
);

AND2x2_ASAP7_75t_SL g704 ( 
.A(n_563),
.B(n_320),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_624),
.B(n_660),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_687),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_570),
.B(n_188),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_591),
.B(n_521),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_660),
.B(n_525),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_642),
.B(n_433),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_681),
.Y(n_711)
);

OAI21xp33_ASAP7_75t_L g712 ( 
.A1(n_625),
.A2(n_414),
.B(n_407),
.Y(n_712)
);

BUFx5_ASAP7_75t_L g713 ( 
.A(n_626),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_629),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_629),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_556),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_642),
.B(n_190),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_634),
.B(n_445),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_681),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_617),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_635),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_614),
.A2(n_310),
.B1(n_299),
.B2(n_267),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_679),
.B(n_525),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_679),
.B(n_522),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_L g725 ( 
.A1(n_623),
.A2(n_290),
.B(n_283),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_635),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_639),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_545),
.B(n_193),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_542),
.B(n_522),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_546),
.A2(n_532),
.B(n_510),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_542),
.B(n_522),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_561),
.A2(n_304),
.B1(n_307),
.B2(n_311),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_550),
.B(n_193),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_665),
.B(n_195),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_614),
.A2(n_296),
.B1(n_297),
.B2(n_302),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_553),
.B(n_522),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_665),
.B(n_543),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_564),
.B(n_582),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_564),
.B(n_522),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_614),
.A2(n_582),
.B1(n_595),
.B2(n_590),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_639),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_638),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_672),
.B(n_195),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_640),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_590),
.B(n_469),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_638),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_621),
.B(n_199),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_684),
.Y(n_748)
);

A2O1A1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_569),
.A2(n_515),
.B(n_513),
.C(n_510),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_665),
.B(n_199),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_644),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_595),
.B(n_471),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_640),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_684),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_551),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_603),
.A2(n_352),
.B1(n_360),
.B2(n_355),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_647),
.Y(n_757)
);

OR2x6_ASAP7_75t_L g758 ( 
.A(n_556),
.B(n_414),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_688),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_622),
.B(n_203),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_603),
.B(n_471),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_567),
.A2(n_313),
.B1(n_323),
.B2(n_326),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_605),
.B(n_606),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_669),
.B(n_203),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_541),
.B(n_211),
.Y(n_765)
);

OAI21xp5_ASAP7_75t_L g766 ( 
.A1(n_605),
.A2(n_515),
.B(n_513),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_551),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_671),
.B(n_541),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_594),
.B(n_211),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_688),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_596),
.A2(n_663),
.B1(n_646),
.B2(n_600),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_606),
.A2(n_418),
.B1(n_443),
.B2(n_439),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_608),
.B(n_471),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_SL g774 ( 
.A1(n_634),
.A2(n_274),
.B1(n_285),
.B2(n_364),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_572),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_608),
.B(n_471),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_613),
.B(n_471),
.Y(n_777)
);

CKINVDCx11_ASAP7_75t_R g778 ( 
.A(n_538),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_572),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_597),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_609),
.B(n_214),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_613),
.A2(n_418),
.B1(n_443),
.B2(n_439),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_647),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_569),
.B(n_214),
.Y(n_784)
);

BUFx8_ASAP7_75t_L g785 ( 
.A(n_579),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_648),
.B(n_471),
.Y(n_786)
);

NOR3xp33_ASAP7_75t_L g787 ( 
.A(n_575),
.B(n_419),
.C(n_438),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_551),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_649),
.Y(n_789)
);

NAND2xp33_ASAP7_75t_L g790 ( 
.A(n_607),
.B(n_335),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_630),
.A2(n_419),
.B1(n_438),
.B2(n_436),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_579),
.B(n_422),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_648),
.B(n_473),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_649),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_653),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_611),
.B(n_219),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_558),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_651),
.B(n_473),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_601),
.A2(n_422),
.B1(n_424),
.B2(n_432),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_651),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_601),
.A2(n_424),
.B1(n_427),
.B2(n_430),
.Y(n_801)
);

NAND2xp33_ASAP7_75t_L g802 ( 
.A(n_674),
.B(n_337),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_631),
.A2(n_220),
.B1(n_276),
.B2(n_340),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_658),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_611),
.B(n_340),
.Y(n_805)
);

NOR2xp67_ASAP7_75t_L g806 ( 
.A(n_558),
.B(n_508),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_653),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_586),
.B(n_341),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_658),
.B(n_473),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_551),
.B(n_631),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_656),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_656),
.B(n_473),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_631),
.B(n_341),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_631),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_559),
.B(n_343),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_633),
.B(n_346),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_657),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_659),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_659),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_666),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_587),
.B(n_540),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_662),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_662),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_633),
.B(n_346),
.Y(n_824)
);

INVxp33_ASAP7_75t_L g825 ( 
.A(n_654),
.Y(n_825)
);

OR2x2_ASAP7_75t_L g826 ( 
.A(n_619),
.B(n_427),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_666),
.A2(n_347),
.B1(n_348),
.B2(n_354),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_673),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_599),
.B(n_347),
.Y(n_829)
);

OAI221xp5_ASAP7_75t_L g830 ( 
.A1(n_654),
.A2(n_429),
.B1(n_430),
.B2(n_508),
.C(n_319),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_599),
.B(n_348),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_597),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_678),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_587),
.B(n_473),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_673),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_675),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_675),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_670),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_678),
.B(n_354),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_587),
.B(n_473),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_680),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_555),
.A2(n_365),
.B1(n_359),
.B2(n_356),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_540),
.B(n_356),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_540),
.B(n_359),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_555),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_670),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_655),
.B(n_429),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_626),
.B(n_365),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_676),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_557),
.B(n_228),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_655),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_557),
.B(n_242),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_632),
.B(n_285),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_715),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_775),
.B(n_632),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_697),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_826),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_710),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_SL g859 ( 
.A1(n_825),
.A2(n_309),
.B1(n_245),
.B2(n_246),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_775),
.B(n_637),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_715),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_697),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_785),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_771),
.B(n_696),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_700),
.Y(n_865)
);

AOI221xp5_ASAP7_75t_L g866 ( 
.A1(n_824),
.A2(n_317),
.B1(n_253),
.B2(n_257),
.C(n_258),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_708),
.B(n_676),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_738),
.B(n_562),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_707),
.A2(n_668),
.B1(n_637),
.B2(n_645),
.Y(n_869)
);

AO22x1_ASAP7_75t_L g870 ( 
.A1(n_824),
.A2(n_315),
.B1(n_263),
.B2(n_269),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_707),
.A2(n_645),
.B1(n_643),
.B2(n_557),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_SL g872 ( 
.A1(n_704),
.A2(n_733),
.B1(n_813),
.B2(n_743),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_785),
.Y(n_873)
);

NOR2xp67_ASAP7_75t_L g874 ( 
.A(n_716),
.B(n_686),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_704),
.A2(n_588),
.B1(n_580),
.B2(n_589),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_700),
.Y(n_876)
);

BUFx5_ASAP7_75t_L g877 ( 
.A(n_820),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_720),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_689),
.A2(n_735),
.B1(n_722),
.B2(n_851),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_720),
.Y(n_880)
);

OR2x6_ASAP7_75t_L g881 ( 
.A(n_718),
.B(n_192),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_725),
.A2(n_588),
.B1(n_580),
.B2(n_589),
.Y(n_882)
);

NOR2x1_ASAP7_75t_L g883 ( 
.A(n_703),
.B(n_643),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_692),
.A2(n_571),
.B1(n_592),
.B2(n_602),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_778),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_743),
.B(n_581),
.Y(n_886)
);

OR2x6_ASAP7_75t_L g887 ( 
.A(n_755),
.B(n_686),
.Y(n_887)
);

INVx1_ASAP7_75t_SL g888 ( 
.A(n_792),
.Y(n_888)
);

AO22x1_ASAP7_75t_L g889 ( 
.A1(n_813),
.A2(n_287),
.B1(n_277),
.B2(n_366),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_833),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_763),
.B(n_562),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_715),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_695),
.B(n_565),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_758),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_751),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_728),
.B(n_548),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_721),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_733),
.A2(n_581),
.B(n_571),
.C(n_576),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_706),
.B(n_565),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_715),
.B(n_546),
.Y(n_900)
);

INVx5_ASAP7_75t_L g901 ( 
.A(n_758),
.Y(n_901)
);

INVx5_ASAP7_75t_L g902 ( 
.A(n_758),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_747),
.A2(n_584),
.B1(n_618),
.B2(n_548),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_742),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_767),
.B(n_788),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_742),
.B(n_546),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_742),
.B(n_620),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_742),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_R g909 ( 
.A(n_845),
.B(n_664),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_759),
.B(n_566),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_847),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_796),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_711),
.B(n_664),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_765),
.B(n_584),
.Y(n_914)
);

INVx5_ASAP7_75t_L g915 ( 
.A(n_780),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_726),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_726),
.Y(n_917)
);

AND2x4_ASAP7_75t_SL g918 ( 
.A(n_797),
.B(n_746),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_746),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_737),
.A2(n_584),
.B1(n_618),
.B2(n_664),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_781),
.A2(n_554),
.B1(n_560),
.B2(n_547),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_SL g922 ( 
.A1(n_774),
.A2(n_329),
.B1(n_303),
.B2(n_325),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_765),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_727),
.Y(n_924)
);

OR2x6_ASAP7_75t_L g925 ( 
.A(n_814),
.B(n_544),
.Y(n_925)
);

INVx5_ASAP7_75t_L g926 ( 
.A(n_780),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_805),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_727),
.Y(n_928)
);

INVxp67_ASAP7_75t_SL g929 ( 
.A(n_714),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_746),
.B(n_620),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_717),
.B(n_327),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_741),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_746),
.Y(n_933)
);

NAND2xp33_ASAP7_75t_SL g934 ( 
.A(n_689),
.B(n_332),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_690),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_719),
.B(n_544),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_781),
.B(n_566),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_693),
.B(n_620),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_779),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_722),
.A2(n_334),
.B1(n_336),
.B2(n_568),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_717),
.B(n_285),
.Y(n_941)
);

NAND3xp33_ASAP7_75t_SL g942 ( 
.A(n_803),
.B(n_842),
.C(n_732),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_714),
.B(n_641),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_741),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_744),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_770),
.B(n_568),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_779),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_744),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_800),
.B(n_576),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_753),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_753),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_804),
.B(n_577),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_748),
.B(n_680),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_735),
.A2(n_592),
.B1(n_593),
.B2(n_577),
.Y(n_954)
);

BUFx2_ASAP7_75t_SL g955 ( 
.A(n_806),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_757),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_754),
.B(n_593),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_768),
.B(n_549),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_779),
.B(n_547),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_757),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_810),
.A2(n_705),
.B1(n_769),
.B2(n_760),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_783),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_783),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_779),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_789),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_789),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_810),
.A2(n_554),
.B1(n_560),
.B2(n_604),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_807),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_740),
.B(n_602),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_815),
.B(n_816),
.Y(n_970)
);

NOR3xp33_ASAP7_75t_SL g971 ( 
.A(n_830),
.B(n_364),
.C(n_1),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_740),
.B(n_604),
.Y(n_972)
);

AND2x6_ASAP7_75t_L g973 ( 
.A(n_780),
.B(n_612),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_794),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_756),
.B(n_682),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_705),
.A2(n_627),
.B1(n_597),
.B2(n_610),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_709),
.B(n_685),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_807),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_794),
.Y(n_979)
);

BUFx12f_ASAP7_75t_SL g980 ( 
.A(n_780),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_817),
.A2(n_641),
.B1(n_597),
.B2(n_610),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_R g982 ( 
.A(n_811),
.B(n_790),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_818),
.A2(n_641),
.B1(n_610),
.B2(n_627),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_762),
.B(n_641),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_795),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_787),
.B(n_641),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_795),
.Y(n_987)
);

NAND2x1_ASAP7_75t_L g988 ( 
.A(n_832),
.B(n_610),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_819),
.A2(n_811),
.B1(n_838),
.B2(n_849),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_694),
.A2(n_549),
.B(n_574),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_691),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_850),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_R g993 ( 
.A(n_802),
.B(n_88),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_846),
.Y(n_994)
);

BUFx4f_ASAP7_75t_L g995 ( 
.A(n_832),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_822),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_698),
.B(n_627),
.Y(n_997)
);

NOR2xp67_ASAP7_75t_L g998 ( 
.A(n_852),
.B(n_89),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_829),
.B(n_549),
.Y(n_999)
);

NOR2x1p5_ASAP7_75t_L g1000 ( 
.A(n_843),
.B(n_650),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_723),
.B(n_574),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_699),
.B(n_574),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_822),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_831),
.B(n_0),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_764),
.B(n_627),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_823),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_844),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_713),
.B(n_574),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_821),
.A2(n_724),
.B(n_840),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_848),
.A2(n_0),
.B(n_4),
.C(n_5),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_713),
.B(n_574),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_828),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_839),
.B(n_583),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_827),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_756),
.B(n_4),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_834),
.A2(n_583),
.B(n_627),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_832),
.B(n_628),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_835),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_848),
.A2(n_628),
.B1(n_636),
.B2(n_610),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_835),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_702),
.B(n_583),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_832),
.B(n_628),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_791),
.A2(n_636),
.B1(n_628),
.B2(n_583),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_734),
.B(n_583),
.Y(n_1024)
);

AND2x6_ASAP7_75t_L g1025 ( 
.A(n_836),
.B(n_636),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_808),
.Y(n_1026)
);

AO22x1_ASAP7_75t_L g1027 ( 
.A1(n_766),
.A2(n_598),
.B1(n_628),
.B2(n_636),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_750),
.B(n_636),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_853),
.B(n_650),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_841),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_837),
.Y(n_1031)
);

AND2x6_ASAP7_75t_SL g1032 ( 
.A(n_745),
.B(n_7),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_970),
.A2(n_701),
.B(n_853),
.C(n_784),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_872),
.A2(n_712),
.B(n_731),
.C(n_736),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_854),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_996),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_888),
.B(n_749),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_964),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_995),
.A2(n_739),
.B(n_729),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_923),
.B(n_841),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_1003),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_895),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_R g1043 ( 
.A(n_980),
.B(n_837),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_879),
.A2(n_776),
.B(n_809),
.C(n_777),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_R g1045 ( 
.A(n_935),
.B(n_773),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_953),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_856),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_862),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_914),
.B(n_713),
.Y(n_1049)
);

AOI222xp33_ASAP7_75t_L g1050 ( 
.A1(n_1015),
.A2(n_772),
.B1(n_782),
.B2(n_791),
.C1(n_799),
.C2(n_801),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_854),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_918),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_879),
.A2(n_761),
.B(n_752),
.C(n_798),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_888),
.B(n_713),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_992),
.B(n_713),
.Y(n_1055)
);

AO21x2_ASAP7_75t_L g1056 ( 
.A1(n_864),
.A2(n_786),
.B(n_793),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_857),
.B(n_713),
.Y(n_1057)
);

OAI21xp33_ASAP7_75t_SL g1058 ( 
.A1(n_864),
.A2(n_801),
.B(n_799),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_961),
.A2(n_730),
.B(n_812),
.C(n_772),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_880),
.Y(n_1060)
);

INVx5_ASAP7_75t_L g1061 ( 
.A(n_973),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_995),
.A2(n_578),
.B(n_650),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_911),
.A2(n_782),
.B1(n_650),
.B2(n_578),
.Y(n_1063)
);

OAI21xp33_ASAP7_75t_L g1064 ( 
.A1(n_941),
.A2(n_650),
.B(n_9),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_901),
.B(n_578),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_1008),
.A2(n_578),
.B(n_661),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_931),
.B(n_598),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_1008),
.A2(n_578),
.B(n_661),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_994),
.Y(n_1069)
);

O2A1O1Ixp5_ASAP7_75t_L g1070 ( 
.A1(n_938),
.A2(n_598),
.B(n_69),
.C(n_134),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_969),
.A2(n_578),
.B1(n_667),
.B2(n_661),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_964),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_863),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_858),
.B(n_7),
.Y(n_1074)
);

AO32x1_ASAP7_75t_L g1075 ( 
.A1(n_940),
.A2(n_598),
.A3(n_12),
.B1(n_13),
.B2(n_32),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_890),
.B(n_11),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_865),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1011),
.A2(n_667),
.B(n_661),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_905),
.B(n_75),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_876),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_964),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_905),
.B(n_84),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_1011),
.A2(n_667),
.B(n_661),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_1014),
.B(n_13),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_878),
.Y(n_1085)
);

BUFx8_ASAP7_75t_L g1086 ( 
.A(n_873),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1007),
.B(n_598),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_897),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_942),
.A2(n_667),
.B(n_661),
.C(n_37),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_934),
.A2(n_598),
.B1(n_36),
.B2(n_38),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_915),
.A2(n_598),
.B(n_99),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_915),
.A2(n_98),
.B(n_176),
.Y(n_1092)
);

OAI22x1_ASAP7_75t_L g1093 ( 
.A1(n_902),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_916),
.Y(n_1094)
);

NAND2x1p5_ASAP7_75t_L g1095 ( 
.A(n_939),
.B(n_103),
.Y(n_1095)
);

NAND2x1p5_ASAP7_75t_L g1096 ( 
.A(n_947),
.B(n_902),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_854),
.Y(n_1097)
);

NAND3xp33_ASAP7_75t_SL g1098 ( 
.A(n_866),
.B(n_45),
.C(n_47),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_902),
.B(n_110),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_908),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_894),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_915),
.A2(n_114),
.B(n_172),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_991),
.B(n_912),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_975),
.B(n_45),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_908),
.Y(n_1105)
);

OR2x6_ASAP7_75t_SL g1106 ( 
.A(n_885),
.B(n_48),
.Y(n_1106)
);

NOR2xp67_ASAP7_75t_SL g1107 ( 
.A(n_955),
.B(n_48),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_926),
.A2(n_117),
.B(n_159),
.Y(n_1108)
);

NOR2xp67_ASAP7_75t_L g1109 ( 
.A(n_937),
.B(n_67),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_874),
.B(n_868),
.Y(n_1110)
);

NAND3xp33_ASAP7_75t_SL g1111 ( 
.A(n_971),
.B(n_49),
.C(n_52),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_917),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_925),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_886),
.A2(n_64),
.B1(n_157),
.B2(n_151),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_868),
.B(n_49),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_883),
.B(n_140),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_908),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_891),
.B(n_52),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_891),
.B(n_53),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_966),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_924),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1004),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1010),
.A2(n_54),
.B(n_55),
.C(n_135),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_927),
.A2(n_137),
.B(n_182),
.C(n_1026),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_925),
.B(n_855),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_867),
.B(n_936),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_974),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_940),
.A2(n_1028),
.B(n_957),
.C(n_1005),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_957),
.A2(n_898),
.B(n_893),
.C(n_899),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_909),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_913),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_867),
.B(n_929),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_969),
.A2(n_972),
.B1(n_981),
.B2(n_983),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_855),
.B(n_860),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_860),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_989),
.A2(n_972),
.B1(n_999),
.B2(n_896),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_928),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_979),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_893),
.A2(n_952),
.B(n_946),
.C(n_910),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_881),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_861),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_932),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_877),
.B(n_997),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_944),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_954),
.A2(n_875),
.B1(n_910),
.B2(n_952),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_887),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_977),
.B(n_968),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1009),
.A2(n_977),
.B(n_899),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1006),
.Y(n_1149)
);

O2A1O1Ixp5_ASAP7_75t_L g1150 ( 
.A1(n_984),
.A2(n_906),
.B(n_907),
.C(n_930),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1013),
.A2(n_1021),
.B(n_1024),
.C(n_958),
.Y(n_1151)
);

OR2x6_ASAP7_75t_L g1152 ( 
.A(n_881),
.B(n_887),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1029),
.A2(n_997),
.B(n_998),
.C(n_967),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_945),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_948),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1002),
.A2(n_1001),
.B(n_900),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_946),
.A2(n_1023),
.B1(n_1019),
.B2(n_976),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_990),
.A2(n_1016),
.B(n_1001),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_859),
.B(n_870),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1023),
.A2(n_1027),
.B(n_943),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_988),
.A2(n_949),
.B(n_1017),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_SL g1162 ( 
.A1(n_861),
.A2(n_892),
.B(n_919),
.C(n_933),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_950),
.Y(n_1163)
);

INVx5_ASAP7_75t_L g1164 ( 
.A(n_973),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_951),
.A2(n_963),
.B(n_985),
.C(n_987),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_903),
.A2(n_959),
.B(n_1022),
.Y(n_1166)
);

INVx5_ASAP7_75t_L g1167 ( 
.A(n_973),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_889),
.B(n_922),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_892),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_968),
.B(n_978),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_956),
.A2(n_965),
.B(n_962),
.C(n_960),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_881),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_986),
.A2(n_978),
.B1(n_882),
.B2(n_1031),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_904),
.A2(n_933),
.B(n_919),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_877),
.B(n_982),
.Y(n_1175)
);

OAI21xp33_ASAP7_75t_L g1176 ( 
.A1(n_993),
.A2(n_887),
.B(n_884),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_877),
.B(n_1031),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1012),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_973),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_877),
.B(n_1018),
.Y(n_1180)
);

BUFx12f_ASAP7_75t_L g1181 ( 
.A(n_1032),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_877),
.B(n_1030),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_1038),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_1042),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1148),
.A2(n_869),
.B(n_871),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1126),
.B(n_1020),
.Y(n_1186)
);

BUFx2_ASAP7_75t_SL g1187 ( 
.A(n_1052),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1132),
.A2(n_1000),
.B1(n_921),
.B2(n_920),
.Y(n_1188)
);

NAND3xp33_ASAP7_75t_L g1189 ( 
.A(n_1168),
.B(n_1025),
.C(n_1159),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1064),
.A2(n_1025),
.B(n_1033),
.C(n_1176),
.Y(n_1190)
);

BUFx4_ASAP7_75t_SL g1191 ( 
.A(n_1073),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1161),
.A2(n_1025),
.B(n_1156),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1045),
.B(n_1025),
.Y(n_1193)
);

NAND3xp33_ASAP7_75t_L g1194 ( 
.A(n_1084),
.B(n_1122),
.C(n_1107),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1069),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1038),
.Y(n_1196)
);

AO21x2_ASAP7_75t_L g1197 ( 
.A1(n_1151),
.A2(n_1148),
.B(n_1160),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1066),
.A2(n_1078),
.B(n_1068),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1139),
.B(n_1110),
.Y(n_1199)
);

AO21x2_ASAP7_75t_L g1200 ( 
.A1(n_1153),
.A2(n_1049),
.B(n_1056),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1083),
.A2(n_1166),
.B(n_1150),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1044),
.A2(n_1053),
.B(n_1059),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1147),
.B(n_1136),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1134),
.B(n_1125),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1175),
.A2(n_1129),
.B(n_1145),
.Y(n_1205)
);

AOI211x1_ASAP7_75t_L g1206 ( 
.A1(n_1098),
.A2(n_1111),
.B(n_1064),
.C(n_1104),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1039),
.A2(n_1174),
.B(n_1165),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1145),
.A2(n_1157),
.B(n_1176),
.Y(n_1208)
);

INVxp67_ASAP7_75t_SL g1209 ( 
.A(n_1180),
.Y(n_1209)
);

AOI21xp33_ASAP7_75t_L g1210 ( 
.A1(n_1058),
.A2(n_1128),
.B(n_1123),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1074),
.B(n_1076),
.Y(n_1211)
);

OA21x2_ASAP7_75t_L g1212 ( 
.A1(n_1034),
.A2(n_1089),
.B(n_1157),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1171),
.A2(n_1182),
.B(n_1177),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1046),
.B(n_1040),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1058),
.A2(n_1133),
.B(n_1109),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1037),
.B(n_1057),
.Y(n_1216)
);

O2A1O1Ixp5_ASAP7_75t_SL g1217 ( 
.A1(n_1114),
.A2(n_1119),
.B(n_1115),
.C(n_1118),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1043),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1055),
.B(n_1077),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1133),
.A2(n_1109),
.B(n_1173),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_1038),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1080),
.B(n_1085),
.Y(n_1222)
);

INVx4_ASAP7_75t_L g1223 ( 
.A(n_1061),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1061),
.A2(n_1167),
.B(n_1164),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1130),
.Y(n_1225)
);

INVx6_ASAP7_75t_L g1226 ( 
.A(n_1086),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1061),
.A2(n_1164),
.B1(n_1167),
.B2(n_1090),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1164),
.A2(n_1167),
.B(n_1143),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1134),
.B(n_1131),
.Y(n_1229)
);

INVx3_ASAP7_75t_SL g1230 ( 
.A(n_1152),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1071),
.A2(n_1062),
.B(n_1173),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1113),
.A2(n_1146),
.B(n_1124),
.C(n_1099),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_1131),
.B(n_1125),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1088),
.B(n_1163),
.Y(n_1234)
);

INVxp67_ASAP7_75t_SL g1235 ( 
.A(n_1179),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1067),
.A2(n_1056),
.B(n_1054),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1071),
.A2(n_1170),
.B(n_1178),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1094),
.B(n_1121),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1116),
.A2(n_1070),
.B(n_1142),
.C(n_1144),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1137),
.B(n_1155),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1154),
.Y(n_1241)
);

AO21x2_ASAP7_75t_L g1242 ( 
.A1(n_1162),
.A2(n_1087),
.B(n_1063),
.Y(n_1242)
);

NAND3xp33_ASAP7_75t_L g1243 ( 
.A(n_1050),
.B(n_1152),
.C(n_1082),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1065),
.A2(n_1050),
.B(n_1179),
.Y(n_1244)
);

AO22x2_ASAP7_75t_L g1245 ( 
.A1(n_1075),
.A2(n_1172),
.B1(n_1116),
.B2(n_1093),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1036),
.B(n_1112),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1041),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1092),
.A2(n_1102),
.B(n_1108),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1047),
.A2(n_1138),
.B(n_1048),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1060),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1135),
.B(n_1082),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1072),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1120),
.A2(n_1127),
.A3(n_1091),
.B(n_1075),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1035),
.B(n_1051),
.Y(n_1254)
);

AO21x2_ASAP7_75t_L g1255 ( 
.A1(n_1079),
.A2(n_1075),
.B(n_1179),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1035),
.B(n_1051),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1072),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1079),
.A2(n_1097),
.B(n_1095),
.Y(n_1258)
);

NAND3xp33_ASAP7_75t_SL g1259 ( 
.A(n_1140),
.B(n_1096),
.C(n_1181),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1141),
.B(n_1169),
.Y(n_1260)
);

AND3x4_ASAP7_75t_L g1261 ( 
.A(n_1106),
.B(n_1086),
.C(n_1101),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1072),
.A2(n_1081),
.B(n_1100),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1100),
.B(n_1105),
.Y(n_1263)
);

AOI21x1_ASAP7_75t_SL g1264 ( 
.A1(n_1105),
.A2(n_1117),
.B(n_1104),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1105),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1117),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1117),
.A2(n_872),
.B(n_1044),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_1042),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1168),
.A2(n_935),
.B1(n_707),
.B2(n_690),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1168),
.A2(n_872),
.B(n_970),
.C(n_677),
.Y(n_1270)
);

AO21x1_ASAP7_75t_L g1271 ( 
.A1(n_1136),
.A2(n_879),
.B(n_1157),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_SL g1272 ( 
.A1(n_1151),
.A2(n_1136),
.B(n_1153),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1126),
.B(n_1132),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1158),
.A2(n_1009),
.B(n_1161),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1046),
.Y(n_1275)
);

AOI21xp33_ASAP7_75t_L g1276 ( 
.A1(n_1064),
.A2(n_872),
.B(n_707),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1045),
.B(n_888),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1158),
.A2(n_1009),
.B(n_1161),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1148),
.A2(n_1049),
.B(n_864),
.Y(n_1279)
);

O2A1O1Ixp5_ASAP7_75t_L g1280 ( 
.A1(n_1168),
.A2(n_707),
.B(n_743),
.C(n_914),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1148),
.A2(n_1049),
.B(n_864),
.Y(n_1281)
);

INVxp67_ASAP7_75t_L g1282 ( 
.A(n_1103),
.Y(n_1282)
);

O2A1O1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1098),
.A2(n_707),
.B(n_677),
.C(n_728),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1126),
.B(n_1132),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1158),
.A2(n_1009),
.B(n_1161),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1158),
.A2(n_1009),
.B(n_1161),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1158),
.A2(n_1009),
.B(n_1161),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1126),
.B(n_1132),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1044),
.A2(n_872),
.B(n_1053),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1044),
.A2(n_872),
.B(n_1053),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1046),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1126),
.B(n_1132),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1045),
.B(n_888),
.Y(n_1293)
);

NOR2xp67_ASAP7_75t_SL g1294 ( 
.A(n_1061),
.B(n_1164),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1151),
.A2(n_1157),
.A3(n_1071),
.B(n_1136),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1038),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1148),
.A2(n_1049),
.B(n_864),
.Y(n_1297)
);

NAND3x1_ASAP7_75t_L g1298 ( 
.A(n_1159),
.B(n_824),
.C(n_683),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1179),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1148),
.A2(n_1049),
.B(n_864),
.Y(n_1300)
);

BUFx4f_ASAP7_75t_L g1301 ( 
.A(n_1038),
.Y(n_1301)
);

INVx5_ASAP7_75t_L g1302 ( 
.A(n_1179),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1069),
.Y(n_1303)
);

NAND3xp33_ASAP7_75t_L g1304 ( 
.A(n_1168),
.B(n_707),
.C(n_872),
.Y(n_1304)
);

INVx4_ASAP7_75t_L g1305 ( 
.A(n_1061),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_1042),
.Y(n_1306)
);

AOI31xp67_ASAP7_75t_L g1307 ( 
.A1(n_1049),
.A2(n_864),
.A3(n_984),
.B(n_886),
.Y(n_1307)
);

NOR2xp67_ASAP7_75t_L g1308 ( 
.A(n_1042),
.B(n_857),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1044),
.A2(n_872),
.B(n_1053),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1045),
.B(n_888),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1126),
.B(n_1132),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1103),
.B(n_923),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1148),
.A2(n_1049),
.B(n_864),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1126),
.B(n_1132),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1148),
.A2(n_1049),
.B(n_864),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1149),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1126),
.B(n_1132),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1134),
.B(n_1125),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1044),
.A2(n_872),
.B(n_1053),
.Y(n_1319)
);

CKINVDCx14_ASAP7_75t_R g1320 ( 
.A(n_1042),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1148),
.A2(n_1049),
.B(n_864),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1042),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1038),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1126),
.B(n_1132),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1148),
.A2(n_1049),
.B(n_864),
.Y(n_1325)
);

AOI211x1_ASAP7_75t_L g1326 ( 
.A1(n_1098),
.A2(n_830),
.B(n_1015),
.C(n_1111),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1126),
.B(n_1132),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1044),
.A2(n_872),
.B(n_1053),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1168),
.A2(n_872),
.B(n_970),
.C(n_677),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1046),
.B(n_888),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1045),
.B(n_888),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1249),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1192),
.A2(n_1278),
.B(n_1274),
.Y(n_1333)
);

OAI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1269),
.A2(n_1304),
.B1(n_1194),
.B2(n_1243),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1301),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1285),
.A2(n_1287),
.B(n_1286),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1195),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1303),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1301),
.Y(n_1339)
);

O2A1O1Ixp5_ASAP7_75t_L g1340 ( 
.A1(n_1280),
.A2(n_1276),
.B(n_1309),
.C(n_1289),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1198),
.A2(n_1201),
.B(n_1207),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1222),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1270),
.B(n_1329),
.Y(n_1343)
);

A2O1A1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1276),
.A2(n_1328),
.B(n_1309),
.C(n_1319),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1298),
.A2(n_1282),
.B1(n_1209),
.B2(n_1189),
.Y(n_1345)
);

AO21x2_ASAP7_75t_L g1346 ( 
.A1(n_1210),
.A2(n_1202),
.B(n_1289),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1271),
.A2(n_1319),
.B1(n_1328),
.B2(n_1290),
.Y(n_1347)
);

AO21x2_ASAP7_75t_L g1348 ( 
.A1(n_1210),
.A2(n_1202),
.B(n_1290),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1330),
.Y(n_1349)
);

AO21x2_ASAP7_75t_L g1350 ( 
.A1(n_1185),
.A2(n_1215),
.B(n_1220),
.Y(n_1350)
);

AO21x2_ASAP7_75t_L g1351 ( 
.A1(n_1215),
.A2(n_1220),
.B(n_1205),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1268),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1283),
.A2(n_1217),
.B(n_1199),
.Y(n_1353)
);

BUFx12f_ASAP7_75t_L g1354 ( 
.A(n_1225),
.Y(n_1354)
);

NAND2x1p5_ASAP7_75t_L g1355 ( 
.A(n_1294),
.B(n_1223),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1204),
.B(n_1318),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1277),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1234),
.Y(n_1358)
);

AO21x2_ASAP7_75t_L g1359 ( 
.A1(n_1199),
.A2(n_1281),
.B(n_1279),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1297),
.A2(n_1300),
.B(n_1313),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1234),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1238),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1312),
.A2(n_1317),
.B1(n_1311),
.B2(n_1292),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1211),
.B(n_1293),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1248),
.A2(n_1237),
.B(n_1231),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1275),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1315),
.A2(n_1325),
.B(n_1321),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_1306),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1310),
.A2(n_1331),
.B1(n_1308),
.B2(n_1251),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1236),
.A2(n_1213),
.B(n_1264),
.Y(n_1370)
);

OA21x2_ASAP7_75t_L g1371 ( 
.A1(n_1208),
.A2(n_1190),
.B(n_1267),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1273),
.A2(n_1327),
.B1(n_1311),
.B2(n_1314),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1191),
.Y(n_1373)
);

NAND2x1p5_ASAP7_75t_L g1374 ( 
.A(n_1223),
.B(n_1305),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1212),
.A2(n_1197),
.B1(n_1245),
.B2(n_1203),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1203),
.A2(n_1244),
.B(n_1239),
.Y(n_1376)
);

OAI22x1_ASAP7_75t_L g1377 ( 
.A1(n_1261),
.A2(n_1230),
.B1(n_1212),
.B2(n_1233),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1291),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1188),
.A2(n_1228),
.B(n_1224),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1284),
.A2(n_1327),
.B(n_1324),
.Y(n_1380)
);

OR2x6_ASAP7_75t_L g1381 ( 
.A(n_1258),
.B(n_1232),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1284),
.A2(n_1292),
.B(n_1288),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1204),
.B(n_1318),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1288),
.B(n_1324),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1263),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1229),
.B(n_1299),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1219),
.A2(n_1227),
.B(n_1216),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1302),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1241),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1238),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1314),
.B(n_1317),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_1320),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1302),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1200),
.A2(n_1197),
.B(n_1227),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1219),
.A2(n_1216),
.B(n_1240),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1186),
.A2(n_1307),
.B(n_1214),
.Y(n_1396)
);

AO31x2_ASAP7_75t_L g1397 ( 
.A1(n_1200),
.A2(n_1186),
.A3(n_1240),
.B(n_1295),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1218),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1193),
.A2(n_1246),
.B(n_1316),
.Y(n_1399)
);

AOI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1326),
.A2(n_1206),
.B1(n_1245),
.B2(n_1259),
.C(n_1187),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1246),
.A2(n_1247),
.B(n_1250),
.Y(n_1401)
);

NAND2x1p5_ASAP7_75t_L g1402 ( 
.A(n_1305),
.B(n_1302),
.Y(n_1402)
);

BUFx12f_ASAP7_75t_L g1403 ( 
.A(n_1226),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_L g1404 ( 
.A(n_1184),
.B(n_1322),
.C(n_1256),
.Y(n_1404)
);

NOR3xp33_ASAP7_75t_L g1405 ( 
.A(n_1235),
.B(n_1260),
.C(n_1256),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1226),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1262),
.A2(n_1254),
.B(n_1260),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1254),
.A2(n_1266),
.B(n_1265),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1183),
.Y(n_1409)
);

BUFx2_ASAP7_75t_R g1410 ( 
.A(n_1255),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1183),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1242),
.A2(n_1295),
.B(n_1253),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1295),
.A2(n_1253),
.B(n_1221),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1196),
.A2(n_1252),
.B(n_1257),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1252),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1252),
.A2(n_1323),
.B1(n_1257),
.B2(n_1296),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1296),
.A2(n_1270),
.B(n_1329),
.C(n_1276),
.Y(n_1417)
);

A2O1A1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1270),
.A2(n_1329),
.B(n_1276),
.C(n_872),
.Y(n_1418)
);

NOR2xp67_ASAP7_75t_L g1419 ( 
.A(n_1225),
.B(n_1042),
.Y(n_1419)
);

NOR2xp67_ASAP7_75t_L g1420 ( 
.A(n_1225),
.B(n_1042),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1280),
.A2(n_707),
.B(n_1304),
.Y(n_1421)
);

INVx2_ASAP7_75t_SL g1422 ( 
.A(n_1191),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1279),
.A2(n_1049),
.B(n_1281),
.Y(n_1423)
);

NOR2x1_ASAP7_75t_R g1424 ( 
.A(n_1226),
.B(n_885),
.Y(n_1424)
);

AO21x2_ASAP7_75t_L g1425 ( 
.A1(n_1210),
.A2(n_1276),
.B(n_1202),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1211),
.B(n_1277),
.Y(n_1426)
);

NAND3xp33_ASAP7_75t_L g1427 ( 
.A(n_1270),
.B(n_707),
.C(n_1329),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1330),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1304),
.B(n_1270),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1218),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1191),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1192),
.A2(n_1278),
.B(n_1274),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1301),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1268),
.Y(n_1434)
);

AOI221xp5_ASAP7_75t_L g1435 ( 
.A1(n_1276),
.A2(n_677),
.B1(n_707),
.B2(n_1283),
.C(n_824),
.Y(n_1435)
);

BUFx12f_ASAP7_75t_L g1436 ( 
.A(n_1225),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1301),
.Y(n_1437)
);

AO21x2_ASAP7_75t_L g1438 ( 
.A1(n_1210),
.A2(n_1276),
.B(n_1202),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1304),
.A2(n_872),
.B1(n_1276),
.B2(n_1098),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1218),
.Y(n_1440)
);

OR2x6_ASAP7_75t_L g1441 ( 
.A(n_1272),
.B(n_1243),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1223),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1270),
.B(n_1329),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1280),
.A2(n_707),
.B(n_1304),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1195),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1195),
.Y(n_1446)
);

AO21x2_ASAP7_75t_L g1447 ( 
.A1(n_1210),
.A2(n_1276),
.B(n_1202),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1218),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1195),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1304),
.A2(n_872),
.B1(n_1276),
.B2(n_1098),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1211),
.B(n_1277),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1211),
.B(n_1277),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1195),
.Y(n_1453)
);

AOI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1199),
.A2(n_1205),
.B(n_1185),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1192),
.A2(n_1278),
.B(n_1274),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1360),
.A2(n_1367),
.B(n_1423),
.Y(n_1456)
);

O2A1O1Ixp5_ASAP7_75t_L g1457 ( 
.A1(n_1429),
.A2(n_1343),
.B(n_1443),
.C(n_1421),
.Y(n_1457)
);

OA22x2_ASAP7_75t_L g1458 ( 
.A1(n_1369),
.A2(n_1377),
.B1(n_1429),
.B2(n_1363),
.Y(n_1458)
);

OA21x2_ASAP7_75t_L g1459 ( 
.A1(n_1394),
.A2(n_1353),
.B(n_1412),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1364),
.B(n_1426),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1349),
.B(n_1428),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1357),
.B(n_1451),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1398),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1452),
.B(n_1366),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1372),
.B(n_1380),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1389),
.Y(n_1466)
);

OA21x2_ASAP7_75t_L g1467 ( 
.A1(n_1340),
.A2(n_1365),
.B(n_1444),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1337),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1347),
.A2(n_1443),
.B1(n_1343),
.B2(n_1439),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1352),
.Y(n_1470)
);

O2A1O1Ixp5_ASAP7_75t_L g1471 ( 
.A1(n_1418),
.A2(n_1427),
.B(n_1344),
.C(n_1334),
.Y(n_1471)
);

OA22x2_ASAP7_75t_L g1472 ( 
.A1(n_1441),
.A2(n_1345),
.B1(n_1382),
.B2(n_1391),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1350),
.A2(n_1351),
.B(n_1359),
.Y(n_1473)
);

O2A1O1Ixp5_ASAP7_75t_L g1474 ( 
.A1(n_1418),
.A2(n_1344),
.B(n_1334),
.C(n_1454),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1338),
.Y(n_1475)
);

NOR2xp67_ASAP7_75t_L g1476 ( 
.A(n_1404),
.B(n_1419),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1356),
.B(n_1383),
.Y(n_1477)
);

O2A1O1Ixp5_ASAP7_75t_L g1478 ( 
.A1(n_1417),
.A2(n_1396),
.B(n_1384),
.C(n_1399),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_SL g1479 ( 
.A1(n_1435),
.A2(n_1417),
.B(n_1393),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1384),
.B(n_1395),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1347),
.A2(n_1439),
.B1(n_1450),
.B2(n_1410),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1415),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1378),
.B(n_1441),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1395),
.B(n_1342),
.Y(n_1484)
);

NOR2x1_ASAP7_75t_L g1485 ( 
.A(n_1381),
.B(n_1420),
.Y(n_1485)
);

O2A1O1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1450),
.A2(n_1441),
.B(n_1381),
.C(n_1400),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1352),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1371),
.A2(n_1358),
.B1(n_1361),
.B2(n_1390),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1411),
.B(n_1405),
.Y(n_1489)
);

OA21x2_ASAP7_75t_L g1490 ( 
.A1(n_1365),
.A2(n_1370),
.B(n_1341),
.Y(n_1490)
);

NOR3xp33_ASAP7_75t_L g1491 ( 
.A(n_1424),
.B(n_1379),
.C(n_1387),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1370),
.A2(n_1341),
.B(n_1379),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1346),
.A2(n_1348),
.B(n_1376),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_SL g1494 ( 
.A1(n_1388),
.A2(n_1393),
.B(n_1376),
.Y(n_1494)
);

O2A1O1Ixp33_ASAP7_75t_L g1495 ( 
.A1(n_1425),
.A2(n_1438),
.B(n_1447),
.C(n_1362),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1408),
.Y(n_1496)
);

AOI21x1_ASAP7_75t_SL g1497 ( 
.A1(n_1447),
.A2(n_1376),
.B(n_1375),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1388),
.A2(n_1393),
.B(n_1355),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_SL g1499 ( 
.A1(n_1388),
.A2(n_1393),
.B(n_1355),
.Y(n_1499)
);

O2A1O1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1445),
.A2(n_1453),
.B(n_1449),
.C(n_1446),
.Y(n_1500)
);

O2A1O1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1371),
.A2(n_1401),
.B(n_1375),
.C(n_1406),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1398),
.A2(n_1448),
.B1(n_1440),
.B2(n_1430),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1409),
.B(n_1416),
.Y(n_1503)
);

AND2x6_ASAP7_75t_L g1504 ( 
.A(n_1388),
.B(n_1442),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1333),
.A2(n_1455),
.B(n_1432),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1397),
.B(n_1413),
.Y(n_1506)
);

NOR2x1_ASAP7_75t_SL g1507 ( 
.A(n_1413),
.B(n_1332),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1414),
.B(n_1448),
.Y(n_1508)
);

AOI21x1_ASAP7_75t_SL g1509 ( 
.A1(n_1392),
.A2(n_1403),
.B(n_1436),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1397),
.B(n_1407),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1440),
.B(n_1442),
.Y(n_1511)
);

OAI31xp33_ASAP7_75t_L g1512 ( 
.A1(n_1422),
.A2(n_1431),
.A3(n_1374),
.B(n_1402),
.Y(n_1512)
);

OA21x2_ASAP7_75t_L g1513 ( 
.A1(n_1333),
.A2(n_1455),
.B(n_1432),
.Y(n_1513)
);

INVxp67_ASAP7_75t_L g1514 ( 
.A(n_1434),
.Y(n_1514)
);

INVx3_ASAP7_75t_SL g1515 ( 
.A(n_1373),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1397),
.B(n_1407),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_SL g1517 ( 
.A1(n_1402),
.A2(n_1335),
.B(n_1437),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1415),
.A2(n_1433),
.B1(n_1339),
.B2(n_1437),
.Y(n_1518)
);

O2A1O1Ixp33_ASAP7_75t_L g1519 ( 
.A1(n_1368),
.A2(n_1433),
.B(n_1339),
.C(n_1437),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1354),
.Y(n_1520)
);

BUFx12f_ASAP7_75t_L g1521 ( 
.A(n_1373),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1336),
.Y(n_1522)
);

O2A1O1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1368),
.A2(n_1354),
.B(n_1436),
.C(n_1434),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1394),
.A2(n_1353),
.B(n_1412),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1398),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1385),
.B(n_1386),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1372),
.B(n_1363),
.Y(n_1527)
);

NOR2xp67_ASAP7_75t_L g1528 ( 
.A(n_1404),
.B(n_1282),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1364),
.B(n_1426),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1347),
.A2(n_1270),
.B1(n_1329),
.B2(n_1298),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1366),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1372),
.B(n_1363),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1349),
.B(n_1428),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1364),
.B(n_1426),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1360),
.A2(n_1272),
.B(n_1367),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1347),
.A2(n_1270),
.B1(n_1329),
.B2(n_1298),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1364),
.B(n_1426),
.Y(n_1537)
);

O2A1O1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1334),
.A2(n_1270),
.B(n_1329),
.C(n_1283),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1484),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1484),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_R g1541 ( 
.A(n_1470),
.B(n_1487),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1459),
.B(n_1524),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1514),
.B(n_1462),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1480),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1460),
.B(n_1529),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1459),
.B(n_1524),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1516),
.B(n_1493),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1508),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1522),
.Y(n_1549)
);

OR2x6_ASAP7_75t_L g1550 ( 
.A(n_1535),
.B(n_1456),
.Y(n_1550)
);

INVxp67_ASAP7_75t_L g1551 ( 
.A(n_1496),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1510),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1510),
.B(n_1507),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1467),
.B(n_1473),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1483),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1491),
.B(n_1466),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1505),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1506),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1469),
.A2(n_1536),
.B1(n_1530),
.B2(n_1481),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1505),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1488),
.B(n_1461),
.Y(n_1561)
);

OAI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1538),
.A2(n_1471),
.B(n_1457),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1488),
.B(n_1533),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1513),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1474),
.A2(n_1478),
.B(n_1532),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1490),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1468),
.B(n_1475),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1538),
.A2(n_1536),
.B(n_1530),
.Y(n_1568)
);

OA21x2_ASAP7_75t_L g1569 ( 
.A1(n_1527),
.A2(n_1532),
.B(n_1465),
.Y(n_1569)
);

AOI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1485),
.A2(n_1469),
.B(n_1527),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1500),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1531),
.Y(n_1572)
);

OAI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1486),
.A2(n_1479),
.B(n_1481),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1495),
.B(n_1492),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1500),
.Y(n_1575)
);

OR2x6_ASAP7_75t_L g1576 ( 
.A(n_1494),
.B(n_1501),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1501),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1472),
.B(n_1458),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1489),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1472),
.B(n_1486),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1458),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1521),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1464),
.B(n_1526),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1503),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1569),
.B(n_1551),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1549),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1552),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1556),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1568),
.A2(n_1528),
.B1(n_1534),
.B2(n_1537),
.Y(n_1589)
);

NAND3xp33_ASAP7_75t_L g1590 ( 
.A(n_1568),
.B(n_1562),
.C(n_1559),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1552),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1569),
.B(n_1476),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1558),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1573),
.A2(n_1502),
.B1(n_1520),
.B2(n_1482),
.Y(n_1594)
);

INVx5_ASAP7_75t_L g1595 ( 
.A(n_1576),
.Y(n_1595)
);

INVx4_ASAP7_75t_L g1596 ( 
.A(n_1576),
.Y(n_1596)
);

AO22x1_ASAP7_75t_L g1597 ( 
.A1(n_1562),
.A2(n_1502),
.B1(n_1504),
.B2(n_1520),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1573),
.B(n_1519),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1557),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1569),
.B(n_1511),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1547),
.B(n_1497),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1547),
.B(n_1542),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1556),
.Y(n_1603)
);

CKINVDCx20_ASAP7_75t_R g1604 ( 
.A(n_1541),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1542),
.B(n_1477),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1561),
.B(n_1525),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1602),
.B(n_1548),
.Y(n_1607)
);

AOI21xp33_ASAP7_75t_SL g1608 ( 
.A1(n_1590),
.A2(n_1523),
.B(n_1580),
.Y(n_1608)
);

INVx6_ASAP7_75t_L g1609 ( 
.A(n_1595),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1586),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1586),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_SL g1612 ( 
.A1(n_1598),
.A2(n_1565),
.B(n_1580),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1588),
.B(n_1553),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1588),
.Y(n_1614)
);

NAND3xp33_ASAP7_75t_L g1615 ( 
.A(n_1590),
.B(n_1581),
.C(n_1578),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1605),
.B(n_1551),
.Y(n_1616)
);

OAI33xp33_ASAP7_75t_L g1617 ( 
.A1(n_1585),
.A2(n_1581),
.A3(n_1575),
.B1(n_1571),
.B2(n_1577),
.B3(n_1544),
.Y(n_1617)
);

BUFx3_ASAP7_75t_L g1618 ( 
.A(n_1604),
.Y(n_1618)
);

OAI221xp5_ASAP7_75t_SL g1619 ( 
.A1(n_1589),
.A2(n_1578),
.B1(n_1576),
.B2(n_1577),
.C(n_1512),
.Y(n_1619)
);

OAI211xp5_ASAP7_75t_SL g1620 ( 
.A1(n_1598),
.A2(n_1523),
.B(n_1561),
.C(n_1563),
.Y(n_1620)
);

NOR4xp25_ASAP7_75t_SL g1621 ( 
.A(n_1588),
.B(n_1579),
.C(n_1571),
.D(n_1575),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1586),
.Y(n_1622)
);

OAI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1594),
.A2(n_1570),
.B(n_1565),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1587),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1604),
.Y(n_1625)
);

OR2x6_ASAP7_75t_SL g1626 ( 
.A(n_1592),
.B(n_1583),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_SL g1627 ( 
.A1(n_1595),
.A2(n_1565),
.B1(n_1576),
.B2(n_1569),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1587),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1594),
.A2(n_1569),
.B1(n_1565),
.B2(n_1579),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1589),
.A2(n_1565),
.B1(n_1543),
.B2(n_1518),
.Y(n_1630)
);

NOR3xp33_ASAP7_75t_L g1631 ( 
.A(n_1597),
.B(n_1570),
.C(n_1518),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1591),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1605),
.B(n_1572),
.Y(n_1633)
);

OAI221xp5_ASAP7_75t_L g1634 ( 
.A1(n_1592),
.A2(n_1563),
.B1(n_1555),
.B2(n_1550),
.C(n_1572),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1602),
.B(n_1548),
.Y(n_1635)
);

AO21x2_ASAP7_75t_L g1636 ( 
.A1(n_1585),
.A2(n_1554),
.B(n_1566),
.Y(n_1636)
);

BUFx6f_ASAP7_75t_L g1637 ( 
.A(n_1595),
.Y(n_1637)
);

INVx4_ASAP7_75t_SL g1638 ( 
.A(n_1603),
.Y(n_1638)
);

AOI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1600),
.A2(n_1545),
.B1(n_1556),
.B2(n_1567),
.C(n_1584),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1605),
.B(n_1584),
.Y(n_1640)
);

AOI33xp33_ASAP7_75t_L g1641 ( 
.A1(n_1601),
.A2(n_1546),
.A3(n_1567),
.B1(n_1584),
.B2(n_1574),
.B3(n_1540),
.Y(n_1641)
);

AOI222xp33_ASAP7_75t_L g1642 ( 
.A1(n_1597),
.A2(n_1546),
.B1(n_1567),
.B2(n_1540),
.C1(n_1539),
.C2(n_1544),
.Y(n_1642)
);

OA21x2_ASAP7_75t_L g1643 ( 
.A1(n_1599),
.A2(n_1554),
.B(n_1566),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1624),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1628),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1637),
.Y(n_1646)
);

AO21x2_ASAP7_75t_L g1647 ( 
.A1(n_1612),
.A2(n_1554),
.B(n_1574),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1615),
.Y(n_1648)
);

OA21x2_ASAP7_75t_L g1649 ( 
.A1(n_1623),
.A2(n_1566),
.B(n_1560),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1638),
.Y(n_1650)
);

INVx4_ASAP7_75t_SL g1651 ( 
.A(n_1609),
.Y(n_1651)
);

OA21x2_ASAP7_75t_L g1652 ( 
.A1(n_1629),
.A2(n_1564),
.B(n_1560),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1643),
.Y(n_1653)
);

INVxp67_ASAP7_75t_L g1654 ( 
.A(n_1615),
.Y(n_1654)
);

INVx5_ASAP7_75t_L g1655 ( 
.A(n_1637),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1626),
.B(n_1603),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1632),
.Y(n_1657)
);

INVx4_ASAP7_75t_SL g1658 ( 
.A(n_1609),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1626),
.B(n_1603),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1614),
.B(n_1601),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1614),
.Y(n_1661)
);

OR2x6_ASAP7_75t_L g1662 ( 
.A(n_1612),
.B(n_1609),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1638),
.B(n_1601),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1610),
.Y(n_1664)
);

CKINVDCx8_ASAP7_75t_R g1665 ( 
.A(n_1638),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1610),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1636),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1611),
.Y(n_1668)
);

AND4x1_ASAP7_75t_L g1669 ( 
.A(n_1631),
.B(n_1517),
.C(n_1498),
.D(n_1499),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1611),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1622),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1638),
.Y(n_1672)
);

AND2x6_ASAP7_75t_SL g1673 ( 
.A(n_1608),
.B(n_1515),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1655),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1656),
.B(n_1613),
.Y(n_1675)
);

AOI211x1_ASAP7_75t_L g1676 ( 
.A1(n_1656),
.A2(n_1634),
.B(n_1633),
.C(n_1616),
.Y(n_1676)
);

NAND2xp33_ASAP7_75t_R g1677 ( 
.A(n_1650),
.B(n_1608),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1664),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1653),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1648),
.B(n_1641),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1664),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1648),
.B(n_1640),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1656),
.B(n_1613),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1666),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1654),
.B(n_1636),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1659),
.B(n_1613),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1659),
.B(n_1613),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1654),
.B(n_1639),
.Y(n_1688)
);

AOI31xp33_ASAP7_75t_L g1689 ( 
.A1(n_1673),
.A2(n_1627),
.A3(n_1630),
.B(n_1617),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1666),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1644),
.B(n_1600),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1659),
.B(n_1607),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1663),
.B(n_1651),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1653),
.Y(n_1694)
);

BUFx2_ASAP7_75t_SL g1695 ( 
.A(n_1665),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1663),
.B(n_1651),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1663),
.B(n_1607),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1644),
.B(n_1630),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1651),
.B(n_1635),
.Y(n_1699)
);

INVx1_ASAP7_75t_SL g1700 ( 
.A(n_1650),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1668),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1668),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1645),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1670),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1651),
.B(n_1635),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1650),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1645),
.B(n_1657),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1653),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1651),
.B(n_1658),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1672),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1670),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1671),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1671),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1673),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1661),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1657),
.B(n_1593),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1715),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1693),
.B(n_1651),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1682),
.B(n_1606),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1715),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1709),
.B(n_1658),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1678),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1688),
.B(n_1660),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1682),
.B(n_1606),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1678),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1680),
.B(n_1660),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1681),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1681),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1684),
.Y(n_1729)
);

NAND3xp33_ASAP7_75t_L g1730 ( 
.A(n_1677),
.B(n_1649),
.C(n_1620),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1684),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1690),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1690),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1703),
.B(n_1661),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1714),
.B(n_1665),
.Y(n_1735)
);

OAI22xp33_ASAP7_75t_SL g1736 ( 
.A1(n_1698),
.A2(n_1619),
.B1(n_1665),
.B2(n_1662),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1695),
.A2(n_1596),
.B1(n_1662),
.B2(n_1647),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1709),
.B(n_1658),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1693),
.B(n_1658),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1707),
.B(n_1606),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1696),
.B(n_1658),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1701),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1700),
.B(n_1660),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1695),
.B(n_1618),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1701),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1689),
.B(n_1618),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1676),
.B(n_1642),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1702),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1696),
.B(n_1658),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1691),
.B(n_1649),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1702),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1704),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1749),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1722),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1725),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1718),
.B(n_1699),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1739),
.B(n_1699),
.Y(n_1757)
);

INVx1_ASAP7_75t_SL g1758 ( 
.A(n_1735),
.Y(n_1758)
);

OAI21x1_ASAP7_75t_L g1759 ( 
.A1(n_1730),
.A2(n_1694),
.B(n_1679),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1750),
.Y(n_1760)
);

INVx1_ASAP7_75t_SL g1761 ( 
.A(n_1744),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1743),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1743),
.B(n_1700),
.Y(n_1763)
);

INVx4_ASAP7_75t_L g1764 ( 
.A(n_1721),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1746),
.A2(n_1662),
.B1(n_1596),
.B2(n_1705),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1736),
.A2(n_1689),
.B(n_1706),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1723),
.B(n_1706),
.Y(n_1767)
);

OAI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1747),
.A2(n_1662),
.B1(n_1655),
.B2(n_1672),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1741),
.B(n_1705),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1734),
.B(n_1710),
.Y(n_1770)
);

OA21x2_ASAP7_75t_L g1771 ( 
.A1(n_1730),
.A2(n_1694),
.B(n_1679),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1721),
.B(n_1692),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1727),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1738),
.B(n_1692),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1728),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_SL g1776 ( 
.A1(n_1736),
.A2(n_1649),
.B1(n_1652),
.B2(n_1710),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1729),
.Y(n_1777)
);

AOI22x1_ASAP7_75t_L g1778 ( 
.A1(n_1738),
.A2(n_1520),
.B1(n_1674),
.B2(n_1672),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1731),
.Y(n_1779)
);

AOI32xp33_ASAP7_75t_L g1780 ( 
.A1(n_1776),
.A2(n_1726),
.A3(n_1749),
.B1(n_1734),
.B2(n_1720),
.Y(n_1780)
);

CKINVDCx14_ASAP7_75t_R g1781 ( 
.A(n_1764),
.Y(n_1781)
);

AOI222xp33_ASAP7_75t_L g1782 ( 
.A1(n_1758),
.A2(n_1717),
.B1(n_1751),
.B2(n_1742),
.C1(n_1752),
.C2(n_1748),
.Y(n_1782)
);

AOI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1766),
.A2(n_1662),
.B1(n_1737),
.B2(n_1647),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1761),
.B(n_1676),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1777),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1766),
.B(n_1655),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1761),
.B(n_1625),
.Y(n_1787)
);

AOI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1776),
.A2(n_1745),
.B1(n_1732),
.B2(n_1733),
.C(n_1685),
.Y(n_1788)
);

OAI222xp33_ASAP7_75t_L g1789 ( 
.A1(n_1758),
.A2(n_1685),
.B1(n_1662),
.B2(n_1674),
.C1(n_1719),
.C2(n_1724),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1753),
.B(n_1697),
.Y(n_1790)
);

AOI322xp5_ASAP7_75t_L g1791 ( 
.A1(n_1767),
.A2(n_1762),
.A3(n_1768),
.B1(n_1774),
.B2(n_1772),
.C1(n_1753),
.C2(n_1757),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1756),
.B(n_1697),
.Y(n_1792)
);

INVxp33_ASAP7_75t_L g1793 ( 
.A(n_1756),
.Y(n_1793)
);

AOI31xp33_ASAP7_75t_L g1794 ( 
.A1(n_1753),
.A2(n_1582),
.A3(n_1740),
.B(n_1675),
.Y(n_1794)
);

AOI31xp33_ASAP7_75t_L g1795 ( 
.A1(n_1770),
.A2(n_1687),
.A3(n_1683),
.B(n_1686),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1772),
.B(n_1675),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_SL g1797 ( 
.A(n_1764),
.B(n_1655),
.Y(n_1797)
);

AOI221xp5_ASAP7_75t_L g1798 ( 
.A1(n_1767),
.A2(n_1667),
.B1(n_1647),
.B2(n_1653),
.C(n_1646),
.Y(n_1798)
);

NOR2x1_ASAP7_75t_L g1799 ( 
.A(n_1771),
.B(n_1625),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1777),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1787),
.B(n_1764),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1793),
.B(n_1764),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1790),
.B(n_1770),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1792),
.B(n_1757),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1781),
.B(n_1769),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1784),
.B(n_1769),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1786),
.A2(n_1771),
.B1(n_1759),
.B2(n_1762),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1799),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1785),
.B(n_1774),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1800),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1796),
.Y(n_1811)
);

NOR2x1_ASAP7_75t_L g1812 ( 
.A(n_1794),
.B(n_1771),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1791),
.B(n_1683),
.Y(n_1813)
);

AOI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1813),
.A2(n_1780),
.B1(n_1788),
.B2(n_1789),
.C(n_1798),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1807),
.A2(n_1783),
.B1(n_1795),
.B2(n_1765),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1805),
.B(n_1782),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1804),
.B(n_1763),
.Y(n_1817)
);

OAI31xp33_ASAP7_75t_SL g1818 ( 
.A1(n_1812),
.A2(n_1806),
.A3(n_1808),
.B(n_1759),
.Y(n_1818)
);

O2A1O1Ixp33_ASAP7_75t_L g1819 ( 
.A1(n_1808),
.A2(n_1789),
.B(n_1771),
.C(n_1797),
.Y(n_1819)
);

NAND3xp33_ASAP7_75t_L g1820 ( 
.A(n_1807),
.B(n_1771),
.C(n_1778),
.Y(n_1820)
);

AOI32xp33_ASAP7_75t_L g1821 ( 
.A1(n_1806),
.A2(n_1759),
.A3(n_1773),
.B1(n_1755),
.B2(n_1775),
.Y(n_1821)
);

OAI21xp33_ASAP7_75t_L g1822 ( 
.A1(n_1801),
.A2(n_1763),
.B(n_1755),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1809),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1809),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1802),
.B(n_1686),
.Y(n_1825)
);

XNOR2x1_ASAP7_75t_L g1826 ( 
.A(n_1816),
.B(n_1803),
.Y(n_1826)
);

OAI321xp33_ASAP7_75t_L g1827 ( 
.A1(n_1814),
.A2(n_1802),
.A3(n_1811),
.B1(n_1810),
.B2(n_1779),
.C(n_1754),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1817),
.Y(n_1828)
);

AOI21xp33_ASAP7_75t_L g1829 ( 
.A1(n_1818),
.A2(n_1819),
.B(n_1815),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1823),
.Y(n_1830)
);

OAI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1818),
.A2(n_1778),
.B1(n_1779),
.B2(n_1775),
.C(n_1773),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1830),
.B(n_1824),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1828),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1826),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1831),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1827),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1829),
.B(n_1825),
.Y(n_1837)
);

XNOR2x1_ASAP7_75t_L g1838 ( 
.A(n_1826),
.B(n_1820),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1834),
.B(n_1822),
.Y(n_1839)
);

OAI31xp33_ASAP7_75t_SL g1840 ( 
.A1(n_1838),
.A2(n_1821),
.A3(n_1777),
.B(n_1754),
.Y(n_1840)
);

NOR2x1_ASAP7_75t_L g1841 ( 
.A(n_1837),
.B(n_1832),
.Y(n_1841)
);

NOR2x1p5_ASAP7_75t_L g1842 ( 
.A(n_1832),
.B(n_1760),
.Y(n_1842)
);

XNOR2xp5_ASAP7_75t_L g1843 ( 
.A(n_1836),
.B(n_1835),
.Y(n_1843)
);

NAND2xp33_ASAP7_75t_R g1844 ( 
.A(n_1833),
.B(n_1621),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1840),
.B(n_1760),
.Y(n_1845)
);

AND3x2_ASAP7_75t_L g1846 ( 
.A(n_1839),
.B(n_1509),
.C(n_1760),
.Y(n_1846)
);

NOR3xp33_ASAP7_75t_L g1847 ( 
.A(n_1841),
.B(n_1463),
.C(n_1687),
.Y(n_1847)
);

OAI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1845),
.A2(n_1843),
.B1(n_1842),
.B2(n_1655),
.Y(n_1848)
);

AOI322xp5_ASAP7_75t_L g1849 ( 
.A1(n_1848),
.A2(n_1847),
.A3(n_1846),
.B1(n_1844),
.B2(n_1667),
.C1(n_1679),
.C2(n_1708),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_SL g1850 ( 
.A1(n_1849),
.A2(n_1662),
.B1(n_1655),
.B2(n_1646),
.Y(n_1850)
);

AOI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1849),
.A2(n_1646),
.B1(n_1655),
.B2(n_1708),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1850),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1851),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1853),
.A2(n_1708),
.B(n_1694),
.Y(n_1854)
);

OAI22x1_ASAP7_75t_L g1855 ( 
.A1(n_1852),
.A2(n_1655),
.B1(n_1669),
.B2(n_1713),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1854),
.A2(n_1711),
.B(n_1704),
.Y(n_1856)
);

INVxp33_ASAP7_75t_L g1857 ( 
.A(n_1856),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1857),
.B(n_1855),
.Y(n_1858)
);

OAI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1858),
.A2(n_1646),
.B1(n_1716),
.B2(n_1712),
.Y(n_1859)
);

OAI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1859),
.A2(n_1716),
.B1(n_1646),
.B2(n_1712),
.Y(n_1860)
);

AOI211xp5_ASAP7_75t_L g1861 ( 
.A1(n_1860),
.A2(n_1646),
.B(n_1713),
.C(n_1711),
.Y(n_1861)
);


endmodule