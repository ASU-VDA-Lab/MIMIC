module real_jpeg_21429_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_0),
.A2(n_10),
.B1(n_26),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_0),
.A2(n_5),
.B1(n_23),
.B2(n_28),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_1),
.A2(n_10),
.B1(n_26),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_1),
.A2(n_5),
.B1(n_23),
.B2(n_30),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_2),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_2),
.B(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_2),
.A2(n_3),
.B1(n_40),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_2),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_2),
.A2(n_40),
.B(n_59),
.C(n_105),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_3),
.A2(n_6),
.B1(n_38),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_3),
.A2(n_10),
.B1(n_26),
.B2(n_40),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_3),
.A2(n_5),
.B1(n_23),
.B2(n_40),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_SL g105 ( 
.A1(n_3),
.A2(n_6),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_3),
.B(n_120),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g129 ( 
.A1(n_3),
.A2(n_5),
.B(n_9),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_3),
.B(n_34),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_3),
.A2(n_7),
.B(n_38),
.C(n_151),
.Y(n_150)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_5),
.A2(n_9),
.B1(n_23),
.B2(n_24),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_5),
.B(n_48),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_7),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_6),
.A2(n_8),
.B1(n_38),
.B2(n_59),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_7),
.A2(n_10),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_9),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g25 ( 
.A1(n_9),
.A2(n_10),
.B1(n_24),
.B2(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_10),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_10),
.A2(n_24),
.B(n_40),
.C(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_89),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_88),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_76),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_15),
.B(n_76),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_65),
.B2(n_75),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_42),
.B2(n_43),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_31),
.B(n_41),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_31),
.Y(n_41)
);

OA22x2_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_27),
.B2(n_29),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_21),
.A2(n_22),
.B1(n_27),
.B2(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_21),
.B(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_22),
.B(n_40),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_23),
.B(n_141),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_26),
.A2(n_35),
.B(n_40),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_56),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_31),
.A2(n_32),
.B1(n_55),
.B2(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_31),
.B(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_31),
.A2(n_32),
.B1(n_70),
.B2(n_97),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_31),
.A2(n_97),
.B(n_153),
.C(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_31),
.A2(n_32),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_31),
.A2(n_56),
.B(n_73),
.C(n_102),
.Y(n_187)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_32),
.B(n_55),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_32),
.B(n_107),
.C(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_39),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_40),
.B(n_69),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_54),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_51),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_55),
.B1(n_56),
.B2(n_64),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_51),
.B1(n_64),
.B2(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_47),
.B(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_50),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_68),
.B1(n_69),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_51),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_71),
.Y(n_70)
);

AOI211xp5_ASAP7_75t_SL g95 ( 
.A1(n_55),
.A2(n_70),
.B(n_74),
.C(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_55),
.A2(n_56),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_72),
.B(n_73),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_67),
.A2(n_70),
.B1(n_97),
.B2(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_67),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_70),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_85),
.B1(n_97),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_70),
.A2(n_97),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_70),
.A2(n_97),
.B1(n_128),
.B2(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_70),
.B(n_107),
.C(n_132),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_70),
.A2(n_97),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_70),
.B(n_159),
.C(n_165),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_73),
.B(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_76),
.Y(n_192)
);

FAx1_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_81),
.CI(n_83),
.CON(n_76),
.SN(n_76)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_79),
.B1(n_102),
.B2(n_108),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_78),
.A2(n_79),
.B1(n_84),
.B2(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_84),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_190),
.B(n_193),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_121),
.B(n_176),
.C(n_189),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_109),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_92),
.B(n_109),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_101),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_94),
.B(n_99),
.C(n_101),
.Y(n_177)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_96),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_97),
.B(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_102),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_103),
.A2(n_104),
.B1(n_107),
.B2(n_116),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_107),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_116),
.B1(n_131),
.B2(n_134),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_107),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_107),
.B(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_107),
.A2(n_116),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_107),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_162)
);

NAND2x1_ASAP7_75t_SL g166 ( 
.A(n_107),
.B(n_150),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_117),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_110),
.A2(n_111),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_112),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_112),
.A2(n_113),
.B1(n_149),
.B2(n_153),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_114),
.A2(n_115),
.B1(n_117),
.B2(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_117),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_175),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_168),
.B(n_174),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_155),
.B(n_167),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_146),
.B(n_154),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_135),
.B(n_145),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_130),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_128),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_131),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_142),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_148),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_149),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_150),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_156),
.B(n_158),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_169),
.B(n_170),
.Y(n_174)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_177),
.B(n_178),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_187),
.B2(n_188),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_181),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_186),
.C(n_188),
.Y(n_191)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_183),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_187),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_191),
.B(n_192),
.Y(n_193)
);


endmodule