module fake_jpeg_2260_n_215 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_215);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_9),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_20),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_13),
.Y(n_75)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_81),
.B(n_82),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_85),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_68),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_SL g89 ( 
.A(n_83),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_75),
.B1(n_76),
.B2(n_74),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_90),
.A2(n_66),
.B1(n_1),
.B2(n_2),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_75),
.B1(n_69),
.B2(n_73),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_92),
.B1(n_67),
.B2(n_55),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_72),
.B1(n_58),
.B2(n_74),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_65),
.B1(n_76),
.B2(n_72),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_63),
.B1(n_77),
.B2(n_55),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_60),
.C(n_58),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_65),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_80),
.B(n_65),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_98),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_82),
.B1(n_78),
.B2(n_61),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_99),
.A2(n_105),
.B1(n_86),
.B2(n_3),
.Y(n_132)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_101),
.Y(n_135)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_117),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_95),
.B1(n_87),
.B2(n_88),
.Y(n_105)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_71),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_63),
.B1(n_55),
.B2(n_66),
.Y(n_109)
);

AO22x2_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_96),
.B1(n_86),
.B2(n_4),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_53),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_54),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_59),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_86),
.B1(n_96),
.B2(n_5),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_98),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_116),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_70),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_106),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_130),
.Y(n_147)
);

BUFx2_ASAP7_75t_SL g119 ( 
.A(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_0),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_109),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

NOR2x1_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_11),
.Y(n_151)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_133),
.B1(n_137),
.B2(n_12),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_103),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_105),
.B1(n_9),
.B2(n_10),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_86),
.B1(n_5),
.B2(n_6),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_136),
.B(n_8),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_86),
.B1(n_6),
.B2(n_7),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_2),
.B(n_8),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_139),
.B(n_125),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_133),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_141),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_149),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_145),
.A2(n_146),
.B1(n_156),
.B2(n_157),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_27),
.B1(n_50),
.B2(n_49),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_151),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_131),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_11),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_154),
.Y(n_173)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_128),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_25),
.B1(n_48),
.B2(n_47),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_23),
.B1(n_46),
.B2(n_43),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_158),
.A2(n_123),
.B(n_28),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_159),
.A2(n_146),
.B1(n_145),
.B2(n_157),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_12),
.B(n_13),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_123),
.B(n_15),
.Y(n_170)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

AND2x4_ASAP7_75t_SL g163 ( 
.A(n_140),
.B(n_123),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_166),
.A2(n_170),
.B(n_178),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_147),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_169),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_SL g172 ( 
.A1(n_155),
.A2(n_22),
.B(n_37),
.C(n_35),
.Y(n_172)
);

OA22x2_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_143),
.B1(n_160),
.B2(n_21),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_52),
.C(n_34),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_30),
.C(n_31),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_179),
.B1(n_156),
.B2(n_174),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_144),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_155),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_190),
.B1(n_179),
.B2(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_171),
.C(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_173),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_17),
.C(n_18),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_176),
.C(n_175),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_172),
.B1(n_191),
.B2(n_184),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_196),
.B(n_198),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_194),
.A2(n_199),
.B(n_182),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_172),
.C(n_163),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_163),
.Y(n_199)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_197),
.A2(n_185),
.B(n_184),
.Y(n_203)
);

OAI31xp33_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_204),
.A3(n_200),
.B(n_172),
.Y(n_205)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_199),
.Y(n_209)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_207),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_209),
.C(n_206),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_204),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_195),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_212),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_187),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_19),
.Y(n_215)
);


endmodule