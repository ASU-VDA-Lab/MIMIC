module fake_jpeg_20498_n_177 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_SL g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_32),
.Y(n_51)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_21),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_37),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_39),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_52),
.B1(n_41),
.B2(n_49),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_44),
.B(n_2),
.Y(n_73)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_42),
.B1(n_46),
.B2(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_14),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_30),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_25),
.B1(n_29),
.B2(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_69),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_55),
.B1(n_61),
.B2(n_65),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_32),
.B1(n_39),
.B2(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_29),
.B1(n_17),
.B2(n_18),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_63),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_60),
.B(n_8),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_20),
.B1(n_22),
.B2(n_19),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_20),
.C(n_22),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_68),
.Y(n_76)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_20),
.B1(n_16),
.B2(n_22),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_19),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_70),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_3),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_3),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_80),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_3),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_5),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_84),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_55),
.B1(n_63),
.B2(n_67),
.Y(n_99)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_7),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_62),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_83),
.B1(n_91),
.B2(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_96),
.B(n_11),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_63),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_106),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_101),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_81),
.B(n_62),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_66),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_104),
.B(n_78),
.Y(n_117)
);

CKINVDCx10_ASAP7_75t_R g101 ( 
.A(n_88),
.Y(n_101)
);

NOR2x1_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_67),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_65),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_109),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_65),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_114),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_77),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_82),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_123),
.C(n_100),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_86),
.B(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_121),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_87),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_79),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_86),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_124),
.Y(n_140)
);

AOI322xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_81),
.A3(n_89),
.B1(n_85),
.B2(n_88),
.C1(n_90),
.C2(n_11),
.Y(n_126)
);

OA21x2_ASAP7_75t_SL g134 ( 
.A1(n_126),
.A2(n_119),
.B(n_128),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_101),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_77),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_123),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_127),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_135),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_141),
.B1(n_124),
.B2(n_115),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_142),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_103),
.C(n_102),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_114),
.B1(n_84),
.B2(n_13),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_141),
.B1(n_125),
.B2(n_139),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_149),
.C(n_151),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

XNOR2x1_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_120),
.Y(n_151)
);

BUFx12_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_152),
.B(n_139),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_155),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_130),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_158),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_137),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_146),
.C(n_149),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_160),
.B(n_163),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_140),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_151),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_152),
.C(n_116),
.Y(n_169)
);

A2O1A1O1Ixp25_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_152),
.B(n_156),
.C(n_140),
.D(n_143),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_166),
.B(n_168),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_121),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_165),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_171),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_164),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_174),
.Y(n_177)
);


endmodule