module fake_jpeg_14151_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp33_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_9),
.B(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_21),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_46),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_69),
.Y(n_72)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_17),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_68),
.Y(n_75)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_56),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_43),
.B(n_59),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_76),
.B(n_81),
.Y(n_85)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_74),
.B(n_78),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_70),
.A2(n_43),
.B(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_45),
.B1(n_61),
.B2(n_51),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_23),
.B1(n_37),
.B2(n_34),
.Y(n_111)
);

OAI22x1_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_45),
.B1(n_57),
.B2(n_47),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_93),
.B1(n_102),
.B2(n_6),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_53),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_56),
.B1(n_2),
.B2(n_3),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_73),
.Y(n_107)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_98),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_1),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_73),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_100),
.Y(n_112)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_97),
.B(n_4),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_107),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_5),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_106),
.A2(n_108),
.B(n_109),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_22),
.C(n_39),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_5),
.Y(n_110)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_102),
.B1(n_10),
.B2(n_11),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_6),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_8),
.B1(n_12),
.B2(n_14),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_7),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_7),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_116),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_87),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_40),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_8),
.B(n_9),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_131),
.B(n_105),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_130),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_12),
.B1(n_16),
.B2(n_20),
.Y(n_131)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_104),
.A3(n_112),
.B1(n_106),
.B2(n_121),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_137),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_109),
.C(n_120),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_136),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_117),
.C(n_118),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_134),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_130),
.B1(n_127),
.B2(n_129),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_124),
.C(n_132),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_142),
.B(n_139),
.Y(n_144)
);

AOI322xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_122),
.A3(n_126),
.B1(n_139),
.B2(n_118),
.C1(n_33),
.C2(n_24),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_25),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_28),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_30),
.Y(n_148)
);


endmodule