module real_jpeg_25446_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_0),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_0),
.B(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_0),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_0),
.B(n_25),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_0),
.B(n_41),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_0),
.B(n_45),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_0),
.B(n_27),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_0),
.B(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_2),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_2),
.B(n_30),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_2),
.B(n_62),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_2),
.B(n_25),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_2),
.B(n_41),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_2),
.B(n_27),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_4),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_4),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_4),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_4),
.B(n_27),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_4),
.B(n_45),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_4),
.B(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g32 ( 
.A(n_6),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_7),
.B(n_27),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_7),
.B(n_45),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_7),
.B(n_16),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_9),
.Y(n_103)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_11),
.B(n_25),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_11),
.B(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_11),
.B(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_11),
.B(n_41),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_11),
.B(n_45),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_11),
.B(n_27),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_11),
.B(n_16),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_13),
.B(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_14),
.B(n_81),
.Y(n_80)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_14),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_25),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_15),
.B(n_41),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_15),
.B(n_27),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_15),
.B(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_16),
.Y(n_106)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_16),
.Y(n_146)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_16),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_112),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_74),
.B2(n_111),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_47),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_33),
.C(n_39),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_23),
.B(n_125),
.Y(n_124)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_23),
.Y(n_203)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_26),
.CI(n_29),
.CON(n_23),
.SN(n_23)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_24),
.B(n_26),
.C(n_29),
.Y(n_96)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_33),
.A2(n_34),
.B1(n_39),
.B2(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_39),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.C(n_44),
.Y(n_39)
);

FAx1_ASAP7_75t_SL g117 ( 
.A(n_40),
.B(n_43),
.CI(n_44),
.CON(n_117),
.SN(n_117)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_45),
.Y(n_182)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_57),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_55),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_66),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_65),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_72),
.C(n_73),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_68),
.B(n_182),
.Y(n_181)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_73),
.Y(n_77)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_94),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.C(n_85),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_76),
.A2(n_78),
.B1(n_79),
.B2(n_115),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_76),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B(n_84),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_83),
.Y(n_84)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_82),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_85),
.B(n_114),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_86),
.B(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_86),
.B(n_193),
.C(n_196),
.Y(n_197)
);

FAx1_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_88),
.CI(n_89),
.CON(n_86),
.SN(n_86)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_151)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_107),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.C(n_123),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_113),
.B(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_116),
.A2(n_123),
.B1(n_124),
.B2(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.C(n_122),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_117),
.B(n_194),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g202 ( 
.A(n_117),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_118),
.B(n_122),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.C(n_121),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_197),
.C(n_198),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_191),
.C(n_192),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_152),
.C(n_165),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_141),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_139),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_132),
.B(n_139),
.C(n_141),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.C(n_137),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_134),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_149),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_150),
.C(n_151),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_143),
.A2(n_144),
.B1(n_147),
.B2(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_164),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_156),
.A2(n_157),
.B1(n_164),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_187),
.C(n_188),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_174),
.C(n_179),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_172),
.C(n_173),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.C(n_183),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);


endmodule