module fake_jpeg_20969_n_177 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_SL g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_30),
.B1(n_29),
.B2(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_20),
.B1(n_30),
.B2(n_29),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_49),
.B1(n_50),
.B2(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_18),
.Y(n_68)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_20),
.B1(n_27),
.B2(n_24),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_20),
.B1(n_27),
.B2(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_55),
.B(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_40),
.B(n_38),
.C(n_16),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_22),
.B(n_23),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_74),
.Y(n_85)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_31),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_41),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g75 ( 
.A(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_48),
.B1(n_43),
.B2(n_51),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_79),
.B1(n_91),
.B2(n_64),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_24),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_51),
.B1(n_41),
.B2(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_92),
.Y(n_97)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_44),
.B1(n_25),
.B2(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_31),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_65),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_93),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_99),
.Y(n_121)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_63),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_107),
.Y(n_128)
);

NOR4xp25_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_25),
.C(n_28),
.D(n_36),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_91),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_65),
.B1(n_71),
.B2(n_64),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_106),
.B1(n_88),
.B2(n_83),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_95),
.B(n_14),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_112),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_75),
.Y(n_111)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_80),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_109),
.Y(n_113)
);

NOR3xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_118),
.C(n_125),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_78),
.B1(n_81),
.B2(n_86),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_116),
.B(n_119),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_115),
.A2(n_120),
.B1(n_116),
.B2(n_102),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_83),
.B1(n_79),
.B2(n_90),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_109),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_76),
.B1(n_58),
.B2(n_90),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_35),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_127),
.Y(n_130)
);

AOI322xp5_ASAP7_75t_SL g125 ( 
.A1(n_107),
.A2(n_14),
.A3(n_13),
.B1(n_10),
.B2(n_9),
.C1(n_7),
.C2(n_8),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_98),
.A2(n_94),
.B1(n_58),
.B2(n_15),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_100),
.B1(n_101),
.B2(n_54),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_112),
.B(n_108),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_135),
.Y(n_144)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_103),
.B(n_102),
.C(n_110),
.D(n_106),
.Y(n_133)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_137),
.C(n_131),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_104),
.B(n_105),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_105),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_141),
.B(n_100),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_137),
.A2(n_119),
.B(n_127),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_149),
.B(n_150),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_132),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_129),
.B(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_17),
.Y(n_159)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_140),
.C(n_36),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_157),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_147),
.A2(n_75),
.B1(n_134),
.B2(n_26),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_159),
.B1(n_149),
.B2(n_150),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_17),
.C(n_21),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_164),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_145),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_165),
.C(n_161),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_154),
.A2(n_158),
.B(n_155),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_1),
.B(n_3),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_7),
.B1(n_8),
.B2(n_4),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_164),
.C(n_35),
.Y(n_170)
);

NOR2x1_ASAP7_75t_SL g167 ( 
.A(n_162),
.B(n_17),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_3),
.B(n_5),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_3),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_169),
.C(n_35),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_172),
.B1(n_5),
.B2(n_6),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_174),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_175),
.A2(n_6),
.B(n_15),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_36),
.Y(n_177)
);


endmodule