module fake_ariane_2712_n_81 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_10, n_81);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_81;

wire n_56;
wire n_60;
wire n_64;
wire n_38;
wire n_47;
wire n_75;
wire n_67;
wire n_34;
wire n_69;
wire n_74;
wire n_33;
wire n_40;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_49;
wire n_20;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_79;
wire n_26;
wire n_46;
wire n_36;
wire n_72;
wire n_44;
wire n_30;
wire n_42;
wire n_31;
wire n_57;
wire n_70;
wire n_48;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_23;
wire n_61;
wire n_22;
wire n_43;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_68;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_35;
wire n_54;
wire n_25;

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

AND2x6_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

AND3x2_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_0),
.C(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_R g33 ( 
.A(n_7),
.B(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_4),
.B(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_24),
.B(n_22),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

OAI21x1_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_24),
.B(n_23),
.Y(n_45)
);

CKINVDCx11_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_39),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_21),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_21),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_1),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_41),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_3),
.B(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_55),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

OAI32xp33_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_53),
.A3(n_32),
.B1(n_47),
.B2(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

AOI221xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_61),
.B1(n_60),
.B2(n_63),
.C(n_62),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_45),
.B(n_34),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_46),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_45),
.B(n_33),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

OAI221xp5_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_34),
.B1(n_30),
.B2(n_25),
.C(n_45),
.Y(n_73)
);

NAND2x1p5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_34),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

NAND4xp75_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_33),
.C(n_25),
.D(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

OAI22x1_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_71),
.B1(n_25),
.B2(n_68),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

OR2x6_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_76),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_79),
.A2(n_25),
.B1(n_73),
.B2(n_80),
.Y(n_81)
);


endmodule