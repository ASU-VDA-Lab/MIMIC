module fake_jpeg_14218_n_97 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_97);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_97;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_13),
.B(n_8),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_10),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_47),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_26),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_1),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_27),
.B1(n_37),
.B2(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_2),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_43),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_55),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_37),
.B1(n_32),
.B2(n_34),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_32),
.B(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_33),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_64),
.B(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_66),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_44),
.B1(n_41),
.B2(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_39),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_2),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_16),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_75),
.Y(n_79)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_77),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_52),
.C(n_17),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_78),
.A2(n_52),
.B(n_6),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_81),
.B(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_3),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_7),
.B(n_11),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_73),
.B(n_15),
.Y(n_89)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_86),
.B(n_89),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_79),
.A2(n_77),
.B1(n_80),
.B2(n_85),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_85),
.B1(n_7),
.B2(n_24),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_89),
.C(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

NOR2xp67_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_90),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_20),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_25),
.Y(n_97)
);


endmodule