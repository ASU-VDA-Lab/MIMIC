module fake_jpeg_1388_n_212 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_212);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_3),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_6),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_8),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_15),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_5),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_35),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_11),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_70),
.Y(n_89)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_75),
.Y(n_86)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_61),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_78),
.B(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_85),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_49),
.B1(n_64),
.B2(n_53),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_69),
.B1(n_67),
.B2(n_52),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_63),
.Y(n_85)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_91),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_70),
.B1(n_60),
.B2(n_57),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_92),
.B1(n_51),
.B2(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_54),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_57),
.B1(n_55),
.B2(n_64),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_51),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_85),
.A2(n_76),
.B1(n_53),
.B2(n_74),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_103),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_66),
.B1(n_81),
.B2(n_2),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_50),
.Y(n_98)
);

XOR2x1_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_106),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_82),
.B1(n_87),
.B2(n_83),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_52),
.B1(n_77),
.B2(n_68),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_101),
.Y(n_118)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

NOR2x1_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_54),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_107),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_68),
.A3(n_56),
.B1(n_67),
.B2(n_69),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_58),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_110),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_62),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_45),
.Y(n_132)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_96),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_65),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_120),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_121),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_81),
.B(n_56),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_42),
.B(n_41),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_5),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_102),
.B(n_43),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_105),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_150),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_155),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_131),
.B(n_3),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_140),
.B(n_148),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_117),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_127),
.B(n_4),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_143),
.B(n_157),
.Y(n_160)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_147),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_39),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_149),
.C(n_150),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_123),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_125),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_122),
.B1(n_114),
.B2(n_115),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_36),
.B1(n_32),
.B2(n_31),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_151),
.A2(n_114),
.B1(n_115),
.B2(n_133),
.Y(n_158)
);

OAI211xp5_ASAP7_75t_SL g152 ( 
.A1(n_129),
.A2(n_30),
.B(n_29),
.C(n_27),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_130),
.B(n_9),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_154),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_26),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_121),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_135),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_159),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_142),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_135),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_18),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_154),
.B(n_136),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_150),
.C(n_155),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_115),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_173),
.Y(n_182)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_128),
.C(n_25),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_137),
.A2(n_12),
.B(n_13),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_177),
.A2(n_178),
.B(n_144),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_24),
.B(n_22),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_179),
.A2(n_187),
.B1(n_163),
.B2(n_174),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_174),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_166),
.A2(n_14),
.B(n_15),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_186),
.B(n_177),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_20),
.B(n_16),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_169),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_176),
.B(n_17),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_188),
.Y(n_196)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_181),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_192),
.B(n_193),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_164),
.C(n_165),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_197),
.C(n_198),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_190),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_170),
.C(n_172),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_182),
.C(n_183),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_201),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_168),
.C(n_175),
.Y(n_203)
);

NOR4xp25_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_161),
.C(n_160),
.D(n_179),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_202),
.A2(n_194),
.B(n_158),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_206),
.B(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_205),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_208),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_199),
.C(n_187),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_210),
.A2(n_196),
.B(n_20),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_211),
.Y(n_212)
);


endmodule