module real_aes_8568_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_310;
wire n_119;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_0), .A2(n_43), .B1(n_136), .B2(n_139), .Y(n_135) );
INVx1_ASAP7_75t_L g111 ( .A(n_1), .Y(n_111) );
INVx1_ASAP7_75t_L g264 ( .A(n_2), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_3), .B(n_124), .Y(n_123) );
AOI21xp33_ASAP7_75t_L g244 ( .A1(n_4), .A2(n_202), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g185 ( .A(n_5), .Y(n_185) );
AND2x6_ASAP7_75t_L g207 ( .A(n_5), .B(n_183), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_5), .B(n_518), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_6), .A2(n_303), .B(n_304), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g81 ( .A1(n_7), .A2(n_82), .B1(n_83), .B2(n_86), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_7), .Y(n_82) );
INVx1_ASAP7_75t_L g251 ( .A(n_8), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_9), .B(n_295), .Y(n_294) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_10), .A2(n_25), .B1(n_101), .B2(n_102), .Y(n_100) );
INVx1_ASAP7_75t_L g200 ( .A(n_11), .Y(n_200) );
INVx1_ASAP7_75t_L g309 ( .A(n_12), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_13), .B(n_215), .Y(n_320) );
AO22x2_ASAP7_75t_L g104 ( .A1(n_14), .A2(n_26), .B1(n_101), .B2(n_105), .Y(n_104) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_15), .A2(n_31), .B1(n_168), .B2(n_171), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_16), .B(n_202), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_17), .B(n_223), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g306 ( .A1(n_18), .A2(n_307), .B(n_308), .C(n_310), .Y(n_306) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_19), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_20), .B(n_249), .Y(n_266) );
AOI22xp33_ASAP7_75t_SL g112 ( .A1(n_21), .A2(n_73), .B1(n_113), .B2(n_119), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_22), .B(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g238 ( .A(n_23), .Y(n_238) );
INVx2_ASAP7_75t_L g205 ( .A(n_24), .Y(n_205) );
OAI221xp5_ASAP7_75t_L g176 ( .A1(n_26), .A2(n_38), .B1(n_47), .B2(n_177), .C(n_178), .Y(n_176) );
INVxp67_ASAP7_75t_L g179 ( .A(n_26), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g276 ( .A1(n_27), .A2(n_207), .B(n_210), .C(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g236 ( .A(n_28), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_29), .A2(n_32), .B1(n_161), .B2(n_164), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_30), .B(n_249), .Y(n_319) );
CKINVDCx16_ASAP7_75t_R g239 ( .A(n_33), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_34), .B(n_202), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_35), .A2(n_210), .B1(n_232), .B2(n_234), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g285 ( .A(n_36), .Y(n_285) );
CKINVDCx16_ASAP7_75t_R g261 ( .A(n_37), .Y(n_261) );
AO22x2_ASAP7_75t_L g108 ( .A1(n_38), .A2(n_57), .B1(n_101), .B2(n_105), .Y(n_108) );
INVxp67_ASAP7_75t_L g180 ( .A(n_38), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_39), .A2(n_219), .B(n_248), .C(n_250), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_40), .Y(n_323) );
INVx1_ASAP7_75t_L g246 ( .A(n_41), .Y(n_246) );
INVx1_ASAP7_75t_L g183 ( .A(n_42), .Y(n_183) );
INVx1_ASAP7_75t_L g199 ( .A(n_44), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_45), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_46), .A2(n_91), .B1(n_92), .B2(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_46), .Y(n_526) );
AO22x2_ASAP7_75t_L g110 ( .A1(n_47), .A2(n_62), .B1(n_101), .B2(n_102), .Y(n_110) );
AOI22xp33_ASAP7_75t_SL g144 ( .A1(n_48), .A2(n_64), .B1(n_145), .B2(n_149), .Y(n_144) );
AOI22xp33_ASAP7_75t_SL g153 ( .A1(n_49), .A2(n_52), .B1(n_154), .B2(n_157), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_SL g214 ( .A1(n_50), .A2(n_215), .B(n_216), .C(n_219), .Y(n_214) );
INVxp67_ASAP7_75t_L g217 ( .A(n_51), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_53), .Y(n_242) );
INVx1_ASAP7_75t_L g316 ( .A(n_54), .Y(n_316) );
INVx1_ASAP7_75t_L g524 ( .A(n_54), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g317 ( .A1(n_55), .A2(n_207), .B(n_210), .C(n_318), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_55), .A2(n_91), .B1(n_92), .B2(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_55), .Y(n_514) );
INVx1_ASAP7_75t_L g90 ( .A(n_56), .Y(n_90) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_58), .B(n_265), .Y(n_278) );
INVx2_ASAP7_75t_L g197 ( .A(n_59), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_60), .B(n_215), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_61), .A2(n_207), .B(n_210), .C(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_63), .B(n_253), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_65), .Y(n_269) );
OAI22xp5_ASAP7_75t_SL g79 ( .A1(n_66), .A2(n_80), .B1(n_81), .B2(n_87), .Y(n_79) );
INVx1_ASAP7_75t_L g87 ( .A(n_66), .Y(n_87) );
A2O1A1Ixp33_ASAP7_75t_L g291 ( .A1(n_66), .A2(n_207), .B(n_210), .C(n_292), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g299 ( .A(n_67), .Y(n_299) );
INVx1_ASAP7_75t_L g213 ( .A(n_68), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g305 ( .A(n_69), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_70), .B(n_265), .Y(n_293) );
INVx1_ASAP7_75t_L g101 ( .A(n_71), .Y(n_101) );
INVx1_ASAP7_75t_L g103 ( .A(n_71), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g83 ( .A1(n_72), .A2(n_75), .B1(n_84), .B2(n_85), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_72), .Y(n_84) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_74), .B(n_195), .Y(n_311) );
INVx1_ASAP7_75t_L g85 ( .A(n_75), .Y(n_85) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_76), .A2(n_202), .B(n_208), .Y(n_201) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_173), .B1(n_186), .B2(n_511), .C(n_512), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_88), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_83), .Y(n_86) );
AOI22xp5_ASAP7_75t_L g88 ( .A1(n_89), .A2(n_90), .B1(n_91), .B2(n_92), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_92), .Y(n_91) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
NAND2xp5_ASAP7_75t_SL g93 ( .A(n_94), .B(n_142), .Y(n_93) );
NOR2xp33_ASAP7_75t_L g94 ( .A(n_95), .B(n_122), .Y(n_94) );
OAI21xp5_ASAP7_75t_SL g95 ( .A1(n_96), .A2(n_111), .B(n_112), .Y(n_95) );
INVx3_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
BUFx3_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x6_ASAP7_75t_L g98 ( .A(n_99), .B(n_106), .Y(n_98) );
AND2x4_ASAP7_75t_L g139 ( .A(n_99), .B(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g99 ( .A(n_100), .B(n_104), .Y(n_99) );
AND2x2_ASAP7_75t_L g118 ( .A(n_100), .B(n_108), .Y(n_118) );
INVx2_ASAP7_75t_L g127 ( .A(n_100), .Y(n_127) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g105 ( .A(n_103), .Y(n_105) );
INVx2_ASAP7_75t_L g117 ( .A(n_104), .Y(n_117) );
AND2x2_ASAP7_75t_L g126 ( .A(n_104), .B(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g134 ( .A(n_104), .B(n_127), .Y(n_134) );
INVx1_ASAP7_75t_L g138 ( .A(n_104), .Y(n_138) );
AND2x6_ASAP7_75t_L g163 ( .A(n_106), .B(n_133), .Y(n_163) );
AND2x4_ASAP7_75t_L g166 ( .A(n_106), .B(n_126), .Y(n_166) );
AND2x2_ASAP7_75t_L g170 ( .A(n_106), .B(n_148), .Y(n_170) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
AND2x2_ASAP7_75t_L g128 ( .A(n_107), .B(n_110), .Y(n_128) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g147 ( .A(n_108), .B(n_141), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_108), .B(n_110), .Y(n_152) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g116 ( .A(n_110), .Y(n_116) );
INVx1_ASAP7_75t_L g141 ( .A(n_110), .Y(n_141) );
BUFx4f_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
INVx1_ASAP7_75t_L g121 ( .A(n_116), .Y(n_121) );
AND2x2_ASAP7_75t_L g148 ( .A(n_117), .B(n_127), .Y(n_148) );
INVx1_ASAP7_75t_L g158 ( .A(n_117), .Y(n_158) );
AND2x4_ASAP7_75t_L g120 ( .A(n_118), .B(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g136 ( .A(n_118), .B(n_137), .Y(n_136) );
BUFx12f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND3xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_129), .C(n_135), .Y(n_122) );
BUFx4f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_128), .Y(n_125) );
AND2x2_ASAP7_75t_L g156 ( .A(n_126), .B(n_147), .Y(n_156) );
AND2x4_ASAP7_75t_L g132 ( .A(n_128), .B(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g172 ( .A(n_128), .B(n_148), .Y(n_172) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx4_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_143), .B(n_159), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_153), .Y(n_143) );
BUFx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x4_ASAP7_75t_L g150 ( .A(n_148), .B(n_151), .Y(n_150) );
BUFx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g157 ( .A(n_151), .B(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx8_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_167), .Y(n_159) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx11_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx6_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_174), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
AND3x1_ASAP7_75t_SL g175 ( .A(n_176), .B(n_181), .C(n_184), .Y(n_175) );
INVxp67_ASAP7_75t_L g518 ( .A(n_176), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_181), .Y(n_519) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_181), .A2(n_203), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g528 ( .A(n_181), .Y(n_528) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_182), .B(n_185), .Y(n_523) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
OR2x2_ASAP7_75t_SL g527 ( .A(n_184), .B(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_SL g187 ( .A(n_188), .B(n_448), .Y(n_187) );
NOR4xp25_ASAP7_75t_L g188 ( .A(n_189), .B(n_378), .C(n_409), .D(n_428), .Y(n_188) );
NAND4xp25_ASAP7_75t_L g189 ( .A(n_190), .B(n_336), .C(n_351), .D(n_369), .Y(n_189) );
AOI222xp33_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_271), .B1(n_312), .B2(n_324), .C1(n_329), .C2(n_331), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_192), .B(n_254), .Y(n_191) );
INVx1_ASAP7_75t_L g392 ( .A(n_192), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_225), .Y(n_192) );
AND2x2_ASAP7_75t_L g255 ( .A(n_193), .B(n_243), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_193), .B(n_258), .Y(n_421) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
OR2x2_ASAP7_75t_L g328 ( .A(n_194), .B(n_227), .Y(n_328) );
AND2x2_ASAP7_75t_L g337 ( .A(n_194), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g363 ( .A(n_194), .Y(n_363) );
AND2x2_ASAP7_75t_L g384 ( .A(n_194), .B(n_227), .Y(n_384) );
BUFx2_ASAP7_75t_L g407 ( .A(n_194), .Y(n_407) );
AND2x2_ASAP7_75t_L g431 ( .A(n_194), .B(n_228), .Y(n_431) );
AND2x2_ASAP7_75t_L g495 ( .A(n_194), .B(n_243), .Y(n_495) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_201), .B(n_222), .Y(n_194) );
INVx4_ASAP7_75t_L g224 ( .A(n_195), .Y(n_224) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g229 ( .A(n_196), .Y(n_229) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
AND2x2_ASAP7_75t_SL g253 ( .A(n_197), .B(n_198), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
BUFx2_ASAP7_75t_L g303 ( .A(n_202), .Y(n_303) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_207), .Y(n_202) );
NAND2x1p5_ASAP7_75t_L g240 ( .A(n_203), .B(n_207), .Y(n_240) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_206), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g211 ( .A(n_205), .Y(n_211) );
INVx1_ASAP7_75t_L g233 ( .A(n_205), .Y(n_233) );
INVx1_ASAP7_75t_L g212 ( .A(n_206), .Y(n_212) );
INVx1_ASAP7_75t_L g215 ( .A(n_206), .Y(n_215) );
INVx3_ASAP7_75t_L g218 ( .A(n_206), .Y(n_218) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_206), .Y(n_235) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_206), .Y(n_249) );
INVx4_ASAP7_75t_SL g221 ( .A(n_207), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_213), .B(n_214), .C(n_221), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_209), .A2(n_221), .B(n_246), .C(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g304 ( .A1(n_209), .A2(n_221), .B(n_305), .C(n_306), .Y(n_304) );
INVx5_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x6_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_211), .Y(n_220) );
BUFx3_ASAP7_75t_L g282 ( .A(n_211), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_218), .B(n_251), .Y(n_250) );
INVx5_ASAP7_75t_L g265 ( .A(n_218), .Y(n_265) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_220), .Y(n_296) );
OAI22xp33_ASAP7_75t_L g230 ( .A1(n_221), .A2(n_231), .B1(n_239), .B2(n_240), .Y(n_230) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_223), .A2(n_244), .B(n_252), .Y(n_243) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_SL g284 ( .A(n_224), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g396 ( .A(n_225), .B(n_327), .Y(n_396) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_226), .B(n_421), .Y(n_420) );
OR2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_243), .Y(n_226) );
OR2x2_ASAP7_75t_L g356 ( .A(n_227), .B(n_259), .Y(n_356) );
AND2x2_ASAP7_75t_L g368 ( .A(n_227), .B(n_327), .Y(n_368) );
BUFx2_ASAP7_75t_L g500 ( .A(n_227), .Y(n_500) );
INVx3_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
OR2x2_ASAP7_75t_L g257 ( .A(n_228), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g350 ( .A(n_228), .B(n_259), .Y(n_350) );
AND2x2_ASAP7_75t_L g403 ( .A(n_228), .B(n_243), .Y(n_403) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_228), .Y(n_439) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_241), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_229), .B(n_242), .Y(n_241) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_229), .A2(n_260), .B(n_268), .Y(n_259) );
INVx2_ASAP7_75t_L g283 ( .A(n_229), .Y(n_283) );
INVx2_ASAP7_75t_L g267 ( .A(n_232), .Y(n_267) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
OAI22xp5_ASAP7_75t_SL g234 ( .A1(n_235), .A2(n_236), .B1(n_237), .B2(n_238), .Y(n_234) );
INVx2_ASAP7_75t_L g237 ( .A(n_235), .Y(n_237) );
INVx4_ASAP7_75t_L g307 ( .A(n_235), .Y(n_307) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_240), .A2(n_261), .B(n_262), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g315 ( .A1(n_240), .A2(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_L g326 ( .A(n_243), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g338 ( .A(n_243), .Y(n_338) );
INVx2_ASAP7_75t_L g349 ( .A(n_243), .Y(n_349) );
BUFx2_ASAP7_75t_L g373 ( .A(n_243), .Y(n_373) );
AND2x2_ASAP7_75t_SL g430 ( .A(n_243), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx4_ASAP7_75t_L g295 ( .A(n_249), .Y(n_295) );
INVx1_ASAP7_75t_L g270 ( .A(n_253), .Y(n_270) );
INVx2_ASAP7_75t_L g289 ( .A(n_253), .Y(n_289) );
OA21x2_ASAP7_75t_L g301 ( .A1(n_253), .A2(n_302), .B(n_311), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
AOI332xp33_ASAP7_75t_L g351 ( .A1(n_255), .A2(n_352), .A3(n_356), .B1(n_357), .B2(n_361), .B3(n_364), .C1(n_365), .C2(n_367), .Y(n_351) );
NAND2x1_ASAP7_75t_L g436 ( .A(n_255), .B(n_327), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_255), .B(n_341), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_SL g369 ( .A1(n_256), .A2(n_370), .B(n_373), .C(n_374), .Y(n_369) );
AND2x2_ASAP7_75t_L g508 ( .A(n_256), .B(n_349), .Y(n_508) );
INVx3_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g405 ( .A(n_257), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g410 ( .A(n_257), .B(n_407), .Y(n_410) );
INVx1_ASAP7_75t_L g341 ( .A(n_258), .Y(n_341) );
AND2x2_ASAP7_75t_L g444 ( .A(n_258), .B(n_403), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_258), .B(n_384), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_258), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_258), .B(n_362), .Y(n_470) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g327 ( .A(n_259), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_265), .B(n_266), .C(n_267), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_270), .B(n_299), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_270), .B(n_323), .Y(n_322) );
OAI31xp33_ASAP7_75t_L g509 ( .A1(n_271), .A2(n_430), .A3(n_437), .B(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_286), .Y(n_271) );
AND2x2_ASAP7_75t_L g312 ( .A(n_272), .B(n_313), .Y(n_312) );
NAND2x1_ASAP7_75t_SL g332 ( .A(n_272), .B(n_333), .Y(n_332) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_272), .Y(n_419) );
AND2x2_ASAP7_75t_L g424 ( .A(n_272), .B(n_335), .Y(n_424) );
INVx3_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_273), .A2(n_337), .B(n_339), .C(n_342), .Y(n_336) );
OR2x2_ASAP7_75t_L g353 ( .A(n_273), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g366 ( .A(n_273), .Y(n_366) );
AND2x2_ASAP7_75t_L g372 ( .A(n_273), .B(n_314), .Y(n_372) );
INVx2_ASAP7_75t_L g390 ( .A(n_273), .Y(n_390) );
AND2x2_ASAP7_75t_L g401 ( .A(n_273), .B(n_355), .Y(n_401) );
AND2x2_ASAP7_75t_L g433 ( .A(n_273), .B(n_391), .Y(n_433) );
AND2x2_ASAP7_75t_L g437 ( .A(n_273), .B(n_360), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_273), .B(n_286), .Y(n_442) );
AND2x2_ASAP7_75t_L g476 ( .A(n_273), .B(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_273), .B(n_379), .Y(n_510) );
OR2x6_ASAP7_75t_L g273 ( .A(n_274), .B(n_284), .Y(n_273) );
AOI21xp5_ASAP7_75t_SL g274 ( .A1(n_275), .A2(n_276), .B(n_283), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_279), .B(n_280), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_280), .A2(n_319), .B(n_320), .Y(n_318) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g310 ( .A(n_282), .Y(n_310) );
INVx1_ASAP7_75t_L g321 ( .A(n_283), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_286), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g418 ( .A(n_286), .Y(n_418) );
AND2x2_ASAP7_75t_L g480 ( .A(n_286), .B(n_401), .Y(n_480) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_300), .Y(n_286) );
OR2x2_ASAP7_75t_L g334 ( .A(n_287), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g344 ( .A(n_287), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_287), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g452 ( .A(n_287), .Y(n_452) );
AND2x2_ASAP7_75t_L g469 ( .A(n_287), .B(n_314), .Y(n_469) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g360 ( .A(n_288), .B(n_300), .Y(n_360) );
AND2x2_ASAP7_75t_L g389 ( .A(n_288), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g400 ( .A(n_288), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_288), .B(n_355), .Y(n_491) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_290), .B(n_298), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_297), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B(n_296), .Y(n_292) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g313 ( .A(n_301), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g335 ( .A(n_301), .Y(n_335) );
AND2x2_ASAP7_75t_L g391 ( .A(n_301), .B(n_355), .Y(n_391) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_303), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_307), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g493 ( .A(n_312), .Y(n_493) );
INVx1_ASAP7_75t_L g497 ( .A(n_313), .Y(n_497) );
INVx2_ASAP7_75t_L g355 ( .A(n_314), .Y(n_355) );
AO21x2_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_321), .B(n_322), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_325), .B(n_328), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_326), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_326), .B(n_431), .Y(n_489) );
OR2x2_ASAP7_75t_L g330 ( .A(n_327), .B(n_328), .Y(n_330) );
INVx1_ASAP7_75t_SL g382 ( .A(n_327), .Y(n_382) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_333), .A2(n_386), .B1(n_388), .B2(n_392), .C(n_393), .Y(n_385) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g413 ( .A(n_334), .B(n_377), .Y(n_413) );
INVx2_ASAP7_75t_L g345 ( .A(n_335), .Y(n_345) );
INVx1_ASAP7_75t_L g371 ( .A(n_335), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_335), .B(n_355), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_335), .B(n_358), .Y(n_465) );
INVx1_ASAP7_75t_L g473 ( .A(n_335), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_337), .B(n_341), .Y(n_387) );
AND2x4_ASAP7_75t_L g362 ( .A(n_338), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g475 ( .A(n_341), .B(n_431), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_346), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_344), .B(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_L g483 ( .A(n_345), .Y(n_483) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g383 ( .A(n_349), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g455 ( .A(n_349), .B(n_431), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_349), .B(n_368), .Y(n_461) );
AOI322xp5_ASAP7_75t_L g415 ( .A1(n_350), .A2(n_384), .A3(n_391), .B1(n_416), .B2(n_419), .C1(n_420), .C2(n_422), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_350), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g481 ( .A(n_353), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g427 ( .A(n_354), .Y(n_427) );
INVx2_ASAP7_75t_L g358 ( .A(n_355), .Y(n_358) );
INVx1_ASAP7_75t_L g417 ( .A(n_355), .Y(n_417) );
CKINVDCx16_ASAP7_75t_R g364 ( .A(n_356), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
AND2x2_ASAP7_75t_L g453 ( .A(n_358), .B(n_366), .Y(n_453) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g365 ( .A(n_360), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g408 ( .A(n_360), .B(n_401), .Y(n_408) );
AND2x2_ASAP7_75t_L g412 ( .A(n_360), .B(n_372), .Y(n_412) );
OAI21xp33_ASAP7_75t_SL g422 ( .A1(n_361), .A2(n_423), .B(n_425), .Y(n_422) );
OAI22xp33_ASAP7_75t_L g492 ( .A1(n_361), .A2(n_493), .B1(n_494), .B2(n_496), .Y(n_492) );
INVx3_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g367 ( .A(n_362), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_362), .B(n_382), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_364), .B(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
INVx1_ASAP7_75t_L g504 ( .A(n_371), .Y(n_504) );
INVx4_ASAP7_75t_L g377 ( .A(n_372), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_372), .B(n_399), .Y(n_447) );
INVx1_ASAP7_75t_SL g459 ( .A(n_373), .Y(n_459) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NOR2xp67_ASAP7_75t_L g472 ( .A(n_377), .B(n_473), .Y(n_472) );
OAI211xp5_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_380), .B(n_385), .C(n_402), .Y(n_378) );
OAI221xp5_ASAP7_75t_SL g498 ( .A1(n_380), .A2(n_418), .B1(n_497), .B2(n_499), .C(n_501), .Y(n_498) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_382), .B(n_495), .Y(n_494) );
OAI31xp33_ASAP7_75t_L g474 ( .A1(n_383), .A2(n_460), .A3(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g414 ( .A(n_384), .Y(n_414) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
INVx1_ASAP7_75t_L g464 ( .A(n_389), .Y(n_464) );
AND2x2_ASAP7_75t_L g477 ( .A(n_391), .B(n_400), .Y(n_477) );
AOI21xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B(n_397), .Y(n_393) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_401), .B(n_504), .Y(n_503) );
OAI21xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B(n_408), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI221xp5_ASAP7_75t_SL g409 ( .A1(n_410), .A2(n_411), .B1(n_413), .B2(n_414), .C(n_415), .Y(n_409) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_410), .A2(n_479), .B(n_481), .C(n_484), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_413), .B(n_463), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g440 ( .A(n_421), .Y(n_440) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g426 ( .A(n_424), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g468 ( .A(n_424), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI211xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_432), .B(n_434), .C(n_443), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI221xp5_ASAP7_75t_L g505 ( .A1(n_432), .A2(n_442), .B1(n_506), .B2(n_507), .C(n_509), .Y(n_505) );
INVx1_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B1(n_438), .B2(n_441), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI21xp5_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_445), .B(n_446), .Y(n_443) );
INVx1_ASAP7_75t_SL g506 ( .A(n_445), .Y(n_506) );
INVxp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NOR4xp25_ASAP7_75t_L g448 ( .A(n_449), .B(n_478), .C(n_498), .D(n_505), .Y(n_448) );
OAI211xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_454), .B(n_456), .C(n_474), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_453), .Y(n_450) );
INVxp67_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_460), .B(n_462), .C(n_466), .Y(n_456) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_SL g485 ( .A(n_463), .Y(n_485) );
OR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
OR2x2_ASAP7_75t_L g496 ( .A(n_464), .B(n_497), .Y(n_496) );
OAI21xp33_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_470), .B(n_471), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_488), .B2(n_490), .C(n_492), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVxp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_495), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OAI322xp33_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_515), .A3(n_519), .B1(n_520), .B2(n_524), .C1(n_525), .C2(n_527), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_522), .Y(n_521) );
endmodule