module fake_jpeg_10308_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_3),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_6),
.B(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_14),
.A2(n_10),
.B1(n_11),
.B2(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

OA22x2_ASAP7_75t_L g19 ( 
.A1(n_16),
.A2(n_17),
.B1(n_15),
.B2(n_11),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_19),
.A2(n_10),
.B1(n_13),
.B2(n_8),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_18),
.B(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_8),
.C(n_7),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_24),
.B(n_25),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_20),
.C(n_17),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_19),
.B1(n_13),
.B2(n_14),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_19),
.C(n_7),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_32),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_19),
.B(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_5),
.C(n_14),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_5),
.Y(n_37)
);

AOI322xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_35),
.A3(n_13),
.B1(n_3),
.B2(n_2),
.C1(n_1),
.C2(n_14),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_1),
.Y(n_40)
);


endmodule