module fake_aes_2800_n_686 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_686);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_686;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g78 ( .A(n_21), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_27), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_13), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_4), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_32), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_12), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_43), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_66), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_15), .Y(n_86) );
BUFx3_ASAP7_75t_L g87 ( .A(n_36), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_49), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_57), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_59), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_15), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_31), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_67), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_53), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_41), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_44), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_73), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_61), .Y(n_98) );
HB1xp67_ASAP7_75t_L g99 ( .A(n_25), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_14), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_45), .B(n_56), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_72), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_7), .Y(n_103) );
INVx2_ASAP7_75t_SL g104 ( .A(n_35), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_6), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_63), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_8), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_37), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_13), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_38), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_55), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_42), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_3), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_22), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_33), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_9), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_30), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_64), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_40), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_12), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_65), .Y(n_121) );
HB1xp67_ASAP7_75t_SL g122 ( .A(n_34), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_47), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_16), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_3), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_81), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_79), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_82), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_82), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_85), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_110), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_113), .B(n_0), .Y(n_133) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_85), .A2(n_28), .B(n_76), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_110), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_88), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_110), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_81), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_113), .B(n_0), .Y(n_139) );
BUFx3_ASAP7_75t_L g140 ( .A(n_87), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_88), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_90), .Y(n_142) );
INVxp67_ASAP7_75t_L g143 ( .A(n_99), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_110), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_90), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_92), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_110), .Y(n_147) );
OAI22xp5_ASAP7_75t_L g148 ( .A1(n_109), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_89), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_87), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_102), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_92), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_93), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_80), .B(n_1), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_93), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_89), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_95), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_119), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_104), .B(n_2), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_102), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_104), .B(n_5), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_95), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_119), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_97), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_97), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_98), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_80), .B(n_125), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_98), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_143), .B(n_106), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_168), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_143), .B(n_125), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_168), .Y(n_172) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_133), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_127), .B(n_100), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_127), .B(n_100), .Y(n_176) );
INVx4_ASAP7_75t_L g177 ( .A(n_140), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_150), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_154), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_154), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_154), .Y(n_181) );
BUFx10_ASAP7_75t_L g182 ( .A(n_161), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_150), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_159), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_159), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_128), .B(n_121), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_128), .B(n_111), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_129), .B(n_121), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_129), .B(n_86), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_144), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_140), .Y(n_191) );
OR2x2_ASAP7_75t_L g192 ( .A(n_133), .B(n_116), .Y(n_192) );
INVx5_ASAP7_75t_L g193 ( .A(n_150), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_144), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_130), .B(n_86), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_150), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_130), .B(n_83), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_141), .Y(n_198) );
INVxp67_ASAP7_75t_SL g199 ( .A(n_139), .Y(n_199) );
NAND2x1p5_ASAP7_75t_L g200 ( .A(n_131), .B(n_83), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_168), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_150), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_141), .Y(n_203) );
BUFx3_ASAP7_75t_L g204 ( .A(n_150), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_141), .Y(n_205) );
INVx4_ASAP7_75t_L g206 ( .A(n_141), .Y(n_206) );
BUFx2_ASAP7_75t_L g207 ( .A(n_139), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_153), .Y(n_208) );
INVx4_ASAP7_75t_L g209 ( .A(n_153), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_131), .B(n_114), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_153), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_167), .B(n_120), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_153), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_144), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_136), .B(n_116), .Y(n_215) );
AND2x6_ASAP7_75t_L g216 ( .A(n_136), .B(n_123), .Y(n_216) );
NAND2x1p5_ASAP7_75t_L g217 ( .A(n_142), .B(n_114), .Y(n_217) );
INVx1_ASAP7_75t_SL g218 ( .A(n_167), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_142), .B(n_145), .Y(n_219) );
OR2x2_ASAP7_75t_L g220 ( .A(n_145), .B(n_120), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_146), .Y(n_221) );
NOR2xp33_ASAP7_75t_SL g222 ( .A(n_148), .B(n_94), .Y(n_222) );
AND3x4_ASAP7_75t_L g223 ( .A(n_148), .B(n_124), .C(n_122), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_146), .B(n_123), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_152), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_152), .B(n_118), .Y(n_226) );
AND2x6_ASAP7_75t_L g227 ( .A(n_155), .B(n_117), .Y(n_227) );
INVx4_ASAP7_75t_L g228 ( .A(n_151), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_144), .Y(n_229) );
NAND2xp33_ASAP7_75t_SL g230 ( .A(n_155), .B(n_157), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_157), .Y(n_231) );
AND2x6_ASAP7_75t_L g232 ( .A(n_184), .B(n_115), .Y(n_232) );
INVx2_ASAP7_75t_SL g233 ( .A(n_218), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_207), .A2(n_166), .B1(n_165), .B2(n_164), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_200), .Y(n_235) );
BUFx6f_ASAP7_75t_SL g236 ( .A(n_175), .Y(n_236) );
INVx5_ASAP7_75t_L g237 ( .A(n_206), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_200), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_199), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_185), .B(n_162), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_173), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_207), .Y(n_242) );
AND3x2_ASAP7_75t_SL g243 ( .A(n_223), .B(n_158), .C(n_156), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_216), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_217), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_179), .B(n_162), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_186), .B(n_164), .Y(n_247) );
INVxp67_ASAP7_75t_L g248 ( .A(n_188), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_230), .A2(n_166), .B1(n_165), .B2(n_91), .Y(n_249) );
AND2x6_ASAP7_75t_L g250 ( .A(n_180), .B(n_118), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_181), .B(n_126), .Y(n_251) );
INVx2_ASAP7_75t_SL g252 ( .A(n_212), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_206), .B(n_163), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_171), .B(n_126), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_217), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_217), .Y(n_256) );
AO22x1_ASAP7_75t_L g257 ( .A1(n_223), .A2(n_78), .B1(n_112), .B2(n_84), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_230), .A2(n_149), .B(n_163), .C(n_158), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_212), .B(n_206), .Y(n_259) );
INVx2_ASAP7_75t_SL g260 ( .A(n_192), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_209), .Y(n_261) );
INVx1_ASAP7_75t_SL g262 ( .A(n_216), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_169), .A2(n_103), .B1(n_105), .B2(n_107), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_191), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_209), .Y(n_265) );
INVx4_ASAP7_75t_SL g266 ( .A(n_216), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_209), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_192), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_175), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_175), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_176), .Y(n_271) );
NOR2xp33_ASAP7_75t_SL g272 ( .A(n_216), .B(n_96), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_216), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_171), .B(n_138), .Y(n_274) );
O2A1O1Ixp5_ASAP7_75t_L g275 ( .A1(n_174), .A2(n_108), .B(n_117), .C(n_115), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_176), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_216), .A2(n_168), .B1(n_163), .B2(n_149), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_176), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_182), .B(n_126), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_221), .B(n_149), .Y(n_280) );
INVx5_ASAP7_75t_L g281 ( .A(n_227), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_191), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_227), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_225), .B(n_156), .Y(n_284) );
AOI21x1_ASAP7_75t_L g285 ( .A1(n_231), .A2(n_134), .B(n_158), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_219), .B(n_138), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_174), .Y(n_287) );
CKINVDCx8_ASAP7_75t_R g288 ( .A(n_227), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_189), .B(n_138), .Y(n_289) );
AND2x2_ASAP7_75t_SL g290 ( .A(n_222), .B(n_134), .Y(n_290) );
INVx3_ASAP7_75t_L g291 ( .A(n_220), .Y(n_291) );
OR2x6_ASAP7_75t_L g292 ( .A(n_220), .B(n_138), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_189), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_182), .B(n_126), .Y(n_294) );
BUFx2_ASAP7_75t_L g295 ( .A(n_227), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_227), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_195), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_195), .B(n_156), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_244), .Y(n_299) );
BUFx12f_ASAP7_75t_L g300 ( .A(n_233), .Y(n_300) );
CKINVDCx20_ASAP7_75t_R g301 ( .A(n_268), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_252), .A2(n_224), .B1(n_226), .B2(n_208), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_244), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_237), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_240), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_240), .B(n_197), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_260), .Y(n_307) );
BUFx3_ASAP7_75t_L g308 ( .A(n_237), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_241), .B(n_197), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_291), .B(n_215), .Y(n_310) );
INVxp67_ASAP7_75t_L g311 ( .A(n_236), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_292), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_245), .B(n_174), .Y(n_313) );
O2A1O1Ixp5_ASAP7_75t_L g314 ( .A1(n_275), .A2(n_177), .B(n_187), .C(n_210), .Y(n_314) );
NAND2x2_ASAP7_75t_L g315 ( .A(n_257), .B(n_204), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_255), .A2(n_227), .B1(n_182), .B2(n_215), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_291), .A2(n_198), .B1(n_213), .B2(n_211), .Y(n_317) );
INVx2_ASAP7_75t_SL g318 ( .A(n_292), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_256), .A2(n_203), .B1(n_205), .B2(n_177), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_292), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_259), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_236), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_237), .Y(n_323) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_274), .A2(n_168), .B(n_132), .C(n_135), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_232), .Y(n_325) );
INVx4_ASAP7_75t_L g326 ( .A(n_244), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_235), .B(n_177), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_273), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_239), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_269), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_270), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_238), .A2(n_168), .B1(n_228), .B2(n_134), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_296), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_266), .B(n_228), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_234), .A2(n_228), .B1(n_134), .B2(n_151), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_248), .B(n_151), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_242), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_232), .A2(n_134), .B1(n_172), .B2(n_201), .Y(n_338) );
CKINVDCx16_ASAP7_75t_R g339 ( .A(n_272), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_261), .Y(n_340) );
BUFx3_ASAP7_75t_L g341 ( .A(n_281), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_288), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_293), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_232), .Y(n_344) );
INVx3_ASAP7_75t_L g345 ( .A(n_281), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_271), .Y(n_346) );
A2O1A1Ixp33_ASAP7_75t_L g347 ( .A1(n_247), .A2(n_135), .B(n_132), .C(n_147), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_265), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_276), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_281), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_339), .A2(n_290), .B1(n_278), .B2(n_298), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_307), .A2(n_250), .B1(n_232), .B2(n_254), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_301), .A2(n_250), .B1(n_254), .B2(n_297), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_301), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_321), .B(n_246), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_343), .A2(n_250), .B1(n_246), .B2(n_289), .Y(n_356) );
AOI22xp5_ASAP7_75t_SL g357 ( .A1(n_320), .A2(n_250), .B1(n_243), .B2(n_279), .Y(n_357) );
NAND2x1_ASAP7_75t_L g358 ( .A(n_299), .B(n_287), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_308), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_306), .B(n_289), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_329), .Y(n_361) );
BUFx4f_ASAP7_75t_L g362 ( .A(n_342), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_340), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_302), .A2(n_263), .B1(n_251), .B2(n_249), .C(n_294), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_340), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_337), .A2(n_251), .B1(n_267), .B2(n_249), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_348), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_348), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_305), .B(n_263), .Y(n_369) );
INVxp67_ASAP7_75t_L g370 ( .A(n_309), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_310), .A2(n_286), .B1(n_258), .B2(n_284), .C(n_280), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_312), .B(n_253), .Y(n_372) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_300), .A2(n_272), .B1(n_262), .B2(n_283), .Y(n_373) );
OAI22x1_ASAP7_75t_L g374 ( .A1(n_338), .A2(n_285), .B1(n_284), .B2(n_280), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_300), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_299), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_330), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_308), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_325), .A2(n_283), .B1(n_262), .B2(n_253), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_318), .B(n_295), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_322), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_327), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_368), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_363), .Y(n_384) );
HB1xp67_ASAP7_75t_SL g385 ( .A(n_375), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_372), .B(n_331), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_364), .A2(n_315), .B1(n_344), .B2(n_346), .Y(n_387) );
BUFx2_ASAP7_75t_L g388 ( .A(n_363), .Y(n_388) );
AO21x2_ASAP7_75t_L g389 ( .A1(n_351), .A2(n_335), .B(n_332), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_372), .B(n_349), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_361), .B(n_317), .Y(n_391) );
AO31x2_ASAP7_75t_L g392 ( .A1(n_374), .A2(n_324), .A3(n_347), .B(n_147), .Y(n_392) );
OA21x2_ASAP7_75t_L g393 ( .A1(n_351), .A2(n_324), .B(n_347), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_368), .B(n_327), .Y(n_394) );
INVx11_ASAP7_75t_L g395 ( .A(n_381), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_355), .B(n_327), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_369), .A2(n_315), .B1(n_317), .B2(n_336), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_374), .A2(n_314), .B(n_313), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_363), .B(n_304), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_352), .A2(n_316), .B1(n_342), .B2(n_323), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_365), .A2(n_313), .B(n_319), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_354), .A2(n_323), .B1(n_304), .B2(n_311), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_365), .B(n_326), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_366), .A2(n_277), .B1(n_264), .B2(n_282), .C(n_160), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_353), .A2(n_342), .B1(n_333), .B2(n_334), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_365), .B(n_326), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_370), .A2(n_342), .B1(n_333), .B2(n_334), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_367), .A2(n_303), .B1(n_299), .B2(n_326), .Y(n_408) );
AOI21x1_ASAP7_75t_L g409 ( .A1(n_358), .A2(n_202), .B(n_178), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_367), .A2(n_299), .B1(n_303), .B2(n_328), .Y(n_410) );
AO21x2_ASAP7_75t_L g411 ( .A1(n_398), .A2(n_373), .B(n_376), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_386), .B(n_361), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_384), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_387), .A2(n_356), .B1(n_382), .B2(n_360), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_383), .B(n_367), .Y(n_415) );
OAI211xp5_ASAP7_75t_L g416 ( .A1(n_402), .A2(n_397), .B(n_407), .C(n_405), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_397), .A2(n_357), .B1(n_360), .B2(n_377), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_384), .Y(n_418) );
OAI211xp5_ASAP7_75t_L g419 ( .A1(n_386), .A2(n_377), .B(n_371), .C(n_378), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_384), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_383), .B(n_357), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_388), .Y(n_422) );
OAI31xp33_ASAP7_75t_L g423 ( .A1(n_396), .A2(n_378), .A3(n_359), .B(n_380), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_388), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_392), .Y(n_425) );
AOI33xp33_ASAP7_75t_L g426 ( .A1(n_390), .A2(n_147), .A3(n_137), .B1(n_132), .B2(n_135), .B3(n_359), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_396), .A2(n_362), .B1(n_379), .B2(n_333), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_391), .A2(n_362), .B1(n_376), .B2(n_358), .Y(n_428) );
OAI33xp33_ASAP7_75t_L g429 ( .A1(n_391), .A2(n_137), .A3(n_101), .B1(n_178), .B2(n_183), .B3(n_196), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_390), .B(n_394), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_394), .A2(n_362), .B1(n_376), .B2(n_303), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g432 ( .A1(n_400), .A2(n_151), .B1(n_160), .B2(n_362), .C(n_137), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_400), .A2(n_160), .B1(n_151), .B2(n_201), .C(n_170), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_398), .A2(n_160), .B1(n_151), .B2(n_201), .C(n_170), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_404), .A2(n_303), .B1(n_328), .B2(n_160), .Y(n_435) );
AOI22xp33_ASAP7_75t_SL g436 ( .A1(n_404), .A2(n_350), .B1(n_345), .B2(n_341), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_401), .A2(n_160), .B1(n_170), .B2(n_172), .C(n_204), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_401), .A2(n_172), .B1(n_202), .B2(n_183), .C(n_196), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_399), .B(n_5), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_399), .B(n_6), .Y(n_440) );
BUFx4f_ASAP7_75t_L g441 ( .A(n_406), .Y(n_441) );
AOI211xp5_ASAP7_75t_L g442 ( .A1(n_406), .A2(n_334), .B(n_144), .C(n_341), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_403), .Y(n_443) );
INVx4_ASAP7_75t_L g444 ( .A(n_403), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_393), .B(n_7), .Y(n_445) );
NAND4xp25_ASAP7_75t_L g446 ( .A(n_417), .B(n_395), .C(n_9), .D(n_10), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_443), .Y(n_447) );
INVx3_ASAP7_75t_L g448 ( .A(n_413), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_445), .B(n_392), .Y(n_449) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_444), .A2(n_395), .B1(n_385), .B2(n_393), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_415), .B(n_392), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_415), .B(n_392), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_413), .B(n_392), .Y(n_453) );
NOR2xp33_ASAP7_75t_SL g454 ( .A(n_441), .B(n_385), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_413), .B(n_392), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_418), .B(n_393), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_445), .B(n_389), .Y(n_457) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_442), .B(n_423), .C(n_419), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_422), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_418), .B(n_389), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_412), .B(n_393), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_418), .B(n_393), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_420), .B(n_389), .Y(n_463) );
INVx1_ASAP7_75t_SL g464 ( .A(n_439), .Y(n_464) );
OAI21xp33_ASAP7_75t_L g465 ( .A1(n_421), .A2(n_144), .B(n_408), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_421), .A2(n_389), .B1(n_408), .B2(n_410), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_430), .B(n_8), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_420), .B(n_410), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_420), .B(n_10), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_422), .Y(n_470) );
INVxp67_ASAP7_75t_SL g471 ( .A(n_441), .Y(n_471) );
OAI31xp33_ASAP7_75t_SL g472 ( .A1(n_416), .A2(n_11), .A3(n_14), .B(n_16), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_424), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_424), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_444), .B(n_11), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_444), .B(n_17), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_439), .B(n_17), .Y(n_477) );
OAI211xp5_ASAP7_75t_SL g478 ( .A1(n_423), .A2(n_345), .B(n_18), .C(n_193), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_425), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_425), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_425), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_411), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_444), .B(n_18), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_441), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_440), .B(n_409), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_428), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_411), .Y(n_487) );
OAI21xp33_ASAP7_75t_SL g488 ( .A1(n_426), .A2(n_345), .B(n_20), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_411), .B(n_19), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_428), .B(n_23), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_435), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_414), .B(n_193), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_442), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_427), .B(n_24), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_436), .B(n_350), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_479), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_447), .B(n_431), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_451), .B(n_433), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_479), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_459), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_451), .B(n_432), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_464), .B(n_435), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_475), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_473), .B(n_429), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_459), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_470), .B(n_437), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_452), .B(n_434), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_448), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_473), .B(n_193), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_484), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_470), .B(n_193), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_480), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_452), .B(n_193), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_449), .B(n_26), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_474), .B(n_438), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_474), .B(n_29), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_457), .B(n_39), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_480), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_481), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_469), .B(n_46), .Y(n_520) );
INVxp67_ASAP7_75t_SL g521 ( .A(n_448), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_481), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_475), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_448), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_457), .B(n_48), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_476), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_446), .A2(n_328), .B1(n_350), .B2(n_229), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_457), .B(n_50), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_446), .A2(n_328), .B1(n_350), .B2(n_229), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g530 ( .A1(n_472), .A2(n_229), .B1(n_214), .B2(n_194), .C(n_190), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_457), .B(n_51), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_469), .B(n_52), .Y(n_532) );
OAI211xp5_ASAP7_75t_L g533 ( .A1(n_483), .A2(n_229), .B(n_214), .C(n_194), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_488), .A2(n_54), .B(n_58), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_483), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_454), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_449), .B(n_60), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_449), .B(n_62), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_449), .B(n_68), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_456), .B(n_69), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_471), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_467), .B(n_70), .Y(n_542) );
OA211x2_ASAP7_75t_L g543 ( .A1(n_465), .A2(n_71), .B(n_74), .C(n_75), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_460), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_456), .B(n_77), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_462), .B(n_190), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_493), .Y(n_547) );
BUFx2_ASAP7_75t_L g548 ( .A(n_468), .Y(n_548) );
INVx2_ASAP7_75t_SL g549 ( .A(n_484), .Y(n_549) );
AOI211x1_ASAP7_75t_SL g550 ( .A1(n_478), .A2(n_190), .B(n_194), .C(n_214), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_461), .B(n_190), .Y(n_551) );
INVx2_ASAP7_75t_SL g552 ( .A(n_485), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_552), .B(n_463), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_547), .B(n_463), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_513), .B(n_485), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_503), .Y(n_556) );
OAI32xp33_ASAP7_75t_L g557 ( .A1(n_535), .A2(n_458), .A3(n_488), .B1(n_493), .B2(n_465), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_496), .Y(n_558) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_521), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_523), .B(n_458), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_527), .A2(n_450), .B1(n_494), .B2(n_477), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_552), .B(n_460), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_513), .Y(n_563) );
XNOR2x1_ASAP7_75t_L g564 ( .A(n_510), .B(n_494), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_548), .B(n_460), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_500), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_496), .Y(n_567) );
INVxp67_ASAP7_75t_L g568 ( .A(n_541), .Y(n_568) );
AO211x2_ASAP7_75t_L g569 ( .A1(n_534), .A2(n_450), .B(n_486), .C(n_492), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_538), .B(n_462), .Y(n_570) );
A2O1A1Ixp33_ASAP7_75t_L g571 ( .A1(n_529), .A2(n_490), .B(n_495), .C(n_489), .Y(n_571) );
AND3x2_ASAP7_75t_L g572 ( .A(n_538), .B(n_490), .C(n_489), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_539), .B(n_455), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_526), .A2(n_466), .B1(n_489), .B2(n_460), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_539), .B(n_455), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_509), .Y(n_576) );
OAI211xp5_ASAP7_75t_SL g577 ( .A1(n_530), .A2(n_486), .B(n_487), .C(n_482), .Y(n_577) );
NAND2xp33_ASAP7_75t_L g578 ( .A(n_510), .B(n_468), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_505), .B(n_453), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_499), .B(n_453), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_512), .B(n_487), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_498), .B(n_489), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_512), .Y(n_583) );
BUFx2_ASAP7_75t_L g584 ( .A(n_549), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_498), .B(n_482), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_501), .B(n_491), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_509), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_518), .Y(n_588) );
NOR2x1_ASAP7_75t_L g589 ( .A(n_533), .B(n_491), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_517), .B(n_190), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_517), .B(n_194), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_536), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_519), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_519), .Y(n_594) );
INVxp67_ASAP7_75t_L g595 ( .A(n_497), .Y(n_595) );
NOR2xp33_ASAP7_75t_SL g596 ( .A(n_549), .B(n_266), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_501), .B(n_194), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_525), .B(n_214), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_544), .B(n_214), .Y(n_599) );
AOI211x1_ASAP7_75t_L g600 ( .A1(n_557), .A2(n_525), .B(n_528), .C(n_531), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_567), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_567), .B(n_522), .Y(n_602) );
AO211x2_ASAP7_75t_L g603 ( .A1(n_569), .A2(n_502), .B(n_532), .C(n_520), .Y(n_603) );
INVx3_ASAP7_75t_L g604 ( .A(n_565), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_566), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_585), .B(n_507), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_586), .B(n_507), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_568), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_580), .B(n_595), .Y(n_609) );
INVxp67_ASAP7_75t_L g610 ( .A(n_560), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_560), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_554), .B(n_504), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_583), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_588), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_593), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_555), .B(n_528), .Y(n_616) );
AOI221xp5_ASAP7_75t_SL g617 ( .A1(n_592), .A2(n_531), .B1(n_542), .B2(n_540), .C(n_545), .Y(n_617) );
OAI21xp5_ASAP7_75t_SL g618 ( .A1(n_572), .A2(n_550), .B(n_514), .Y(n_618) );
NAND2xp67_ASAP7_75t_L g619 ( .A(n_562), .B(n_545), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_558), .B(n_504), .Y(n_620) );
NOR2x1_ASAP7_75t_L g621 ( .A(n_571), .B(n_514), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_594), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_553), .B(n_537), .Y(n_623) );
OA211x2_ASAP7_75t_L g624 ( .A1(n_596), .A2(n_543), .B(n_516), .C(n_506), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_553), .B(n_556), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_564), .B(n_514), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_571), .B(n_537), .Y(n_627) );
XNOR2x1_ASAP7_75t_L g628 ( .A(n_564), .B(n_537), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_584), .B(n_524), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_563), .B(n_511), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_578), .Y(n_631) );
XNOR2x2_ASAP7_75t_L g632 ( .A(n_561), .B(n_511), .Y(n_632) );
XNOR2xp5_ASAP7_75t_L g633 ( .A(n_572), .B(n_540), .Y(n_633) );
OAI211xp5_ASAP7_75t_SL g634 ( .A1(n_578), .A2(n_515), .B(n_551), .C(n_524), .Y(n_634) );
INVxp67_ASAP7_75t_L g635 ( .A(n_597), .Y(n_635) );
OAI21xp5_ASAP7_75t_SL g636 ( .A1(n_574), .A2(n_546), .B(n_508), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_581), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_579), .Y(n_638) );
O2A1O1Ixp33_ASAP7_75t_L g639 ( .A1(n_577), .A2(n_551), .B(n_508), .C(n_546), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g640 ( .A1(n_582), .A2(n_229), .B1(n_576), .B2(n_587), .C(n_559), .Y(n_640) );
OAI22xp33_ASAP7_75t_L g641 ( .A1(n_559), .A2(n_589), .B1(n_569), .B2(n_565), .Y(n_641) );
AOI211xp5_ASAP7_75t_SL g642 ( .A1(n_565), .A2(n_590), .B(n_598), .C(n_591), .Y(n_642) );
O2A1O1Ixp33_ASAP7_75t_L g643 ( .A1(n_599), .A2(n_562), .B(n_573), .C(n_575), .Y(n_643) );
OAI211xp5_ASAP7_75t_L g644 ( .A1(n_570), .A2(n_560), .B(n_472), .C(n_571), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_599), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_553), .B(n_562), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_567), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_557), .A2(n_571), .B(n_569), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_553), .B(n_562), .Y(n_649) );
CKINVDCx14_ASAP7_75t_R g650 ( .A(n_584), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_567), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_650), .Y(n_652) );
OAI21xp5_ASAP7_75t_L g653 ( .A1(n_648), .A2(n_621), .B(n_641), .Y(n_653) );
INVxp33_ASAP7_75t_SL g654 ( .A(n_626), .Y(n_654) );
XNOR2xp5_ASAP7_75t_L g655 ( .A(n_628), .B(n_632), .Y(n_655) );
OAI211xp5_ASAP7_75t_SL g656 ( .A1(n_611), .A2(n_610), .B(n_644), .C(n_618), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_650), .B(n_649), .Y(n_657) );
OAI22xp33_ASAP7_75t_SL g658 ( .A1(n_627), .A2(n_631), .B1(n_611), .B2(n_610), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_L g659 ( .A1(n_608), .A2(n_640), .B(n_639), .C(n_634), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_642), .A2(n_633), .B(n_603), .Y(n_660) );
OAI21xp33_ASAP7_75t_L g661 ( .A1(n_636), .A2(n_619), .B(n_612), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_633), .A2(n_602), .B(n_643), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_617), .A2(n_606), .B1(n_638), .B2(n_607), .Y(n_663) );
XNOR2x1_ASAP7_75t_L g664 ( .A(n_609), .B(n_624), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_625), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_652), .Y(n_666) );
NAND4xp25_ASAP7_75t_L g667 ( .A(n_653), .B(n_600), .C(n_630), .D(n_612), .Y(n_667) );
OAI22x1_ASAP7_75t_L g668 ( .A1(n_655), .A2(n_604), .B1(n_651), .B2(n_601), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_656), .A2(n_607), .B1(n_606), .B2(n_605), .C(n_637), .Y(n_669) );
AOI211xp5_ASAP7_75t_L g670 ( .A1(n_658), .A2(n_620), .B(n_635), .C(n_647), .Y(n_670) );
OAI221xp5_ASAP7_75t_L g671 ( .A1(n_660), .A2(n_604), .B1(n_620), .B2(n_602), .C(n_645), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_662), .A2(n_623), .B1(n_616), .B2(n_629), .Y(n_672) );
AOI211xp5_ASAP7_75t_L g673 ( .A1(n_662), .A2(n_615), .B(n_613), .C(n_614), .Y(n_673) );
INVxp67_ASAP7_75t_L g674 ( .A(n_666), .Y(n_674) );
OAI211xp5_ASAP7_75t_L g675 ( .A1(n_673), .A2(n_659), .B(n_663), .C(n_661), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_670), .B(n_654), .Y(n_676) );
NOR3xp33_ASAP7_75t_L g677 ( .A(n_671), .B(n_657), .C(n_664), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_674), .Y(n_678) );
OAI322xp33_ASAP7_75t_L g679 ( .A1(n_676), .A2(n_668), .A3(n_665), .B1(n_667), .B2(n_669), .C1(n_672), .C2(n_622), .Y(n_679) );
NAND3x1_ASAP7_75t_L g680 ( .A(n_677), .B(n_649), .C(n_646), .Y(n_680) );
INVx3_ASAP7_75t_L g681 ( .A(n_678), .Y(n_681) );
OR3x1_ASAP7_75t_L g682 ( .A(n_680), .B(n_679), .C(n_675), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_681), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_683), .Y(n_684) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_684), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_685), .A2(n_681), .B(n_682), .Y(n_686) );
endmodule