module fake_jpeg_24318_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_1),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_31),
.B1(n_19),
.B2(n_32),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_50),
.B1(n_38),
.B2(n_37),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_31),
.B1(n_19),
.B2(n_23),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_48),
.B(n_27),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_23),
.C(n_31),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_22),
.B1(n_23),
.B2(n_31),
.Y(n_50)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_26),
.B1(n_21),
.B2(n_30),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_58),
.B1(n_27),
.B2(n_35),
.Y(n_74)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_65),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_16),
.B1(n_27),
.B2(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_16),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_67),
.B(n_68),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_21),
.C(n_26),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_38),
.B1(n_37),
.B2(n_21),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_70),
.B(n_88),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_71),
.B(n_73),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_77),
.B1(n_89),
.B2(n_99),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_12),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_75),
.B(n_86),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_44),
.B1(n_22),
.B2(n_40),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_79),
.A2(n_108),
.B(n_49),
.Y(n_124)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_80),
.A2(n_85),
.B1(n_102),
.B2(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_26),
.Y(n_81)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_1),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_61),
.B(n_29),
.C(n_34),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_18),
.Y(n_87)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_48),
.A2(n_46),
.B1(n_55),
.B2(n_59),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_90),
.B(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_18),
.Y(n_91)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_18),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_17),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_44),
.B(n_41),
.C(n_40),
.Y(n_94)
);

FAx1_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_56),
.CI(n_53),
.CON(n_109),
.SN(n_109)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_17),
.Y(n_96)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_41),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_106),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_44),
.B1(n_41),
.B2(n_40),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_20),
.B1(n_35),
.B2(n_25),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_104),
.Y(n_113)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_53),
.A2(n_44),
.B1(n_22),
.B2(n_40),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_49),
.A2(n_35),
.B1(n_20),
.B2(n_17),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_109),
.A2(n_78),
.B(n_95),
.C(n_100),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_112),
.A2(n_124),
.B(n_94),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_114),
.B(n_126),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_30),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_SL g162 ( 
.A(n_115),
.B(n_134),
.C(n_12),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_56),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_130),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_93),
.B(n_25),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_12),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_67),
.B(n_53),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_138),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_78),
.B(n_25),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_141),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_142),
.A2(n_149),
.B(n_150),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_89),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_144),
.C(n_157),
.Y(n_185)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_82),
.B(n_94),
.C(n_74),
.D(n_77),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_73),
.B(n_86),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_162),
.B(n_115),
.Y(n_190)
);

AOI22x1_ASAP7_75t_L g146 ( 
.A1(n_109),
.A2(n_99),
.B1(n_75),
.B2(n_103),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_117),
.B1(n_110),
.B2(n_133),
.Y(n_175)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_95),
.B(n_105),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_151),
.B(n_155),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_112),
.A2(n_83),
.B(n_90),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_152),
.A2(n_158),
.B(n_149),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_136),
.A2(n_80),
.B1(n_85),
.B2(n_102),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_154),
.A2(n_163),
.B1(n_167),
.B2(n_131),
.Y(n_174)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_125),
.C(n_128),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_111),
.A2(n_88),
.B1(n_83),
.B2(n_106),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_156),
.A2(n_125),
.B1(n_122),
.B2(n_127),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_107),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_69),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_41),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_121),
.Y(n_171)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_28),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_160),
.B(n_115),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_110),
.B(n_92),
.C(n_97),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_113),
.C(n_131),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_30),
.B1(n_28),
.B2(n_13),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_166),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_138),
.B(n_28),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_168),
.B(n_170),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_SL g169 ( 
.A1(n_109),
.A2(n_24),
.B(n_34),
.Y(n_169)
);

XNOR2x1_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_109),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_123),
.B(n_11),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_197),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_172),
.A2(n_120),
.B1(n_164),
.B2(n_166),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_134),
.B(n_126),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_173),
.A2(n_188),
.B(n_200),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_174),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_179),
.B1(n_151),
.B2(n_34),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_176),
.Y(n_216)
);

OA21x2_ASAP7_75t_L g177 ( 
.A1(n_146),
.A2(n_133),
.B(n_134),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_177),
.A2(n_190),
.B(n_202),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_126),
.Y(n_178)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_119),
.B1(n_117),
.B2(n_121),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_158),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_180),
.B(n_192),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_127),
.B1(n_113),
.B2(n_128),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_184),
.A2(n_186),
.B1(n_203),
.B2(n_24),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_130),
.Y(n_187)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_150),
.C(n_143),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_161),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_193),
.Y(n_231)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_195),
.Y(n_230)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_198),
.Y(n_205)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_144),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_160),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_201),
.A2(n_1),
.B(n_2),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_150),
.A2(n_120),
.B(n_29),
.Y(n_202)
);

AO22x1_ASAP7_75t_SL g203 ( 
.A1(n_150),
.A2(n_92),
.B1(n_84),
.B2(n_104),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_214),
.C(n_215),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_165),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_210),
.Y(n_239)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_223),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_186),
.B1(n_189),
.B2(n_200),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_141),
.C(n_129),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_24),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_129),
.C(n_34),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_222),
.C(n_228),
.Y(n_235)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_221),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_24),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_129),
.C(n_29),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_172),
.B(n_182),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_180),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_225),
.Y(n_256)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_184),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_29),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_229),
.A2(n_188),
.B(n_175),
.Y(n_237)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_249),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_225),
.A2(n_195),
.B1(n_197),
.B2(n_203),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_252),
.B1(n_205),
.B2(n_221),
.Y(n_260)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_187),
.C(n_202),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_241),
.C(n_217),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_206),
.C(n_215),
.Y(n_241)
);

XNOR2x1_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_173),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_242),
.B(n_231),
.Y(n_271)
);

AO21x1_ASAP7_75t_L g243 ( 
.A1(n_216),
.A2(n_190),
.B(n_177),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_210),
.B(n_201),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_177),
.Y(n_244)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_244),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_212),
.A2(n_177),
.B1(n_173),
.B2(n_176),
.Y(n_246)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_246),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_213),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_248),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_230),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_208),
.B(n_199),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_255),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_181),
.Y(n_251)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_205),
.A2(n_227),
.B1(n_204),
.B2(n_224),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

AO221x1_ASAP7_75t_L g269 ( 
.A1(n_253),
.A2(n_219),
.B1(n_218),
.B2(n_228),
.C(n_211),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_208),
.B(n_178),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_261),
.Y(n_282)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_242),
.B(n_207),
.CI(n_171),
.CON(n_258),
.SN(n_258)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_264),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_260),
.A2(n_238),
.B1(n_254),
.B2(n_220),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_232),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_204),
.C(n_207),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_239),
.B(n_209),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_274),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_232),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_271),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_272),
.B(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_181),
.C(n_196),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_196),
.C(n_193),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_235),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_259),
.A2(n_245),
.B(n_239),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_278),
.A2(n_280),
.B(n_281),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_268),
.A2(n_248),
.B1(n_234),
.B2(n_256),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_288),
.B1(n_291),
.B2(n_292),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_262),
.A2(n_237),
.B(n_243),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_L g285 ( 
.A1(n_270),
.A2(n_256),
.B(n_247),
.Y(n_285)
);

AO21x1_ASAP7_75t_L g307 ( 
.A1(n_285),
.A2(n_13),
.B(n_11),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_255),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_293),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_267),
.A2(n_236),
.B1(n_253),
.B2(n_252),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_289),
.B(n_263),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_273),
.B1(n_277),
.B2(n_264),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_274),
.A2(n_260),
.B1(n_246),
.B2(n_257),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_250),
.Y(n_293)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_294),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_263),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_295),
.B(n_302),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_272),
.Y(n_297)
);

AOI32xp33_ASAP7_75t_L g315 ( 
.A1(n_297),
.A2(n_293),
.A3(n_10),
.B1(n_6),
.B2(n_7),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_282),
.C(n_283),
.Y(n_311)
);

NOR4xp25_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_271),
.C(n_275),
.D(n_258),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_10),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_254),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_304),
.B(n_306),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_258),
.B(n_15),
.C(n_14),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_305),
.A2(n_308),
.B(n_14),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_15),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_307),
.B(n_13),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_284),
.A2(n_3),
.B(n_4),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_303),
.A2(n_292),
.B(n_282),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_303),
.B(n_309),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_311),
.B(n_299),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_307),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_283),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_313),
.B(n_314),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_305),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_316),
.B(n_317),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_10),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_322),
.Y(n_329)
);

AOI322xp5_ASAP7_75t_L g327 ( 
.A1(n_323),
.A2(n_324),
.A3(n_326),
.B1(n_318),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_327)
);

MAJx2_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_295),
.C(n_300),
.Y(n_325)
);

MAJx2_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_8),
.C(n_5),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_318),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

AOI322xp5_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_4),
.A3(n_5),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_325),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_4),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_330),
.B(n_331),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_332),
.A2(n_329),
.B(n_7),
.Y(n_334)
);

AO21x1_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_333),
.B(n_8),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_335),
.Y(n_336)
);


endmodule