module real_aes_16730_n_329 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_329);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_329;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_1328;
wire n_571;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1632;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1638;
wire n_1072;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_1672;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1595;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_1352;
wire n_729;
wire n_394;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g1159 ( .A(n_0), .Y(n_1159) );
AO22x1_ASAP7_75t_L g1183 ( .A1(n_0), .A2(n_216), .B1(n_450), .B2(n_1184), .Y(n_1183) );
AND2x2_ASAP7_75t_L g420 ( .A(n_1), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g445 ( .A(n_1), .Y(n_445) );
AND2x2_ASAP7_75t_L g456 ( .A(n_1), .B(n_238), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_1), .B(n_444), .Y(n_889) );
INVx1_ASAP7_75t_L g1168 ( .A(n_2), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_2), .A2(n_112), .B1(n_455), .B2(n_622), .Y(n_1182) );
AOI22xp33_ASAP7_75t_SL g520 ( .A1(n_3), .A2(n_293), .B1(n_370), .B2(n_498), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g547 ( .A1(n_3), .A2(n_5), .B1(n_548), .B2(n_550), .C(n_553), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g1269 ( .A1(n_4), .A2(n_45), .B1(n_613), .B2(n_914), .Y(n_1269) );
INVxp67_ASAP7_75t_SL g1295 ( .A(n_4), .Y(n_1295) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_5), .A2(n_9), .B1(n_366), .B2(n_384), .Y(n_530) );
AOI22xp33_ASAP7_75t_SL g363 ( .A1(n_6), .A2(n_290), .B1(n_364), .B2(n_370), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_6), .A2(n_244), .B1(n_434), .B2(n_438), .C(n_442), .Y(n_433) );
INVx1_ASAP7_75t_L g1074 ( .A(n_7), .Y(n_1074) );
CKINVDCx5p33_ASAP7_75t_R g1303 ( .A(n_8), .Y(n_1303) );
A2O1A1Ixp33_ASAP7_75t_L g565 ( .A1(n_9), .A2(n_566), .B(n_570), .C(n_579), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g1141 ( .A1(n_10), .A2(n_201), .B1(n_398), .B2(n_657), .Y(n_1141) );
INVx1_ASAP7_75t_L g821 ( .A(n_11), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g1440 ( .A1(n_11), .A2(n_195), .B1(n_1414), .B2(n_1428), .Y(n_1440) );
AOI22xp33_ASAP7_75t_SL g1356 ( .A1(n_12), .A2(n_208), .B1(n_382), .B2(n_604), .Y(n_1356) );
INVxp67_ASAP7_75t_SL g1377 ( .A(n_12), .Y(n_1377) );
AOI221xp5_ASAP7_75t_L g833 ( .A1(n_13), .A2(n_283), .B1(n_704), .B2(n_834), .C(n_835), .Y(n_833) );
AOI22xp33_ASAP7_75t_SL g853 ( .A1(n_13), .A2(n_302), .B1(n_343), .B2(n_387), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_14), .A2(n_268), .B1(n_608), .B2(n_612), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_14), .A2(n_80), .B1(n_621), .B2(n_622), .C(n_623), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_15), .A2(n_304), .B1(n_555), .B2(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g752 ( .A(n_15), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g1432 ( .A1(n_16), .A2(n_89), .B1(n_1414), .B2(n_1416), .Y(n_1432) );
AOI22xp33_ASAP7_75t_L g1529 ( .A1(n_17), .A2(n_312), .B1(n_1406), .B2(n_1411), .Y(n_1529) );
INVx2_ASAP7_75t_L g360 ( .A(n_18), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_19), .A2(n_108), .B1(n_1314), .B2(n_1316), .Y(n_1313) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_19), .A2(n_152), .B1(n_463), .B2(n_839), .Y(n_1329) );
INVx1_ASAP7_75t_L g773 ( .A(n_20), .Y(n_773) );
OAI222xp33_ASAP7_75t_L g803 ( .A1(n_20), .A2(n_155), .B1(n_634), .B2(n_655), .C1(n_804), .C2(n_809), .Y(n_803) );
INVx1_ASAP7_75t_L g1120 ( .A(n_21), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_22), .A2(n_212), .B1(n_387), .B2(n_606), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_22), .A2(n_126), .B1(n_625), .B2(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g1659 ( .A(n_23), .Y(n_1659) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_24), .A2(n_250), .B1(n_447), .B2(n_557), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_24), .A2(n_245), .B1(n_613), .B2(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g1118 ( .A(n_25), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_25), .A2(n_65), .B1(n_1133), .B2(n_1134), .Y(n_1132) );
AOI22xp5_ASAP7_75t_L g1437 ( .A1(n_26), .A2(n_204), .B1(n_1406), .B2(n_1411), .Y(n_1437) );
OAI22xp33_ASAP7_75t_L g1324 ( .A1(n_27), .A2(n_193), .B1(n_538), .B2(n_1023), .Y(n_1324) );
INVx1_ASAP7_75t_L g1331 ( .A(n_27), .Y(n_1331) );
AOI22xp33_ASAP7_75t_SL g1320 ( .A1(n_28), .A2(n_83), .B1(n_384), .B2(n_612), .Y(n_1320) );
AOI22xp33_ASAP7_75t_SL g1337 ( .A1(n_28), .A2(n_226), .B1(n_626), .B2(n_627), .Y(n_1337) );
OAI22xp5_ASAP7_75t_L g1027 ( .A1(n_29), .A2(n_284), .B1(n_484), .B2(n_672), .Y(n_1027) );
CKINVDCx5p33_ASAP7_75t_R g660 ( .A(n_30), .Y(n_660) );
HB1xp67_ASAP7_75t_L g1391 ( .A(n_31), .Y(n_1391) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_31), .B(n_1389), .Y(n_1407) );
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_32), .A2(n_175), .B1(n_1414), .B2(n_1528), .Y(n_1527) );
OAI22xp5_ASAP7_75t_SL g1630 ( .A1(n_33), .A2(n_269), .B1(n_1631), .B2(n_1632), .Y(n_1630) );
INVxp67_ASAP7_75t_SL g1662 ( .A(n_33), .Y(n_1662) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_34), .A2(n_205), .B1(n_387), .B2(n_1017), .Y(n_1019) );
AOI221xp5_ASAP7_75t_L g1046 ( .A1(n_34), .A2(n_298), .B1(n_471), .B2(n_1047), .C(n_1049), .Y(n_1046) );
CKINVDCx5p33_ASAP7_75t_R g1342 ( .A(n_35), .Y(n_1342) );
INVxp67_ASAP7_75t_L g337 ( .A(n_36), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g1446 ( .A1(n_36), .A2(n_190), .B1(n_1414), .B2(n_1416), .Y(n_1446) );
AOI22xp5_ASAP7_75t_L g842 ( .A1(n_37), .A2(n_302), .B1(n_447), .B2(n_733), .Y(n_842) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_37), .A2(n_283), .B1(n_387), .B2(n_780), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_38), .A2(n_53), .B1(n_350), .B2(n_921), .Y(n_980) );
INVx1_ASAP7_75t_L g990 ( .A(n_38), .Y(n_990) );
INVx1_ASAP7_75t_L g1013 ( .A(n_39), .Y(n_1013) );
OAI221xp5_ASAP7_75t_L g1039 ( .A1(n_39), .A2(n_231), .B1(n_710), .B2(n_1040), .C(n_1041), .Y(n_1039) );
INVx1_ASAP7_75t_L g898 ( .A(n_40), .Y(n_898) );
INVx1_ASAP7_75t_L g800 ( .A(n_41), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g864 ( .A1(n_42), .A2(n_50), .B1(n_865), .B2(n_866), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_42), .A2(n_148), .B1(n_387), .B2(n_920), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_43), .A2(n_88), .B1(n_349), .B2(n_522), .Y(n_521) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_43), .A2(n_183), .B1(n_438), .B2(n_572), .C(n_573), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g969 ( .A1(n_44), .A2(n_319), .B1(n_372), .B2(n_970), .C(n_971), .Y(n_969) );
AOI221xp5_ASAP7_75t_L g988 ( .A1(n_44), .A2(n_105), .B1(n_704), .B2(n_729), .C(n_989), .Y(n_988) );
AOI221xp5_ASAP7_75t_L g1285 ( .A1(n_45), .A2(n_93), .B1(n_548), .B2(n_1131), .C(n_1286), .Y(n_1285) );
AOI22xp33_ASAP7_75t_L g1354 ( .A1(n_46), .A2(n_265), .B1(n_386), .B2(n_1237), .Y(n_1354) );
INVx1_ASAP7_75t_L g1373 ( .A(n_46), .Y(n_1373) );
INVx1_ASAP7_75t_L g736 ( .A(n_47), .Y(n_736) );
OAI21xp5_ASAP7_75t_L g846 ( .A1(n_48), .A2(n_671), .B(n_847), .Y(n_846) );
NAND5xp2_ASAP7_75t_L g1210 ( .A(n_49), .B(n_1211), .C(n_1233), .D(n_1244), .E(n_1249), .Y(n_1210) );
INVx1_ASAP7_75t_L g1257 ( .A(n_49), .Y(n_1257) );
AOI22xp33_ASAP7_75t_SL g910 ( .A1(n_50), .A2(n_158), .B1(n_911), .B2(n_912), .Y(n_910) );
INVx1_ASAP7_75t_L g735 ( .A(n_51), .Y(n_735) );
INVx1_ASAP7_75t_L g799 ( .A(n_52), .Y(n_799) );
INVx1_ASAP7_75t_L g985 ( .A(n_53), .Y(n_985) );
INVxp67_ASAP7_75t_L g1301 ( .A(n_54), .Y(n_1301) );
AOI22xp5_ASAP7_75t_L g1422 ( .A1(n_54), .A2(n_150), .B1(n_1414), .B2(n_1416), .Y(n_1422) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_55), .Y(n_426) );
INVx1_ASAP7_75t_L g1350 ( .A(n_56), .Y(n_1350) );
INVx1_ASAP7_75t_L g597 ( .A(n_57), .Y(n_597) );
OAI222xp33_ASAP7_75t_L g633 ( .A1(n_57), .A2(n_327), .B1(n_634), .B2(n_635), .C1(n_646), .C2(n_654), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_58), .A2(n_246), .B1(n_1271), .B2(n_1273), .Y(n_1270) );
AOI22xp33_ASAP7_75t_L g1287 ( .A1(n_58), .A2(n_128), .B1(n_447), .B2(n_556), .Y(n_1287) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_59), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g1216 ( .A1(n_60), .A2(n_156), .B1(n_455), .B2(n_622), .C(n_835), .Y(n_1216) );
AOI22xp33_ASAP7_75t_L g1238 ( .A1(n_60), .A2(n_223), .B1(n_387), .B2(n_1239), .Y(n_1238) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_61), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_62), .A2(n_223), .B1(n_733), .B2(n_1184), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_62), .A2(n_156), .B1(n_387), .B2(n_1237), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_63), .A2(n_146), .B1(n_342), .B2(n_386), .Y(n_385) );
AOI21xp33_ASAP7_75t_L g468 ( .A1(n_63), .A2(n_469), .B(n_471), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_64), .A2(n_823), .B1(n_824), .B2(n_858), .Y(n_822) );
INVxp67_ASAP7_75t_SL g858 ( .A(n_64), .Y(n_858) );
INVx1_ASAP7_75t_L g1107 ( .A(n_65), .Y(n_1107) );
INVx1_ASAP7_75t_L g517 ( .A(n_66), .Y(n_517) );
AOI221xp5_ASAP7_75t_L g867 ( .A1(n_67), .A2(n_306), .B1(n_868), .B2(n_869), .C(n_871), .Y(n_867) );
AOI221xp5_ASAP7_75t_L g915 ( .A1(n_67), .A2(n_271), .B1(n_758), .B2(n_916), .C(n_918), .Y(n_915) );
AOI22xp33_ASAP7_75t_SL g1352 ( .A1(n_68), .A2(n_160), .B1(n_364), .B2(n_758), .Y(n_1352) );
INVxp67_ASAP7_75t_SL g1376 ( .A(n_68), .Y(n_1376) );
OAI211xp5_ASAP7_75t_SL g960 ( .A1(n_69), .A2(n_930), .B(n_937), .C(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g995 ( .A(n_69), .Y(n_995) );
INVx1_ASAP7_75t_L g831 ( .A(n_70), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_71), .Y(n_396) );
OAI21xp5_ASAP7_75t_SL g483 ( .A1(n_72), .A2(n_484), .B(n_496), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g1224 ( .A(n_73), .Y(n_1224) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_74), .A2(n_220), .B1(n_604), .B2(n_914), .Y(n_1066) );
AOI22xp33_ASAP7_75t_SL g1091 ( .A1(n_74), .A2(n_267), .B1(n_466), .B2(n_555), .Y(n_1091) );
INVxp67_ASAP7_75t_SL g903 ( .A(n_75), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_75), .A2(n_313), .B1(n_923), .B2(n_926), .Y(n_922) );
AOI22xp33_ASAP7_75t_SL g1020 ( .A1(n_76), .A2(n_321), .B1(n_613), .B2(n_1021), .Y(n_1020) );
AOI221xp5_ASAP7_75t_L g1033 ( .A1(n_76), .A2(n_132), .B1(n_442), .B2(n_459), .C(n_1034), .Y(n_1033) );
AOI22xp33_ASAP7_75t_SL g381 ( .A1(n_77), .A2(n_244), .B1(n_366), .B2(n_382), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_77), .A2(n_290), .B1(n_463), .B2(n_466), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g1275 ( .A1(n_78), .A2(n_93), .B1(n_914), .B2(n_1276), .Y(n_1275) );
INVxp67_ASAP7_75t_SL g1296 ( .A(n_78), .Y(n_1296) );
INVx1_ASAP7_75t_L g832 ( .A(n_79), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_80), .A2(n_119), .B1(n_606), .B2(n_608), .Y(n_605) );
AOI22xp33_ASAP7_75t_SL g1065 ( .A1(n_81), .A2(n_211), .B1(n_912), .B2(n_1063), .Y(n_1065) );
INVx1_ASAP7_75t_L g1086 ( .A(n_81), .Y(n_1086) );
AOI22xp33_ASAP7_75t_SL g1635 ( .A1(n_82), .A2(n_147), .B1(n_450), .B2(n_797), .Y(n_1635) );
INVxp67_ASAP7_75t_SL g1655 ( .A(n_82), .Y(n_1655) );
AOI221xp5_ASAP7_75t_L g1328 ( .A1(n_83), .A2(n_295), .B1(n_553), .B2(n_622), .C(n_1049), .Y(n_1328) );
INVx1_ASAP7_75t_L g1379 ( .A(n_84), .Y(n_1379) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_85), .A2(n_256), .B1(n_613), .B2(n_686), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_85), .A2(n_254), .B1(n_549), .B2(n_553), .C(n_704), .Y(n_703) );
OAI21xp33_ASAP7_75t_L g656 ( .A1(n_86), .A2(n_657), .B(n_658), .Y(n_656) );
INVx1_ASAP7_75t_L g684 ( .A(n_87), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_87), .A2(n_275), .B1(n_463), .B2(n_557), .Y(n_705) );
AOI22xp33_ASAP7_75t_SL g554 ( .A1(n_88), .A2(n_123), .B1(n_555), .B2(n_556), .Y(n_554) );
AOI22xp33_ASAP7_75t_SL g785 ( .A1(n_90), .A2(n_301), .B1(n_613), .B2(n_686), .Y(n_785) );
INVxp67_ASAP7_75t_SL g792 ( .A(n_90), .Y(n_792) );
INVx1_ASAP7_75t_L g1117 ( .A(n_91), .Y(n_1117) );
AOI221xp5_ASAP7_75t_L g1127 ( .A1(n_91), .A2(n_213), .B1(n_434), .B2(n_471), .C(n_621), .Y(n_1127) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_92), .Y(n_427) );
XNOR2xp5_ASAP7_75t_L g723 ( .A(n_94), .B(n_724), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g1405 ( .A1(n_95), .A2(n_202), .B1(n_1406), .B2(n_1411), .Y(n_1405) );
OAI211xp5_ASAP7_75t_L g1220 ( .A1(n_96), .A2(n_1087), .B(n_1221), .C(n_1223), .Y(n_1220) );
INVx1_ASAP7_75t_L g1253 ( .A(n_96), .Y(n_1253) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_97), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_97), .A2(n_109), .B1(n_475), .B2(n_478), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g1640 ( .A1(n_98), .A2(n_222), .B1(n_450), .B2(n_465), .Y(n_1640) );
AOI22xp33_ASAP7_75t_L g1652 ( .A1(n_98), .A2(n_240), .B1(n_366), .B2(n_914), .Y(n_1652) );
AOI21xp33_ASAP7_75t_L g742 ( .A1(n_99), .A2(n_704), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g751 ( .A(n_99), .Y(n_751) );
INVx1_ASAP7_75t_L g669 ( .A(n_100), .Y(n_669) );
INVx1_ASAP7_75t_L g1623 ( .A(n_101), .Y(n_1623) );
INVx1_ASAP7_75t_L g1389 ( .A(n_102), .Y(n_1389) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_103), .A2(n_239), .B1(n_553), .B2(n_729), .C(n_730), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_103), .A2(n_162), .B1(n_371), .B2(n_613), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_104), .A2(n_168), .B1(n_784), .B2(n_1237), .Y(n_1353) );
INVx1_ASAP7_75t_L g1374 ( .A(n_104), .Y(n_1374) );
INVx1_ASAP7_75t_L g976 ( .A(n_105), .Y(n_976) );
OAI22xp33_ASAP7_75t_L g1102 ( .A1(n_106), .A2(n_278), .B1(n_532), .B2(n_1103), .Y(n_1102) );
INVx1_ASAP7_75t_L g1137 ( .A(n_106), .Y(n_1137) );
OAI222xp33_ASAP7_75t_L g1173 ( .A1(n_107), .A2(n_305), .B1(n_933), .B2(n_935), .C1(n_1174), .C2(n_1176), .Y(n_1173) );
INVx1_ASAP7_75t_L g1187 ( .A(n_107), .Y(n_1187) );
AOI21xp33_ASAP7_75t_L g1336 ( .A1(n_108), .A2(n_436), .B(n_835), .Y(n_1336) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_109), .Y(n_405) );
INVx1_ASAP7_75t_L g1267 ( .A(n_110), .Y(n_1267) );
OAI221xp5_ASAP7_75t_L g1291 ( .A1(n_110), .A2(n_111), .B1(n_710), .B2(n_1040), .C(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1266 ( .A(n_111), .Y(n_1266) );
INVx1_ASAP7_75t_L g1164 ( .A(n_112), .Y(n_1164) );
OAI211xp5_ASAP7_75t_L g1625 ( .A1(n_113), .A2(n_805), .B(n_1626), .C(n_1627), .Y(n_1625) );
INVxp33_ASAP7_75t_SL g1644 ( .A(n_113), .Y(n_1644) );
CKINVDCx5p33_ASAP7_75t_R g692 ( .A(n_114), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g940 ( .A1(n_115), .A2(n_153), .B1(n_941), .B2(n_944), .Y(n_940) );
INVxp67_ASAP7_75t_SL g947 ( .A(n_115), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g1426 ( .A1(n_116), .A2(n_297), .B1(n_1406), .B2(n_1411), .Y(n_1426) );
INVx1_ASAP7_75t_L g1109 ( .A(n_117), .Y(n_1109) );
AOI221xp5_ASAP7_75t_L g1130 ( .A1(n_117), .A2(n_262), .B1(n_572), .B2(n_621), .C(n_1131), .Y(n_1130) );
INVx1_ASAP7_75t_L g840 ( .A(n_118), .Y(n_840) );
INVx1_ASAP7_75t_L g644 ( .A(n_119), .Y(n_644) );
INVx1_ASAP7_75t_L g679 ( .A(n_120), .Y(n_679) );
AOI21xp33_ASAP7_75t_L g715 ( .A1(n_120), .A2(n_471), .B(n_704), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_121), .A2(n_151), .B1(n_671), .B2(n_672), .Y(n_670) );
OAI211xp5_ASAP7_75t_L g701 ( .A1(n_121), .A2(n_618), .B(n_702), .C(n_706), .Y(n_701) );
INVx1_ASAP7_75t_L g1346 ( .A(n_122), .Y(n_1346) );
OAI222xp33_ASAP7_75t_L g1370 ( .A1(n_122), .A2(n_191), .B1(n_654), .B2(n_1371), .C1(n_1372), .C2(n_1375), .Y(n_1370) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_123), .A2(n_183), .B1(n_349), .B2(n_526), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g1436 ( .A1(n_124), .A2(n_207), .B1(n_1414), .B2(n_1416), .Y(n_1436) );
AOI221xp5_ASAP7_75t_L g841 ( .A1(n_125), .A2(n_245), .B1(n_442), .B2(n_552), .C(n_729), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_125), .A2(n_250), .B1(n_371), .B2(n_613), .Y(n_852) );
AOI22xp33_ASAP7_75t_SL g603 ( .A1(n_126), .A2(n_215), .B1(n_387), .B2(n_604), .Y(n_603) );
OAI22xp33_ASAP7_75t_L g959 ( .A1(n_127), .A2(n_326), .B1(n_941), .B2(n_944), .Y(n_959) );
INVxp33_ASAP7_75t_SL g999 ( .A(n_127), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1274 ( .A1(n_128), .A2(n_159), .B1(n_1271), .B2(n_1273), .Y(n_1274) );
INVx1_ASAP7_75t_L g1056 ( .A(n_129), .Y(n_1056) );
OAI221xp5_ASAP7_75t_L g1084 ( .A1(n_129), .A2(n_130), .B1(n_634), .B2(n_655), .C(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_L g1057 ( .A(n_130), .Y(n_1057) );
CKINVDCx5p33_ASAP7_75t_R g962 ( .A(n_131), .Y(n_962) );
AOI22xp33_ASAP7_75t_SL g1015 ( .A1(n_132), .A2(n_174), .B1(n_613), .B2(n_914), .Y(n_1015) );
AOI22xp5_ASAP7_75t_L g1441 ( .A1(n_133), .A2(n_221), .B1(n_1406), .B2(n_1411), .Y(n_1441) );
INVx1_ASAP7_75t_L g966 ( .A(n_134), .Y(n_966) );
AOI221xp5_ASAP7_75t_L g983 ( .A1(n_134), .A2(n_233), .B1(n_704), .B2(n_729), .C(n_984), .Y(n_983) );
AOI221xp5_ASAP7_75t_L g882 ( .A1(n_135), .A2(n_148), .B1(n_866), .B2(n_883), .C(n_885), .Y(n_882) );
AOI221xp5_ASAP7_75t_L g913 ( .A1(n_135), .A2(n_306), .B1(n_613), .B2(n_788), .C(n_914), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_136), .A2(n_298), .B1(n_781), .B2(n_1017), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_136), .A2(n_205), .B1(n_449), .B2(n_1032), .Y(n_1031) );
OAI22xp33_ASAP7_75t_L g1278 ( .A1(n_137), .A2(n_264), .B1(n_532), .B2(n_538), .Y(n_1278) );
INVx1_ASAP7_75t_L g1290 ( .A(n_137), .Y(n_1290) );
INVx1_ASAP7_75t_L g826 ( .A(n_138), .Y(n_826) );
INVx1_ASAP7_75t_L g1360 ( .A(n_139), .Y(n_1360) );
INVx1_ASAP7_75t_L g1306 ( .A(n_140), .Y(n_1306) );
OAI221xp5_ASAP7_75t_SL g1333 ( .A1(n_140), .A2(n_242), .B1(n_654), .B2(n_710), .C(n_1334), .Y(n_1333) );
CKINVDCx5p33_ASAP7_75t_R g1026 ( .A(n_141), .Y(n_1026) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_142), .A2(n_314), .B1(n_634), .B2(n_655), .C(n_738), .Y(n_737) );
OAI22xp33_ASAP7_75t_L g759 ( .A1(n_142), .A2(n_314), .B1(n_596), .B2(n_698), .Y(n_759) );
INVx1_ASAP7_75t_L g661 ( .A(n_143), .Y(n_661) );
AO22x1_ASAP7_75t_L g341 ( .A1(n_144), .A2(n_181), .B1(n_342), .B2(n_349), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_144), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g1248 ( .A(n_145), .Y(n_1248) );
AOI22xp33_ASAP7_75t_SL g446 ( .A1(n_146), .A2(n_181), .B1(n_447), .B2(n_449), .Y(n_446) );
INVx1_ASAP7_75t_L g1651 ( .A(n_147), .Y(n_1651) );
CKINVDCx5p33_ASAP7_75t_R g1629 ( .A(n_149), .Y(n_1629) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_152), .A2(n_285), .B1(n_1316), .B2(n_1318), .Y(n_1317) );
INVxp67_ASAP7_75t_SL g894 ( .A(n_153), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g1281 ( .A1(n_154), .A2(n_172), .B1(n_484), .B2(n_672), .Y(n_1281) );
OAI211xp5_ASAP7_75t_L g1283 ( .A1(n_154), .A2(n_618), .B(n_1284), .C(n_1288), .Y(n_1283) );
INVx1_ASAP7_75t_L g771 ( .A(n_155), .Y(n_771) );
INVx1_ASAP7_75t_L g1161 ( .A(n_157), .Y(n_1161) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_157), .A2(n_247), .B1(n_733), .B2(n_1184), .Y(n_1195) );
INVx1_ASAP7_75t_L g886 ( .A(n_158), .Y(n_886) );
AOI221xp5_ASAP7_75t_L g1297 ( .A1(n_159), .A2(n_246), .B1(n_471), .B2(n_621), .C(n_1298), .Y(n_1297) );
AOI221xp5_ASAP7_75t_L g1365 ( .A1(n_160), .A2(n_208), .B1(n_623), .B2(n_1366), .C(n_1367), .Y(n_1365) );
CKINVDCx5p33_ASAP7_75t_R g1628 ( .A(n_161), .Y(n_1628) );
AOI22xp33_ASAP7_75t_SL g744 ( .A1(n_162), .A2(n_291), .B1(n_447), .B2(n_450), .Y(n_744) );
OAI211xp5_ASAP7_75t_L g726 ( .A1(n_163), .A2(n_618), .B(n_727), .C(n_734), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_163), .A2(n_308), .B1(n_671), .B2(n_672), .Y(n_762) );
INVx1_ASAP7_75t_L g1638 ( .A(n_164), .Y(n_1638) );
AOI22xp33_ASAP7_75t_SL g1062 ( .A1(n_165), .A2(n_272), .B1(n_912), .B2(n_1063), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_165), .A2(n_211), .B1(n_557), .B2(n_626), .Y(n_1080) );
OAI211xp5_ASAP7_75t_L g1212 ( .A1(n_166), .A2(n_1213), .B(n_1214), .C(n_1219), .Y(n_1212) );
NOR2xp33_ASAP7_75t_L g1232 ( .A(n_166), .B(n_398), .Y(n_1232) );
XNOR2x2_ASAP7_75t_L g1007 ( .A(n_167), .B(n_1008), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1368 ( .A1(n_168), .A2(n_265), .B1(n_1032), .B2(n_1134), .Y(n_1368) );
INVx2_ASAP7_75t_L g1409 ( .A(n_169), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1412 ( .A(n_169), .B(n_1410), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_169), .B(n_276), .Y(n_1417) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_170), .A2(n_318), .B1(n_780), .B2(n_781), .Y(n_779) );
INVx1_ASAP7_75t_L g808 ( .A(n_170), .Y(n_808) );
AOI22xp5_ASAP7_75t_L g1421 ( .A1(n_171), .A2(n_257), .B1(n_1406), .B2(n_1411), .Y(n_1421) );
INVx1_ASAP7_75t_L g708 ( .A(n_173), .Y(n_708) );
INVxp67_ASAP7_75t_SL g1042 ( .A(n_174), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_176), .A2(n_266), .B1(n_398), .B2(n_484), .Y(n_542) );
OAI211xp5_ASAP7_75t_L g544 ( .A1(n_176), .A2(n_545), .B(n_546), .C(n_558), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_177), .Y(n_417) );
XOR2x2_ASAP7_75t_L g1261 ( .A(n_178), .B(n_1262), .Y(n_1261) );
OAI22xp33_ASAP7_75t_L g1022 ( .A1(n_179), .A2(n_249), .B1(n_538), .B2(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g1036 ( .A(n_179), .Y(n_1036) );
INVx1_ASAP7_75t_L g1323 ( .A(n_180), .Y(n_1323) );
AOI22xp5_ASAP7_75t_L g1427 ( .A1(n_182), .A2(n_282), .B1(n_1414), .B2(n_1428), .Y(n_1427) );
INVx1_ASAP7_75t_L g1202 ( .A(n_184), .Y(n_1202) );
INVx1_ASAP7_75t_L g1359 ( .A(n_185), .Y(n_1359) );
AOI22xp33_ASAP7_75t_L g1215 ( .A1(n_186), .A2(n_261), .B1(n_465), .B2(n_733), .Y(n_1215) );
AOI22xp33_ASAP7_75t_SL g1240 ( .A1(n_186), .A2(n_274), .B1(n_613), .B2(n_856), .Y(n_1240) );
AOI22xp33_ASAP7_75t_SL g685 ( .A1(n_187), .A2(n_254), .B1(n_613), .B2(n_686), .Y(n_685) );
AOI22xp33_ASAP7_75t_SL g716 ( .A1(n_187), .A2(n_256), .B1(n_447), .B2(n_466), .Y(n_716) );
INVx1_ASAP7_75t_L g820 ( .A(n_188), .Y(n_820) );
INVx1_ASAP7_75t_L g1113 ( .A(n_189), .Y(n_1113) );
INVx1_ASAP7_75t_L g1347 ( .A(n_191), .Y(n_1347) );
INVx1_ASAP7_75t_L g600 ( .A(n_192), .Y(n_600) );
OAI211xp5_ASAP7_75t_L g617 ( .A1(n_192), .A2(n_618), .B(n_619), .C(n_629), .Y(n_617) );
INVx1_ASAP7_75t_L g1332 ( .A(n_193), .Y(n_1332) );
CKINVDCx5p33_ASAP7_75t_R g1163 ( .A(n_194), .Y(n_1163) );
CKINVDCx5p33_ASAP7_75t_R g739 ( .A(n_196), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g1075 ( .A1(n_197), .A2(n_323), .B1(n_538), .B2(n_1023), .Y(n_1075) );
INVx1_ASAP7_75t_L g1082 ( .A(n_197), .Y(n_1082) );
CKINVDCx5p33_ASAP7_75t_R g1227 ( .A(n_198), .Y(n_1227) );
INVx2_ASAP7_75t_L g358 ( .A(n_199), .Y(n_358) );
INVx1_ASAP7_75t_L g380 ( .A(n_199), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_199), .B(n_360), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_200), .Y(n_630) );
OAI211xp5_ASAP7_75t_L g1128 ( .A1(n_201), .A2(n_618), .B(n_1129), .C(n_1136), .Y(n_1128) );
INVx1_ASAP7_75t_L g1171 ( .A(n_203), .Y(n_1171) );
NAND2xp33_ASAP7_75t_SL g1196 ( .A(n_203), .B(n_455), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_206), .A2(n_292), .B1(n_691), .B2(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g806 ( .A(n_206), .Y(n_806) );
AOI22xp33_ASAP7_75t_SL g777 ( .A1(n_209), .A2(n_235), .B1(n_613), .B2(n_778), .Y(n_777) );
INVxp67_ASAP7_75t_SL g810 ( .A(n_209), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g1431 ( .A1(n_210), .A2(n_289), .B1(n_1406), .B2(n_1411), .Y(n_1431) );
INVx1_ASAP7_75t_L g639 ( .A(n_212), .Y(n_639) );
INVx1_ASAP7_75t_L g1114 ( .A(n_213), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g1230 ( .A1(n_214), .A2(n_280), .B1(n_1221), .B2(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1251 ( .A(n_214), .Y(n_1251) );
INVx1_ASAP7_75t_L g647 ( .A(n_215), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g1172 ( .A1(n_216), .A2(n_788), .B(n_921), .Y(n_1172) );
INVx1_ASAP7_75t_L g1198 ( .A(n_217), .Y(n_1198) );
OAI21xp5_ASAP7_75t_L g814 ( .A1(n_218), .A2(n_671), .B(n_815), .Y(n_814) );
BUFx3_ASAP7_75t_L g348 ( .A(n_219), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g1079 ( .A1(n_220), .A2(n_228), .B1(n_549), .B2(n_553), .C(n_704), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g1656 ( .A1(n_222), .A2(n_258), .B1(n_914), .B2(n_1657), .Y(n_1656) );
CKINVDCx5p33_ASAP7_75t_R g963 ( .A(n_224), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_225), .A2(n_229), .B1(n_596), .B2(n_1101), .Y(n_1100) );
OAI221xp5_ASAP7_75t_L g1125 ( .A1(n_225), .A2(n_229), .B1(n_654), .B2(n_710), .C(n_1126), .Y(n_1125) );
AOI22xp33_ASAP7_75t_SL g1312 ( .A1(n_226), .A2(n_295), .B1(n_382), .B2(n_612), .Y(n_1312) );
INVx1_ASAP7_75t_L g1153 ( .A(n_227), .Y(n_1153) );
NOR2xp33_ASAP7_75t_L g1155 ( .A(n_227), .B(n_941), .Y(n_1155) );
AOI22xp33_ASAP7_75t_SL g1061 ( .A1(n_228), .A2(n_267), .B1(n_364), .B2(n_914), .Y(n_1061) );
AOI21xp33_ASAP7_75t_L g1639 ( .A1(n_230), .A2(n_704), .B(n_835), .Y(n_1639) );
INVx1_ASAP7_75t_L g1649 ( .A(n_230), .Y(n_1649) );
INVx1_ASAP7_75t_L g1012 ( .A(n_231), .Y(n_1012) );
INVx1_ASAP7_75t_L g1097 ( .A(n_232), .Y(n_1097) );
AOI21xp33_ASAP7_75t_L g979 ( .A1(n_233), .A2(n_528), .B(n_918), .Y(n_979) );
AOI22xp5_ASAP7_75t_L g1413 ( .A1(n_234), .A2(n_248), .B1(n_1414), .B2(n_1416), .Y(n_1413) );
XOR2x2_ASAP7_75t_L g1618 ( .A(n_234), .B(n_1619), .Y(n_1618) );
AOI22xp33_ASAP7_75t_L g1666 ( .A1(n_234), .A2(n_1667), .B1(n_1670), .B2(n_1673), .Y(n_1666) );
AOI21xp33_ASAP7_75t_L g794 ( .A1(n_235), .A2(n_442), .B(n_795), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_236), .B(n_1052), .Y(n_1051) );
AOI22xp5_ASAP7_75t_L g1069 ( .A1(n_236), .A2(n_1070), .B1(n_1071), .B2(n_1092), .Y(n_1069) );
INVx1_ASAP7_75t_L g1094 ( .A(n_236), .Y(n_1094) );
OAI22xp33_ASAP7_75t_L g531 ( .A1(n_237), .A2(n_253), .B1(n_532), .B2(n_538), .Y(n_531) );
INVx1_ASAP7_75t_L g559 ( .A(n_237), .Y(n_559) );
INVx1_ASAP7_75t_L g421 ( .A(n_238), .Y(n_421) );
BUFx3_ASAP7_75t_L g444 ( .A(n_238), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_239), .A2(n_291), .B1(n_613), .B2(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g1634 ( .A(n_240), .B(n_704), .Y(n_1634) );
INVxp67_ASAP7_75t_SL g1310 ( .A(n_241), .Y(n_1310) );
OAI211xp5_ASAP7_75t_SL g1326 ( .A1(n_241), .A2(n_545), .B(n_1327), .C(n_1330), .Y(n_1326) );
INVx1_ASAP7_75t_L g1308 ( .A(n_242), .Y(n_1308) );
CKINVDCx5p33_ASAP7_75t_R g968 ( .A(n_243), .Y(n_968) );
INVx1_ASAP7_75t_L g1169 ( .A(n_247), .Y(n_1169) );
INVx1_ASAP7_75t_L g1037 ( .A(n_249), .Y(n_1037) );
CKINVDCx5p33_ASAP7_75t_R g1068 ( .A(n_251), .Y(n_1068) );
INVx1_ASAP7_75t_L g518 ( .A(n_252), .Y(n_518) );
INVx1_ASAP7_75t_L g562 ( .A(n_253), .Y(n_562) );
INVx1_ASAP7_75t_L g707 ( .A(n_255), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g1636 ( .A(n_258), .B(n_1034), .Y(n_1636) );
INVx1_ASAP7_75t_L g950 ( .A(n_259), .Y(n_950) );
XNOR2x2_ASAP7_75t_L g512 ( .A(n_260), .B(n_513), .Y(n_512) );
AOI22xp33_ASAP7_75t_SL g1235 ( .A1(n_261), .A2(n_328), .B1(n_613), .B2(n_686), .Y(n_1235) );
INVx1_ASAP7_75t_L g1121 ( .A(n_262), .Y(n_1121) );
INVx1_ASAP7_75t_L g346 ( .A(n_263), .Y(n_346) );
INVx1_ASAP7_75t_L g354 ( .A(n_263), .Y(n_354) );
INVx1_ASAP7_75t_L g1289 ( .A(n_264), .Y(n_1289) );
INVx1_ASAP7_75t_L g653 ( .A(n_268), .Y(n_653) );
OAI21xp33_ASAP7_75t_L g1642 ( .A1(n_269), .A2(n_1246), .B(n_1643), .Y(n_1642) );
INVx1_ASAP7_75t_L g775 ( .A(n_270), .Y(n_775) );
INVx1_ASAP7_75t_L g887 ( .A(n_271), .Y(n_887) );
AOI21xp33_ASAP7_75t_L g1088 ( .A1(n_272), .A2(n_471), .B(n_1089), .Y(n_1088) );
CKINVDCx5p33_ASAP7_75t_R g1152 ( .A(n_273), .Y(n_1152) );
AOI221xp5_ASAP7_75t_SL g1218 ( .A1(n_274), .A2(n_328), .B1(n_436), .B2(n_442), .C(n_455), .Y(n_1218) );
INVx1_ASAP7_75t_L g695 ( .A(n_275), .Y(n_695) );
INVx1_ASAP7_75t_L g1410 ( .A(n_276), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1415 ( .A(n_276), .B(n_1409), .Y(n_1415) );
INVx1_ASAP7_75t_L g845 ( .A(n_277), .Y(n_845) );
INVx1_ASAP7_75t_L g1138 ( .A(n_278), .Y(n_1138) );
XNOR2xp5_ASAP7_75t_L g1671 ( .A(n_279), .B(n_1672), .Y(n_1671) );
INVx1_ASAP7_75t_L g1243 ( .A(n_280), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1447 ( .A1(n_281), .A2(n_315), .B1(n_1406), .B2(n_1411), .Y(n_1447) );
XNOR2xp5_ASAP7_75t_L g951 ( .A(n_282), .B(n_952), .Y(n_951) );
OAI211xp5_ASAP7_75t_L g1029 ( .A1(n_284), .A2(n_545), .B(n_1030), .C(n_1035), .Y(n_1029) );
INVx1_ASAP7_75t_L g1335 ( .A(n_285), .Y(n_1335) );
INVx1_ASAP7_75t_L g844 ( .A(n_286), .Y(n_844) );
INVxp67_ASAP7_75t_SL g1059 ( .A(n_287), .Y(n_1059) );
OAI211xp5_ASAP7_75t_L g1077 ( .A1(n_287), .A2(n_618), .B(n_1078), .C(n_1081), .Y(n_1077) );
CKINVDCx16_ASAP7_75t_R g1175 ( .A(n_288), .Y(n_1175) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_292), .A2(n_318), .B1(n_557), .B2(n_797), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_293), .B(n_575), .Y(n_574) );
OAI21xp33_ASAP7_75t_L g1357 ( .A1(n_294), .A2(n_484), .B(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g954 ( .A(n_296), .Y(n_954) );
INVx1_ASAP7_75t_L g974 ( .A(n_299), .Y(n_974) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_300), .Y(n_511) );
INVxp67_ASAP7_75t_SL g812 ( .A(n_301), .Y(n_812) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_303), .Y(n_424) );
INVx1_ASAP7_75t_L g756 ( .A(n_304), .Y(n_756) );
NOR2xp33_ASAP7_75t_R g1189 ( .A(n_305), .B(n_1190), .Y(n_1189) );
INVx1_ASAP7_75t_L g1148 ( .A(n_307), .Y(n_1148) );
INVxp67_ASAP7_75t_SL g901 ( .A(n_309), .Y(n_901) );
OAI221xp5_ASAP7_75t_L g932 ( .A1(n_309), .A2(n_311), .B1(n_933), .B2(n_935), .C(n_937), .Y(n_932) );
INVx1_ASAP7_75t_L g761 ( .A(n_310), .Y(n_761) );
OAI221xp5_ASAP7_75t_L g873 ( .A1(n_311), .A2(n_313), .B1(n_874), .B2(n_879), .C(n_880), .Y(n_873) );
INVx2_ASAP7_75t_L g362 ( .A(n_316), .Y(n_362) );
INVx1_ASAP7_75t_L g379 ( .A(n_316), .Y(n_379) );
INVx1_ASAP7_75t_L g403 ( .A(n_316), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g1280 ( .A(n_317), .Y(n_1280) );
INVx1_ASAP7_75t_L g986 ( .A(n_319), .Y(n_986) );
CKINVDCx5p33_ASAP7_75t_R g1140 ( .A(n_320), .Y(n_1140) );
INVxp67_ASAP7_75t_SL g1045 ( .A(n_321), .Y(n_1045) );
OAI22xp33_ASAP7_75t_SL g697 ( .A1(n_322), .A2(n_325), .B1(n_596), .B2(n_698), .Y(n_697) );
OAI221xp5_ASAP7_75t_L g709 ( .A1(n_322), .A2(n_325), .B1(n_655), .B2(n_710), .C(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g1083 ( .A(n_323), .Y(n_1083) );
XNOR2xp5_ASAP7_75t_L g666 ( .A(n_324), .B(n_667), .Y(n_666) );
INVxp67_ASAP7_75t_SL g957 ( .A(n_326), .Y(n_957) );
INVx1_ASAP7_75t_L g594 ( .A(n_327), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_1383), .B(n_1399), .Y(n_329) );
XNOR2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_1001), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
XNOR2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_662), .Y(n_332) );
XNOR2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_590), .Y(n_333) );
OAI22x1_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B1(n_512), .B2(n_589), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
XNOR2x1_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
AND3x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_414), .C(n_502), .Y(n_338) );
NOR2xp33_ASAP7_75t_SL g339 ( .A(n_340), .B(n_388), .Y(n_339) );
OAI21xp5_ASAP7_75t_SL g340 ( .A1(n_341), .A2(n_355), .B(n_373), .Y(n_340) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g501 ( .A(n_343), .B(n_500), .Y(n_501) );
INVx2_ASAP7_75t_SL g750 ( .A(n_343), .Y(n_750) );
INVx2_ASAP7_75t_SL g1116 ( .A(n_343), .Y(n_1116) );
INVx3_ASAP7_75t_L g1272 ( .A(n_343), .Y(n_1272) );
INVx3_ASAP7_75t_L g1319 ( .A(n_343), .Y(n_1319) );
BUFx8_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g524 ( .A(n_344), .Y(n_524) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_344), .Y(n_528) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_344), .Y(n_691) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
INVxp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g369 ( .A(n_346), .Y(n_369) );
AND2x4_ASAP7_75t_L g367 ( .A(n_347), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_348), .Y(n_351) );
AND2x4_ASAP7_75t_L g372 ( .A(n_348), .B(n_353), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_348), .B(n_354), .Y(n_508) );
OR2x2_ASAP7_75t_L g535 ( .A(n_348), .B(n_369), .Y(n_535) );
BUFx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx12f_ASAP7_75t_L g387 ( .A(n_350), .Y(n_387) );
INVx5_ASAP7_75t_L g782 ( .A(n_350), .Y(n_782) );
BUFx2_ASAP7_75t_L g912 ( .A(n_350), .Y(n_912) );
AND2x4_ASAP7_75t_L g945 ( .A(n_350), .B(n_943), .Y(n_945) );
BUFx3_ASAP7_75t_L g1273 ( .A(n_350), .Y(n_1273) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx2_ASAP7_75t_L g408 ( .A(n_351), .Y(n_408) );
NAND2x1p5_ASAP7_75t_L g491 ( .A(n_351), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g413 ( .A(n_352), .Y(n_413) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g492 ( .A(n_354), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_363), .Y(n_355) );
AOI33xp33_ASAP7_75t_L g519 ( .A1(n_356), .A2(n_520), .A3(n_521), .B1(n_525), .B2(n_529), .B3(n_530), .Y(n_519) );
AOI33xp33_ASAP7_75t_L g602 ( .A1(n_356), .A2(n_603), .A3(n_605), .B1(n_610), .B2(n_611), .B3(n_614), .Y(n_602) );
AOI33xp33_ASAP7_75t_L g1311 ( .A1(n_356), .A2(n_688), .A3(n_1312), .B1(n_1313), .B2(n_1317), .B3(n_1320), .Y(n_1311) );
AOI33xp33_ASAP7_75t_L g1351 ( .A1(n_356), .A2(n_1352), .A3(n_1353), .B1(n_1354), .B2(n_1355), .B3(n_1356), .Y(n_1351) );
BUFx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI33xp33_ASAP7_75t_L g776 ( .A1(n_357), .A2(n_777), .A3(n_779), .B1(n_783), .B2(n_785), .B3(n_786), .Y(n_776) );
AOI33xp33_ASAP7_75t_L g851 ( .A1(n_357), .A2(n_852), .A3(n_853), .B1(n_854), .B2(n_855), .B3(n_857), .Y(n_851) );
AOI33xp33_ASAP7_75t_L g1014 ( .A1(n_357), .A2(n_529), .A3(n_1015), .B1(n_1016), .B2(n_1019), .B3(n_1020), .Y(n_1014) );
AOI33xp33_ASAP7_75t_L g1060 ( .A1(n_357), .A2(n_614), .A3(n_1061), .B1(n_1062), .B2(n_1065), .B3(n_1066), .Y(n_1060) );
AOI33xp33_ASAP7_75t_L g1234 ( .A1(n_357), .A2(n_1235), .A3(n_1236), .B1(n_1238), .B2(n_1240), .B3(n_1241), .Y(n_1234) );
AOI33xp33_ASAP7_75t_L g1268 ( .A1(n_357), .A2(n_529), .A3(n_1269), .B1(n_1270), .B2(n_1274), .B3(n_1275), .Y(n_1268) );
AND3x4_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .C(n_361), .Y(n_357) );
INVx1_ASAP7_75t_L g394 ( .A(n_358), .Y(n_394) );
NAND2xp33_ASAP7_75t_SL g677 ( .A(n_358), .B(n_360), .Y(n_677) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_358), .B(n_359), .Y(n_1165) );
BUFx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx3_ASAP7_75t_L g377 ( .A(n_360), .Y(n_377) );
INVx2_ASAP7_75t_SL g482 ( .A(n_361), .Y(n_482) );
INVx1_ASAP7_75t_L g588 ( .A(n_361), .Y(n_588) );
OAI31xp33_ASAP7_75t_SL g958 ( .A1(n_361), .A2(n_959), .A3(n_960), .B(n_964), .Y(n_958) );
OAI31xp33_ASAP7_75t_L g1154 ( .A1(n_361), .A2(n_1155), .A3(n_1156), .B(n_1173), .Y(n_1154) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx2_ASAP7_75t_L g720 ( .A(n_362), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_362), .B(n_456), .Y(n_876) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g1277 ( .A(n_366), .Y(n_1277) );
BUFx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2x1p5_ASAP7_75t_L g399 ( .A(n_367), .B(n_393), .Y(n_399) );
INVx8_ASAP7_75t_L g499 ( .A(n_367), .Y(n_499) );
BUFx3_ASAP7_75t_L g921 ( .A(n_367), .Y(n_921) );
AND2x2_ASAP7_75t_L g924 ( .A(n_367), .B(n_925), .Y(n_924) );
HB1xp67_ASAP7_75t_L g1657 ( .A(n_367), .Y(n_1657) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g390 ( .A(n_371), .B(n_391), .Y(n_390) );
BUFx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx2_ASAP7_75t_L g384 ( .A(n_372), .Y(n_384) );
INVx2_ASAP7_75t_L g609 ( .A(n_372), .Y(n_609) );
BUFx2_ASAP7_75t_L g686 ( .A(n_372), .Y(n_686) );
BUFx3_ASAP7_75t_L g914 ( .A(n_372), .Y(n_914) );
AND2x2_ASAP7_75t_L g927 ( .A(n_372), .B(n_925), .Y(n_927) );
BUFx2_ASAP7_75t_L g1021 ( .A(n_372), .Y(n_1021) );
NAND3xp33_ASAP7_75t_L g373 ( .A(n_374), .B(n_381), .C(n_385), .Y(n_373) );
INVx1_ASAP7_75t_L g1122 ( .A(n_374), .Y(n_1122) );
BUFx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g529 ( .A(n_375), .Y(n_529) );
BUFx2_ASAP7_75t_L g614 ( .A(n_375), .Y(n_614) );
BUFx2_ASAP7_75t_L g1355 ( .A(n_375), .Y(n_1355) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx3_ASAP7_75t_L g688 ( .A(n_376), .Y(n_688) );
NAND3x1_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .C(n_380), .Y(n_376) );
AND2x4_ASAP7_75t_L g393 ( .A(n_377), .B(n_394), .Y(n_393) );
NAND2x1p5_ASAP7_75t_L g788 ( .A(n_377), .B(n_380), .Y(n_788) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g392 ( .A(n_379), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_379), .B(n_420), .Y(n_897) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND3xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_395), .C(n_404), .Y(n_388) );
AND4x1_ASAP7_75t_L g769 ( .A(n_389), .B(n_770), .C(n_774), .D(n_776), .Y(n_769) );
INVx1_ASAP7_75t_L g1024 ( .A(n_389), .Y(n_1024) );
NAND4xp25_ASAP7_75t_SL g1054 ( .A(n_389), .B(n_1055), .C(n_1058), .D(n_1060), .Y(n_1054) );
NAND4xp25_ASAP7_75t_SL g1304 ( .A(n_389), .B(n_1305), .C(n_1309), .D(n_1311), .Y(n_1304) );
NAND2xp5_ASAP7_75t_SL g1348 ( .A(n_389), .B(n_1349), .Y(n_1348) );
INVx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_390), .Y(n_539) );
INVx3_ASAP7_75t_L g615 ( .A(n_390), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g746 ( .A(n_390), .B(n_747), .C(n_759), .Y(n_746) );
AOI211xp5_ASAP7_75t_L g848 ( .A1(n_390), .A2(n_397), .B(n_840), .C(n_849), .Y(n_848) );
AOI221xp5_ASAP7_75t_L g1242 ( .A1(n_390), .A2(n_699), .B1(n_772), .B2(n_1224), .C(n_1243), .Y(n_1242) );
AND2x2_ASAP7_75t_L g406 ( .A(n_391), .B(n_407), .Y(n_406) );
AND2x4_ASAP7_75t_L g410 ( .A(n_391), .B(n_411), .Y(n_410) );
NAND2x1_ASAP7_75t_L g596 ( .A(n_391), .B(n_407), .Y(n_596) );
AND2x4_ASAP7_75t_SL g699 ( .A(n_391), .B(n_411), .Y(n_699) );
AND2x4_ASAP7_75t_SL g772 ( .A(n_391), .B(n_407), .Y(n_772) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_391), .B(n_407), .Y(n_1307) );
AND2x4_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
OR2x2_ASAP7_75t_L g509 ( .A(n_392), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g892 ( .A(n_392), .Y(n_892) );
AND2x6_ASAP7_75t_L g934 ( .A(n_393), .B(n_407), .Y(n_934) );
AND2x2_ASAP7_75t_L g936 ( .A(n_393), .B(n_413), .Y(n_936) );
INVx1_ASAP7_75t_L g939 ( .A(n_393), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
AOI221xp5_ASAP7_75t_SL g432 ( .A1(n_396), .A2(n_433), .B1(n_446), .B2(n_453), .C(n_454), .Y(n_432) );
INVx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx5_ASAP7_75t_L g601 ( .A(n_398), .Y(n_601) );
OR2x6_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
OR2x2_ASAP7_75t_L g672 ( .A(n_399), .B(n_400), .Y(n_672) );
INVx2_ASAP7_75t_L g931 ( .A(n_399), .Y(n_931) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g485 ( .A(n_401), .B(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g879 ( .A(n_401), .B(n_486), .Y(n_879) );
INVx1_ASAP7_75t_L g907 ( .A(n_401), .Y(n_907) );
BUFx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g494 ( .A(n_402), .Y(n_494) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B1(n_409), .B2(n_410), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_406), .A2(n_410), .B1(n_517), .B2(n_518), .Y(n_516) );
AO22x1_ASAP7_75t_L g1345 ( .A1(n_406), .A2(n_410), .B1(n_1346), .B2(n_1347), .Y(n_1345) );
INVx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_410), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_410), .A2(n_595), .B1(n_1012), .B2(n_1013), .Y(n_1011) );
AOI22xp5_ASAP7_75t_L g1055 ( .A1(n_410), .A2(n_595), .B1(n_1056), .B2(n_1057), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_410), .A2(n_595), .B1(n_1266), .B2(n_1267), .Y(n_1265) );
AOI22xp5_ASAP7_75t_L g1305 ( .A1(n_410), .A2(n_1306), .B1(n_1307), .B2(n_1308), .Y(n_1305) );
AOI221x1_ASAP7_75t_L g1645 ( .A1(n_410), .A2(n_595), .B1(n_1623), .B2(n_1628), .C(n_1646), .Y(n_1645) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AOI21xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_482), .B(n_483), .Y(n_414) );
NAND3xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_432), .C(n_457), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_427), .B2(n_428), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_417), .A2(n_427), .B1(n_497), .B2(n_501), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_418), .A2(n_428), .B1(n_707), .B2(n_708), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_418), .A2(n_428), .B1(n_799), .B2(n_800), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_418), .A2(n_428), .B1(n_844), .B2(n_845), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_418), .A2(n_428), .B1(n_1082), .B2(n_1083), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1330 ( .A1(n_418), .A2(n_1038), .B1(n_1331), .B2(n_1332), .Y(n_1330) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g561 ( .A(n_419), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_419), .A2(n_428), .B1(n_735), .B2(n_736), .Y(n_734) );
AND2x4_ASAP7_75t_L g906 ( .A(n_419), .B(n_907), .Y(n_906) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
AND2x4_ASAP7_75t_L g428 ( .A(n_420), .B(n_429), .Y(n_428) );
AND2x4_ASAP7_75t_L g453 ( .A(n_420), .B(n_450), .Y(n_453) );
AND2x4_ASAP7_75t_SL g477 ( .A(n_420), .B(n_455), .Y(n_477) );
AND2x2_ASAP7_75t_L g838 ( .A(n_420), .B(n_839), .Y(n_838) );
AND2x2_ASAP7_75t_L g949 ( .A(n_420), .B(n_429), .Y(n_949) );
BUFx2_ASAP7_75t_L g1229 ( .A(n_420), .Y(n_1229) );
INVx3_ASAP7_75t_L g448 ( .A(n_422), .Y(n_448) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_422), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_422), .B(n_456), .Y(n_510) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_425), .Y(n_422) );
OR2x2_ASAP7_75t_L g643 ( .A(n_423), .B(n_426), .Y(n_643) );
HB1xp67_ASAP7_75t_L g1226 ( .A(n_423), .Y(n_1226) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g430 ( .A(n_424), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g441 ( .A(n_424), .B(n_426), .Y(n_441) );
INVx2_ASAP7_75t_L g452 ( .A(n_424), .Y(n_452) );
INVx1_ASAP7_75t_L g488 ( .A(n_424), .Y(n_488) );
OR2x2_ASAP7_75t_L g578 ( .A(n_424), .B(n_426), .Y(n_578) );
NAND2x1_ASAP7_75t_L g638 ( .A(n_424), .B(n_426), .Y(n_638) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g431 ( .A(n_426), .Y(n_431) );
AND2x2_ASAP7_75t_L g451 ( .A(n_426), .B(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_L g481 ( .A(n_426), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_426), .B(n_452), .Y(n_569) );
INVx1_ASAP7_75t_L g564 ( .A(n_428), .Y(n_564) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_428), .Y(n_631) );
BUFx6f_ASAP7_75t_L g1038 ( .A(n_428), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1363 ( .A1(n_428), .A2(n_560), .B1(n_1359), .B2(n_1360), .Y(n_1363) );
INVx2_ASAP7_75t_L g461 ( .A(n_429), .Y(n_461) );
INVx1_ASAP7_75t_L g731 ( .A(n_429), .Y(n_731) );
BUFx6f_ASAP7_75t_L g795 ( .A(n_429), .Y(n_795) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g437 ( .A(n_430), .Y(n_437) );
BUFx3_ASAP7_75t_L g704 ( .A(n_430), .Y(n_704) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g1298 ( .A(n_435), .Y(n_1298) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_436), .Y(n_572) );
INVx1_ASAP7_75t_L g1048 ( .A(n_436), .Y(n_1048) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g622 ( .A(n_437), .Y(n_622) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g834 ( .A(n_439), .Y(n_834) );
INVx1_ASAP7_75t_L g1366 ( .A(n_439), .Y(n_1366) );
BUFx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_441), .Y(n_455) );
INVx4_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx4_ASAP7_75t_L g553 ( .A(n_443), .Y(n_553) );
INVx1_ASAP7_75t_SL g623 ( .A(n_443), .Y(n_623) );
AND2x2_ASAP7_75t_SL g872 ( .A(n_443), .B(n_494), .Y(n_872) );
AND2x4_ASAP7_75t_L g991 ( .A(n_443), .B(n_992), .Y(n_991) );
NAND4xp25_ASAP7_75t_L g1633 ( .A(n_443), .B(n_1634), .C(n_1635), .D(n_1636), .Y(n_1633) );
AND2x4_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx2_ASAP7_75t_L g473 ( .A(n_444), .Y(n_473) );
AND2x4_ASAP7_75t_L g472 ( .A(n_445), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g1395 ( .A(n_445), .Y(n_1395) );
INVx2_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g555 ( .A(n_448), .Y(n_555) );
INVx1_ASAP7_75t_L g797 ( .A(n_448), .Y(n_797) );
INVx2_ASAP7_75t_L g1032 ( .A(n_448), .Y(n_1032) );
INVx1_ASAP7_75t_L g1133 ( .A(n_448), .Y(n_1133) );
INVx2_ASAP7_75t_L g1184 ( .A(n_448), .Y(n_1184) );
BUFx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g628 ( .A(n_450), .Y(n_628) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g467 ( .A(n_451), .Y(n_467) );
BUFx3_ASAP7_75t_L g557 ( .A(n_451), .Y(n_557) );
BUFx3_ASAP7_75t_L g733 ( .A(n_451), .Y(n_733) );
INVx3_ASAP7_75t_L g545 ( .A(n_453), .Y(n_545) );
INVx2_ASAP7_75t_SL g618 ( .A(n_453), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_453), .B(n_775), .Y(n_801) );
NAND2xp5_ASAP7_75t_R g1369 ( .A(n_453), .B(n_1350), .Y(n_1369) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_454), .A2(n_547), .B(n_554), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_454), .A2(n_620), .B(n_624), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_454), .A2(n_703), .B(n_705), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_454), .A2(n_728), .B(n_732), .Y(n_727) );
INVx1_ASAP7_75t_L g802 ( .A(n_454), .Y(n_802) );
AOI221xp5_ASAP7_75t_L g837 ( .A1(n_454), .A2(n_838), .B1(n_840), .B2(n_841), .C(n_842), .Y(n_837) );
AOI21xp5_ASAP7_75t_L g1030 ( .A1(n_454), .A2(n_1031), .B(n_1033), .Y(n_1030) );
AOI21xp5_ASAP7_75t_L g1078 ( .A1(n_454), .A2(n_1079), .B(n_1080), .Y(n_1078) );
AOI21xp5_ASAP7_75t_L g1129 ( .A1(n_454), .A2(n_1130), .B(n_1132), .Y(n_1129) );
AOI21xp5_ASAP7_75t_SL g1284 ( .A1(n_454), .A2(n_1285), .B(n_1287), .Y(n_1284) );
AOI21xp5_ASAP7_75t_L g1327 ( .A1(n_454), .A2(n_1328), .B(n_1329), .Y(n_1327) );
AOI21xp5_ASAP7_75t_L g1364 ( .A1(n_454), .A2(n_1365), .B(n_1368), .Y(n_1364) );
AND2x6_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g470 ( .A(n_455), .Y(n_470) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_455), .Y(n_549) );
BUFx3_ASAP7_75t_L g621 ( .A(n_455), .Y(n_621) );
BUFx3_ASAP7_75t_L g729 ( .A(n_455), .Y(n_729) );
BUFx3_ASAP7_75t_L g1034 ( .A(n_455), .Y(n_1034) );
BUFx3_ASAP7_75t_L g1049 ( .A(n_455), .Y(n_1049) );
AND2x2_ASAP7_75t_L g479 ( .A(n_456), .B(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_456), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g582 ( .A(n_456), .Y(n_582) );
AOI31xp33_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_462), .A3(n_468), .B(n_474), .Y(n_457) );
BUFx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g552 ( .A(n_461), .Y(n_552) );
INVx2_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_465), .Y(n_626) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx3_ASAP7_75t_L g839 ( .A(n_467), .Y(n_839) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g645 ( .A(n_471), .Y(n_645) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g573 ( .A(n_472), .Y(n_573) );
INVx1_ASAP7_75t_L g743 ( .A(n_472), .Y(n_743) );
INVx3_ASAP7_75t_L g835 ( .A(n_472), .Y(n_835) );
OAI221xp5_ASAP7_75t_L g1372 ( .A1(n_472), .A2(n_640), .B1(n_870), .B2(n_1373), .C(n_1374), .Y(n_1372) );
INVxp67_ASAP7_75t_L g1398 ( .A(n_473), .Y(n_1398) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AOI222xp33_ASAP7_75t_L g830 ( .A1(n_476), .A2(n_479), .B1(n_831), .B2(n_832), .C1(n_833), .C2(n_836), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g1622 ( .A(n_476), .B(n_1623), .Y(n_1622) );
BUFx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g584 ( .A(n_477), .Y(n_584) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g1223 ( .A1(n_480), .A2(n_1224), .B1(n_1225), .B2(n_1227), .Y(n_1223) );
AOI22xp33_ASAP7_75t_L g1627 ( .A1(n_480), .A2(n_1225), .B1(n_1628), .B2(n_1629), .Y(n_1627) );
BUFx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g581 ( .A(n_481), .Y(n_581) );
INVx1_ASAP7_75t_L g878 ( .A(n_481), .Y(n_878) );
O2A1O1Ixp5_ASAP7_75t_L g616 ( .A1(n_482), .A2(n_617), .B(n_633), .C(n_656), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g1028 ( .A1(n_482), .A2(n_1029), .B(n_1039), .Y(n_1028) );
OAI21xp5_ASAP7_75t_L g1282 ( .A1(n_482), .A2(n_1283), .B(n_1291), .Y(n_1282) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_484), .Y(n_657) );
INVx2_ASAP7_75t_L g1073 ( .A(n_484), .Y(n_1073) );
AND2x4_ASAP7_75t_L g484 ( .A(n_485), .B(n_489), .Y(n_484) );
AND2x4_ASAP7_75t_L g671 ( .A(n_485), .B(n_489), .Y(n_671) );
INVx2_ASAP7_75t_SL g997 ( .A(n_485), .Y(n_997) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g1250 ( .A(n_489), .Y(n_1250) );
OR2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_493), .Y(n_489) );
INVx3_ASAP7_75t_L g978 ( .A(n_490), .Y(n_978) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g938 ( .A(n_491), .Y(n_938) );
INVx1_ASAP7_75t_L g500 ( .A(n_493), .Y(n_500) );
OR2x2_ASAP7_75t_L g505 ( .A(n_493), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g537 ( .A(n_493), .Y(n_537) );
OR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
OR2x2_ASAP7_75t_L g676 ( .A(n_494), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g993 ( .A(n_494), .Y(n_993) );
INVx1_ASAP7_75t_L g925 ( .A(n_495), .Y(n_925) );
INVx1_ASAP7_75t_L g943 ( .A(n_495), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_497), .A2(n_501), .B1(n_630), .B2(n_632), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_497), .A2(n_501), .B1(n_707), .B2(n_708), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_497), .A2(n_501), .B1(n_735), .B2(n_736), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_497), .A2(n_817), .B1(n_844), .B2(n_845), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_497), .A2(n_501), .B1(n_1359), .B2(n_1360), .Y(n_1358) );
AND2x4_ASAP7_75t_L g497 ( .A(n_498), .B(n_500), .Y(n_497) );
AND2x4_ASAP7_75t_L g816 ( .A(n_498), .B(n_500), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g1174 ( .A1(n_498), .A2(n_856), .B1(n_1152), .B2(n_1175), .Y(n_1174) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx3_ASAP7_75t_L g604 ( .A(n_499), .Y(n_604) );
INVx8_ASAP7_75t_L g613 ( .A(n_499), .Y(n_613) );
CKINVDCx5p33_ASAP7_75t_R g970 ( .A(n_499), .Y(n_970) );
INVx2_ASAP7_75t_L g538 ( .A(n_501), .Y(n_538) );
INVx2_ASAP7_75t_L g1103 ( .A(n_501), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_511), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_503), .A2(n_541), .B(n_542), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_503), .B(n_660), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_503), .A2(n_669), .B(n_670), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_503), .A2(n_761), .B(n_762), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_503), .B(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_503), .B(n_826), .Y(n_825) );
AOI21xp33_ASAP7_75t_SL g1025 ( .A1(n_503), .A2(n_1026), .B(n_1027), .Y(n_1025) );
NAND2xp33_ASAP7_75t_L g1067 ( .A(n_503), .B(n_1068), .Y(n_1067) );
AOI21xp33_ASAP7_75t_L g1139 ( .A1(n_503), .A2(n_1140), .B(n_1141), .Y(n_1139) );
AOI21xp33_ASAP7_75t_SL g1279 ( .A1(n_503), .A2(n_1280), .B(n_1281), .Y(n_1279) );
AOI211x1_ASAP7_75t_L g1302 ( .A1(n_503), .A2(n_1303), .B(n_1304), .C(n_1321), .Y(n_1302) );
AOI211x1_ASAP7_75t_L g1341 ( .A1(n_503), .A2(n_1342), .B(n_1343), .C(n_1357), .Y(n_1341) );
INVx8_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_509), .Y(n_504) );
INVx1_ASAP7_75t_L g1252 ( .A(n_505), .Y(n_1252) );
BUFx3_ASAP7_75t_L g967 ( .A(n_506), .Y(n_967) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_507), .Y(n_694) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g683 ( .A(n_508), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_509), .B(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_L g893 ( .A(n_510), .Y(n_893) );
INVx1_ASAP7_75t_L g589 ( .A(n_512), .Y(n_589) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_540), .C(n_543), .Y(n_513) );
NOR3xp33_ASAP7_75t_L g514 ( .A(n_515), .B(n_531), .C(n_539), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_519), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_517), .A2(n_518), .B1(n_580), .B2(n_583), .Y(n_579) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OAI221xp5_ASAP7_75t_L g678 ( .A1(n_524), .A2(n_679), .B1(n_680), .B2(n_684), .C(n_685), .Y(n_678) );
INVx3_ASAP7_75t_L g818 ( .A(n_524), .Y(n_818) );
INVx1_ASAP7_75t_L g911 ( .A(n_524), .Y(n_911) );
OR2x6_ASAP7_75t_SL g941 ( .A(n_524), .B(n_942), .Y(n_941) );
BUFx2_ASAP7_75t_L g1315 ( .A(n_524), .Y(n_1315) );
INVx8_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g607 ( .A(n_527), .Y(n_607) );
OAI221xp5_ASAP7_75t_L g1654 ( .A1(n_527), .A2(n_967), .B1(n_1638), .B2(n_1655), .C(n_1656), .Y(n_1654) );
INVx5_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx3_ASAP7_75t_L g917 ( .A(n_528), .Y(n_917) );
INVx2_ASAP7_75t_SL g1064 ( .A(n_528), .Y(n_1064) );
INVx2_ASAP7_75t_SL g1167 ( .A(n_528), .Y(n_1167) );
NAND2xp5_ASAP7_75t_L g1660 ( .A(n_532), .B(n_905), .Y(n_1660) );
OR2x6_ASAP7_75t_L g532 ( .A(n_533), .B(n_536), .Y(n_532) );
OR2x2_ASAP7_75t_L g1023 ( .A(n_533), .B(n_536), .Y(n_1023) );
INVx2_ASAP7_75t_SL g1112 ( .A(n_533), .Y(n_1112) );
INVx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx4f_ASAP7_75t_L g1158 ( .A(n_535), .Y(n_1158) );
INVxp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g817 ( .A(n_537), .B(n_818), .Y(n_817) );
NOR3xp33_ASAP7_75t_L g673 ( .A(n_539), .B(n_674), .C(n_697), .Y(n_673) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_565), .B(n_585), .Y(n_543) );
BUFx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
HB1xp67_ASAP7_75t_L g1286 ( .A(n_552), .Y(n_1286) );
HB1xp67_ASAP7_75t_SL g1131 ( .A(n_553), .Y(n_1131) );
BUFx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_SL g1135 ( .A(n_557), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B1(n_562), .B2(n_563), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_560), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g1035 ( .A1(n_560), .A2(n_1036), .B1(n_1037), .B2(n_1038), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_560), .A2(n_631), .B1(n_1137), .B2(n_1138), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1288 ( .A1(n_560), .A2(n_1038), .B1(n_1289), .B2(n_1290), .Y(n_1288) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx5_ASAP7_75t_L g1378 ( .A(n_566), .Y(n_1378) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g652 ( .A(n_567), .Y(n_652) );
INVx2_ASAP7_75t_L g813 ( .A(n_567), .Y(n_813) );
INVx2_ASAP7_75t_SL g1044 ( .A(n_567), .Y(n_1044) );
INVx4_ASAP7_75t_L g1632 ( .A(n_567), .Y(n_1632) );
INVx8_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx2_ASAP7_75t_L g884 ( .A(n_568), .Y(n_884) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_574), .Y(n_570) );
INVx1_ASAP7_75t_L g811 ( .A(n_575), .Y(n_811) );
INVxp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x6_ASAP7_75t_L g1397 ( .A(n_576), .B(n_1398), .Y(n_1397) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx3_ASAP7_75t_L g649 ( .A(n_577), .Y(n_649) );
BUFx4f_ASAP7_75t_L g1222 ( .A(n_577), .Y(n_1222) );
INVx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g655 ( .A(n_580), .Y(n_655) );
INVx2_ASAP7_75t_L g1040 ( .A(n_580), .Y(n_1040) );
NOR2x1_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx1_ASAP7_75t_L g1228 ( .A(n_582), .Y(n_1228) );
INVx2_ASAP7_75t_L g634 ( .A(n_583), .Y(n_634) );
INVx2_ASAP7_75t_L g710 ( .A(n_583), .Y(n_710) );
INVx1_ASAP7_75t_L g1371 ( .A(n_583), .Y(n_1371) );
INVx4_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OAI21xp5_ASAP7_75t_L g1124 ( .A1(n_585), .A2(n_1125), .B(n_1128), .Y(n_1124) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
A2O1A1Ixp33_ASAP7_75t_L g908 ( .A1(n_587), .A2(n_909), .B(n_928), .C(n_946), .Y(n_908) );
HB1xp67_ASAP7_75t_L g1641 ( .A(n_587), .Y(n_1641) );
BUFx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
BUFx2_ASAP7_75t_L g745 ( .A(n_588), .Y(n_745) );
AOI21x1_ASAP7_75t_L g1211 ( .A1(n_588), .A2(n_1212), .B(n_1232), .Y(n_1211) );
XOR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_661), .Y(n_590) );
NAND3x1_ASAP7_75t_SL g591 ( .A(n_592), .B(n_616), .C(n_659), .Y(n_591) );
AND4x1_ASAP7_75t_L g592 ( .A(n_593), .B(n_599), .C(n_602), .D(n_615), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B1(n_597), .B2(n_598), .Y(n_593) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g1101 ( .A(n_598), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_601), .B(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_601), .B(n_1059), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_601), .B(n_1310), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_601), .B(n_1350), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1661 ( .A(n_601), .B(n_1662), .Y(n_1661) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_607), .A2(n_1111), .B1(n_1113), .B2(n_1114), .Y(n_1110) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g758 ( .A(n_609), .Y(n_758) );
INVx1_ASAP7_75t_L g778 ( .A(n_609), .Y(n_778) );
INVx2_ASAP7_75t_L g856 ( .A(n_609), .Y(n_856) );
BUFx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_SL g1123 ( .A(n_615), .Y(n_1123) );
AND5x1_ASAP7_75t_L g1619 ( .A(n_615), .B(n_1620), .C(n_1645), .D(n_1658), .E(n_1661), .Y(n_1619) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI221xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_639), .B1(n_640), .B2(n_644), .C(n_645), .Y(n_635) );
BUFx2_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_SL g741 ( .A(n_637), .Y(n_741) );
OR2x2_ASAP7_75t_L g900 ( .A(n_637), .B(n_897), .Y(n_900) );
OR2x2_ASAP7_75t_L g1190 ( .A(n_637), .B(n_897), .Y(n_1190) );
BUFx3_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_638), .Y(n_714) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx4_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
BUFx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
BUFx3_ASAP7_75t_L g807 ( .A(n_643), .Y(n_807) );
INVx1_ASAP7_75t_L g1194 ( .A(n_643), .Y(n_1194) );
BUFx2_ASAP7_75t_L g1631 ( .A(n_643), .Y(n_1631) );
OAI221xp5_ASAP7_75t_L g804 ( .A1(n_645), .A2(n_805), .B1(n_806), .B2(n_807), .C(n_808), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B1(n_650), .B2(n_653), .Y(n_646) );
INVx1_ASAP7_75t_L g866 ( .A(n_648), .Y(n_866) );
OAI221xp5_ASAP7_75t_L g1041 ( .A1(n_648), .A2(n_1042), .B1(n_1043), .B2(n_1045), .C(n_1046), .Y(n_1041) );
OAI221xp5_ASAP7_75t_SL g1126 ( .A1(n_648), .A2(n_650), .B1(n_1113), .B2(n_1120), .C(n_1127), .Y(n_1126) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_649), .A2(n_813), .B1(n_985), .B2(n_986), .Y(n_984) );
OAI22x1_ASAP7_75t_SL g989 ( .A1(n_649), .A2(n_813), .B1(n_968), .B2(n_990), .Y(n_989) );
BUFx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g865 ( .A(n_651), .Y(n_865) );
OAI221xp5_ASAP7_75t_L g1292 ( .A1(n_651), .A2(n_1293), .B1(n_1295), .B2(n_1296), .C(n_1297), .Y(n_1292) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
BUFx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
XNOR2x1_ASAP7_75t_L g663 ( .A(n_664), .B(n_765), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AO22x2_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_722), .B1(n_723), .B2(n_764), .Y(n_665) );
INVx1_ASAP7_75t_L g764 ( .A(n_666), .Y(n_764) );
AND4x1_ASAP7_75t_L g667 ( .A(n_668), .B(n_673), .C(n_700), .D(n_721), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_672), .B(n_1200), .Y(n_1199) );
OAI22xp5_ASAP7_75t_SL g674 ( .A1(n_675), .A2(n_678), .B1(n_687), .B2(n_689), .Y(n_674) );
BUFx4f_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
BUFx8_ASAP7_75t_L g748 ( .A(n_676), .Y(n_748) );
BUFx2_ASAP7_75t_L g1647 ( .A(n_676), .Y(n_1647) );
BUFx2_ASAP7_75t_L g918 ( .A(n_677), .Y(n_918) );
OAI221xp5_ASAP7_75t_L g749 ( .A1(n_680), .A2(n_750), .B1(n_751), .B2(n_752), .C(n_753), .Y(n_749) );
INVx3_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
BUFx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
CKINVDCx5p33_ASAP7_75t_R g754 ( .A(n_688), .Y(n_754) );
INVx2_ASAP7_75t_L g1653 ( .A(n_688), .Y(n_1653) );
OAI221xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_692), .B1(n_693), .B2(n_695), .C(n_696), .Y(n_689) );
INVx1_ASAP7_75t_L g780 ( .A(n_690), .Y(n_780) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g1018 ( .A(n_691), .Y(n_1018) );
BUFx6f_ASAP7_75t_L g1237 ( .A(n_691), .Y(n_1237) );
BUFx6f_ASAP7_75t_L g1239 ( .A(n_691), .Y(n_1239) );
OAI211xp5_ASAP7_75t_L g711 ( .A1(n_692), .A2(n_712), .B(n_715), .C(n_716), .Y(n_711) );
OAI221xp5_ASAP7_75t_L g755 ( .A1(n_693), .A2(n_739), .B1(n_750), .B2(n_756), .C(n_757), .Y(n_755) );
CKINVDCx8_ASAP7_75t_R g693 ( .A(n_694), .Y(n_693) );
INVx3_ASAP7_75t_L g1106 ( .A(n_694), .Y(n_1106) );
INVx3_ASAP7_75t_L g1160 ( .A(n_694), .Y(n_1160) );
INVx3_ASAP7_75t_L g1650 ( .A(n_694), .Y(n_1650) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_699), .A2(n_771), .B1(n_772), .B2(n_773), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_699), .A2(n_772), .B1(n_831), .B2(n_832), .Y(n_850) );
OAI21xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_709), .B(n_717), .Y(n_700) );
INVx1_ASAP7_75t_L g1090 ( .A(n_704), .Y(n_1090) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g805 ( .A(n_713), .Y(n_805) );
INVx2_ASAP7_75t_L g1087 ( .A(n_713), .Y(n_1087) );
INVx4_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
BUFx4f_ASAP7_75t_L g793 ( .A(n_714), .Y(n_793) );
BUFx4f_ASAP7_75t_L g870 ( .A(n_714), .Y(n_870) );
OR2x6_ASAP7_75t_L g880 ( .A(n_714), .B(n_881), .Y(n_880) );
BUFx4f_ASAP7_75t_L g1231 ( .A(n_714), .Y(n_1231) );
OAI21xp5_ASAP7_75t_L g1076 ( .A1(n_717), .A2(n_1077), .B(n_1084), .Y(n_1076) );
OAI21xp5_ASAP7_75t_L g1361 ( .A1(n_717), .A2(n_1362), .B(n_1370), .Y(n_1361) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g828 ( .A(n_718), .Y(n_828) );
BUFx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g1204 ( .A(n_719), .B(n_945), .Y(n_1204) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OR2x6_ASAP7_75t_L g787 ( .A(n_720), .B(n_788), .Y(n_787) );
AND2x4_ASAP7_75t_L g888 ( .A(n_720), .B(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AND4x1_ASAP7_75t_L g724 ( .A(n_725), .B(n_746), .C(n_760), .D(n_763), .Y(n_724) );
OAI21xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_737), .B(n_745), .Y(n_725) );
INVx2_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
OAI211xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .B(n_742), .C(n_744), .Y(n_738) );
OAI211xp5_ASAP7_75t_L g1334 ( .A1(n_740), .A2(n_1335), .B(n_1336), .C(n_1337), .Y(n_1334) );
OAI211xp5_ASAP7_75t_L g1637 ( .A1(n_740), .A2(n_1638), .B(n_1639), .C(n_1640), .Y(n_1637) );
INVx5_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
O2A1O1Ixp5_ASAP7_75t_SL g789 ( .A1(n_745), .A2(n_790), .B(n_803), .C(n_814), .Y(n_789) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_748), .A2(n_749), .B1(n_754), .B2(n_755), .Y(n_747) );
OAI33xp33_ASAP7_75t_L g1104 ( .A1(n_748), .A2(n_1105), .A3(n_1110), .B1(n_1115), .B2(n_1119), .B3(n_1122), .Y(n_1104) );
XOR2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_859), .Y(n_765) );
XNOR2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_822), .Y(n_766) );
XOR2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_821), .Y(n_767) );
NAND3xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_789), .C(n_819), .Y(n_768) );
INVx2_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g784 ( .A(n_782), .Y(n_784) );
INVx1_ASAP7_75t_L g1316 ( .A(n_782), .Y(n_1316) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_SL g857 ( .A(n_787), .Y(n_857) );
INVx1_ASAP7_75t_L g1241 ( .A(n_787), .Y(n_1241) );
INVx3_ASAP7_75t_L g972 ( .A(n_788), .Y(n_972) );
NAND4xp25_ASAP7_75t_L g790 ( .A(n_791), .B(n_798), .C(n_801), .D(n_802), .Y(n_790) );
OAI211xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_793), .B(n_794), .C(n_796), .Y(n_791) );
BUFx3_ASAP7_75t_L g1367 ( .A(n_795), .Y(n_1367) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_799), .A2(n_800), .B1(n_816), .B2(n_817), .Y(n_815) );
INVx2_ASAP7_75t_L g868 ( .A(n_807), .Y(n_868) );
OAI221xp5_ASAP7_75t_L g885 ( .A1(n_807), .A2(n_870), .B1(n_886), .B2(n_887), .C(n_888), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_809) );
AOI222xp33_ASAP7_75t_L g1249 ( .A1(n_816), .A2(n_1227), .B1(n_1250), .B2(n_1251), .C1(n_1252), .C2(n_1253), .Y(n_1249) );
INVx2_ASAP7_75t_SL g1246 ( .A(n_817), .Y(n_1246) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
NAND3xp33_ASAP7_75t_L g824 ( .A(n_825), .B(n_827), .C(n_848), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_829), .B(n_846), .Y(n_827) );
OAI21xp33_ASAP7_75t_L g1325 ( .A1(n_828), .A2(n_1326), .B(n_1333), .Y(n_1325) );
NAND3xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_837), .C(n_843), .Y(n_829) );
INVx2_ASAP7_75t_L g1213 ( .A(n_838), .Y(n_1213) );
AND2x4_ASAP7_75t_L g895 ( .A(n_839), .B(n_896), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
XNOR2x1_ASAP7_75t_L g859 ( .A(n_860), .B(n_951), .Y(n_859) );
XNOR2x1_ASAP7_75t_L g860 ( .A(n_861), .B(n_950), .Y(n_860) );
OR2x2_ASAP7_75t_L g861 ( .A(n_862), .B(n_908), .Y(n_861) );
NAND3xp33_ASAP7_75t_SL g862 ( .A(n_863), .B(n_890), .C(n_902), .Y(n_862) );
AOI211xp5_ASAP7_75t_SL g863 ( .A1(n_864), .A2(n_867), .B(n_873), .C(n_882), .Y(n_863) );
INVxp67_ASAP7_75t_SL g869 ( .A(n_870), .Y(n_869) );
OAI21xp5_ASAP7_75t_L g1191 ( .A1(n_871), .A2(n_880), .B(n_1192), .Y(n_1191) );
INVx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g996 ( .A(n_874), .Y(n_996) );
INVx2_ASAP7_75t_SL g1188 ( .A(n_874), .Y(n_1188) );
NAND2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_877), .Y(n_874) );
INVx1_ASAP7_75t_L g881 ( .A(n_875), .Y(n_881) );
INVx2_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx2_ASAP7_75t_SL g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_SL g1186 ( .A(n_879), .Y(n_1186) );
CKINVDCx5p33_ASAP7_75t_R g1000 ( .A(n_880), .Y(n_1000) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
HB1xp67_ASAP7_75t_L g987 ( .A(n_888), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_888), .B(n_1182), .Y(n_1181) );
AOI222xp33_ASAP7_75t_L g890 ( .A1(n_891), .A2(n_894), .B1(n_895), .B2(n_898), .C1(n_899), .C2(n_901), .Y(n_890) );
AOI21xp33_ASAP7_75t_SL g998 ( .A1(n_891), .A2(n_999), .B(n_1000), .Y(n_998) );
AND2x4_ASAP7_75t_L g891 ( .A(n_892), .B(n_893), .Y(n_891) );
AOI222xp33_ASAP7_75t_L g994 ( .A1(n_895), .A2(n_962), .B1(n_974), .B2(n_995), .C1(n_996), .C2(n_997), .Y(n_994) );
INVx1_ASAP7_75t_L g1200 ( .A(n_895), .Y(n_1200) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
AOI211xp5_ASAP7_75t_L g928 ( .A1(n_898), .A2(n_929), .B(n_932), .C(n_940), .Y(n_928) );
AOI222xp33_ASAP7_75t_L g982 ( .A1(n_899), .A2(n_963), .B1(n_983), .B2(n_987), .C1(n_988), .C2(n_991), .Y(n_982) );
INVx2_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .Y(n_902) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx3_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
HB1xp67_ASAP7_75t_L g953 ( .A(n_906), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_906), .A2(n_948), .B1(n_1152), .B2(n_1153), .Y(n_1151) );
AND2x4_ASAP7_75t_L g948 ( .A(n_907), .B(n_949), .Y(n_948) );
AOI221xp5_ASAP7_75t_L g909 ( .A1(n_910), .A2(n_913), .B1(n_915), .B2(n_919), .C(n_922), .Y(n_909) );
INVx2_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
OAI221xp5_ASAP7_75t_L g965 ( .A1(n_917), .A2(n_966), .B1(n_967), .B2(n_968), .C(n_969), .Y(n_965) );
OAI221xp5_ASAP7_75t_L g1162 ( .A1(n_917), .A2(n_938), .B1(n_1163), .B2(n_1164), .C(n_1165), .Y(n_1162) );
BUFx2_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx2_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
AOI22xp5_ASAP7_75t_L g973 ( .A1(n_924), .A2(n_927), .B1(n_954), .B2(n_974), .Y(n_973) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx2_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx4_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_934), .A2(n_936), .B1(n_962), .B2(n_963), .Y(n_961) );
INVx2_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
OAI221xp5_ASAP7_75t_L g1156 ( .A1(n_937), .A2(n_1157), .B1(n_1162), .B2(n_1166), .C(n_1170), .Y(n_1156) );
OR2x6_ASAP7_75t_L g937 ( .A(n_938), .B(n_939), .Y(n_937) );
INVx2_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
HB1xp67_ASAP7_75t_L g1177 ( .A(n_943), .Y(n_1177) );
INVx3_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_947), .B(n_948), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_948), .B(n_957), .Y(n_956) );
INVx2_ASAP7_75t_L g1247 ( .A(n_948), .Y(n_1247) );
AOI211x1_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_954), .B(n_955), .C(n_981), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_956), .B(n_958), .Y(n_955) );
NAND3xp33_ASAP7_75t_L g964 ( .A(n_965), .B(n_973), .C(n_975), .Y(n_964) );
INVx3_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
OAI211xp5_ASAP7_75t_L g975 ( .A1(n_976), .A2(n_977), .B(n_979), .C(n_980), .Y(n_975) );
OAI21xp5_ASAP7_75t_SL g1170 ( .A1(n_977), .A2(n_1171), .B(n_1172), .Y(n_1170) );
INVx3_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx2_ASAP7_75t_L g1108 ( .A(n_978), .Y(n_1108) );
NAND3xp33_ASAP7_75t_L g981 ( .A(n_982), .B(n_994), .C(n_998), .Y(n_981) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
XNOR2xp5_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1143), .Y(n_1001) );
INVx2_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
AO22x2_ASAP7_75t_L g1003 ( .A1(n_1004), .A2(n_1005), .B1(n_1096), .B2(n_1142), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
OAI22xp5_ASAP7_75t_L g1005 ( .A1(n_1006), .A2(n_1007), .B1(n_1050), .B2(n_1095), .Y(n_1005) );
INVx2_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
NAND3xp33_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1025), .C(n_1028), .Y(n_1008) );
NOR3xp33_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1022), .C(n_1024), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1014), .Y(n_1010) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
HB1xp67_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx2_ASAP7_75t_L g1095 ( .A(n_1050), .Y(n_1095) );
NAND2x1p5_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1069), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1067), .Y(n_1052) );
INVxp67_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
NOR2xp33_ASAP7_75t_SL g1092 ( .A(n_1054), .B(n_1093), .Y(n_1092) );
INVx2_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1067), .B(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1076), .Y(n_1071) );
AOI21xp5_ASAP7_75t_L g1072 ( .A1(n_1073), .A2(n_1074), .B(n_1075), .Y(n_1072) );
AOI21xp5_ASAP7_75t_L g1322 ( .A1(n_1073), .A2(n_1323), .B(n_1324), .Y(n_1322) );
OAI211xp5_ASAP7_75t_L g1085 ( .A1(n_1086), .A2(n_1087), .B(n_1088), .C(n_1091), .Y(n_1085) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1096), .Y(n_1142) );
XNOR2xp5_ASAP7_75t_SL g1096 ( .A(n_1097), .B(n_1098), .Y(n_1096) );
AND3x2_ASAP7_75t_L g1098 ( .A(n_1099), .B(n_1124), .C(n_1139), .Y(n_1098) );
NOR4xp25_ASAP7_75t_L g1099 ( .A(n_1100), .B(n_1102), .C(n_1104), .D(n_1123), .Y(n_1099) );
OAI22xp33_ASAP7_75t_L g1105 ( .A1(n_1106), .A2(n_1107), .B1(n_1108), .B2(n_1109), .Y(n_1105) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_1106), .A2(n_1116), .B1(n_1117), .B2(n_1118), .Y(n_1115) );
OAI22xp5_ASAP7_75t_L g1166 ( .A1(n_1106), .A2(n_1167), .B1(n_1168), .B2(n_1169), .Y(n_1166) );
OAI22xp33_ASAP7_75t_L g1119 ( .A1(n_1108), .A2(n_1111), .B1(n_1120), .B2(n_1121), .Y(n_1119) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
NOR3xp33_ASAP7_75t_L g1263 ( .A(n_1123), .B(n_1264), .C(n_1278), .Y(n_1263) );
INVx1_ASAP7_75t_SL g1134 ( .A(n_1135), .Y(n_1134) );
AOI22xp5_ASAP7_75t_L g1143 ( .A1(n_1144), .A2(n_1299), .B1(n_1381), .B2(n_1382), .Y(n_1143) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1144), .Y(n_1381) );
XNOR2xp5_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1205), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
HB1xp67_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
XNOR2xp5_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1149), .Y(n_1147) );
NOR2x1_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1178), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1154), .Y(n_1150) );
OAI22xp5_ASAP7_75t_L g1157 ( .A1(n_1158), .A2(n_1159), .B1(n_1160), .B2(n_1161), .Y(n_1157) );
OAI211xp5_ASAP7_75t_L g1192 ( .A1(n_1163), .A2(n_1193), .B(n_1195), .C(n_1196), .Y(n_1192) );
OAI221xp5_ASAP7_75t_L g1648 ( .A1(n_1167), .A2(n_1649), .B1(n_1650), .B2(n_1651), .C(n_1652), .Y(n_1648) );
AOI22xp5_ASAP7_75t_L g1185 ( .A1(n_1175), .A2(n_1186), .B1(n_1187), .B2(n_1188), .Y(n_1185) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
NAND3xp33_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1197), .C(n_1201), .Y(n_1178) );
NOR3xp33_ASAP7_75t_SL g1179 ( .A(n_1180), .B(n_1189), .C(n_1191), .Y(n_1179) );
OAI21xp5_ASAP7_75t_SL g1180 ( .A1(n_1181), .A2(n_1183), .B(n_1185), .Y(n_1180) );
INVx2_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1199), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1201 ( .A(n_1202), .B(n_1203), .Y(n_1201) );
XNOR2xp5_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1261), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
HB1xp67_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
NAND3xp33_ASAP7_75t_L g1209 ( .A(n_1210), .B(n_1254), .C(n_1258), .Y(n_1209) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1211), .Y(n_1255) );
AOI22xp5_ASAP7_75t_L g1214 ( .A1(n_1215), .A2(n_1216), .B1(n_1217), .B2(n_1218), .Y(n_1214) );
AOI22xp5_ASAP7_75t_L g1219 ( .A1(n_1220), .A2(n_1228), .B1(n_1229), .B2(n_1230), .Y(n_1219) );
INVx3_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
BUFx6f_ASAP7_75t_L g1294 ( .A(n_1222), .Y(n_1294) );
INVx4_ASAP7_75t_L g1626 ( .A(n_1222), .Y(n_1626) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
AOI22xp5_ASAP7_75t_L g1624 ( .A1(n_1228), .A2(n_1229), .B1(n_1625), .B2(n_1630), .Y(n_1624) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1233), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1234), .B(n_1242), .Y(n_1233) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1244), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1248), .Y(n_1244) );
NAND2x1_ASAP7_75t_L g1245 ( .A(n_1246), .B(n_1247), .Y(n_1245) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1249), .Y(n_1259) );
AOI22xp5_ASAP7_75t_L g1643 ( .A1(n_1250), .A2(n_1252), .B1(n_1629), .B2(n_1644), .Y(n_1643) );
OAI21xp5_ASAP7_75t_L g1254 ( .A1(n_1255), .A2(n_1256), .B(n_1257), .Y(n_1254) );
OAI21xp33_ASAP7_75t_L g1258 ( .A1(n_1257), .A2(n_1259), .B(n_1260), .Y(n_1258) );
NAND3xp33_ASAP7_75t_L g1262 ( .A(n_1263), .B(n_1279), .C(n_1282), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1268), .Y(n_1264) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
OAI22xp5_ASAP7_75t_L g1375 ( .A1(n_1293), .A2(n_1376), .B1(n_1377), .B2(n_1378), .Y(n_1375) );
INVx2_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1299), .Y(n_1382) );
OAI22xp5_ASAP7_75t_L g1299 ( .A1(n_1300), .A2(n_1338), .B1(n_1339), .B2(n_1380), .Y(n_1299) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1300), .Y(n_1380) );
XNOR2x2_ASAP7_75t_L g1300 ( .A(n_1301), .B(n_1302), .Y(n_1300) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1325), .Y(n_1321) );
INVx2_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
XOR2x2_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1379), .Y(n_1339) );
NAND2xp5_ASAP7_75t_SL g1340 ( .A(n_1341), .B(n_1361), .Y(n_1340) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1344), .B(n_1351), .Y(n_1343) );
NOR2xp33_ASAP7_75t_L g1344 ( .A(n_1345), .B(n_1348), .Y(n_1344) );
NAND3xp33_ASAP7_75t_SL g1362 ( .A(n_1363), .B(n_1364), .C(n_1369), .Y(n_1362) );
BUFx4f_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
INVx3_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
OR2x2_ASAP7_75t_L g1385 ( .A(n_1386), .B(n_1392), .Y(n_1385) );
NOR2xp33_ASAP7_75t_L g1665 ( .A(n_1386), .B(n_1395), .Y(n_1665) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
NOR2xp33_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1390), .Y(n_1387) );
NOR2xp33_ASAP7_75t_L g1669 ( .A(n_1388), .B(n_1391), .Y(n_1669) );
INVx1_ASAP7_75t_L g1675 ( .A(n_1388), .Y(n_1675) );
HB1xp67_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
NOR2xp33_ASAP7_75t_L g1677 ( .A(n_1391), .B(n_1675), .Y(n_1677) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_1394), .B(n_1396), .Y(n_1393) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
AND2x4_ASAP7_75t_SL g1664 ( .A(n_1396), .B(n_1665), .Y(n_1664) );
INVx3_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
OAI221xp5_ASAP7_75t_L g1399 ( .A1(n_1400), .A2(n_1614), .B1(n_1617), .B2(n_1663), .C(n_1666), .Y(n_1399) );
AOI211xp5_ASAP7_75t_L g1400 ( .A1(n_1401), .A2(n_1526), .B(n_1530), .C(n_1589), .Y(n_1400) );
NAND5xp2_ASAP7_75t_L g1401 ( .A(n_1402), .B(n_1461), .C(n_1477), .D(n_1496), .E(n_1518), .Y(n_1401) );
AOI211xp5_ASAP7_75t_L g1402 ( .A1(n_1403), .A2(n_1433), .B(n_1442), .C(n_1454), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1404), .B(n_1418), .Y(n_1403) );
INVx2_ASAP7_75t_L g1452 ( .A(n_1404), .Y(n_1452) );
AND2x2_ASAP7_75t_L g1471 ( .A(n_1404), .B(n_1420), .Y(n_1471) );
AOI311xp33_ASAP7_75t_L g1496 ( .A1(n_1404), .A2(n_1497), .A3(n_1502), .B(n_1506), .C(n_1514), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1522 ( .A(n_1404), .B(n_1455), .Y(n_1522) );
OR2x2_ASAP7_75t_L g1548 ( .A(n_1404), .B(n_1549), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1568 ( .A(n_1404), .B(n_1429), .Y(n_1568) );
NAND2xp5_ASAP7_75t_L g1587 ( .A(n_1404), .B(n_1425), .Y(n_1587) );
OR2x2_ASAP7_75t_L g1604 ( .A(n_1404), .B(n_1425), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1405), .B(n_1413), .Y(n_1404) );
AND2x4_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1408), .Y(n_1406) );
AND2x6_ASAP7_75t_L g1411 ( .A(n_1407), .B(n_1412), .Y(n_1411) );
AND2x6_ASAP7_75t_L g1414 ( .A(n_1407), .B(n_1415), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_1407), .B(n_1417), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_1407), .B(n_1417), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1528 ( .A(n_1407), .B(n_1417), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1409), .B(n_1410), .Y(n_1408) );
INVx2_ASAP7_75t_L g1616 ( .A(n_1414), .Y(n_1616) );
OAI21xp5_ASAP7_75t_L g1674 ( .A1(n_1415), .A2(n_1675), .B(n_1676), .Y(n_1674) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1419), .B(n_1423), .Y(n_1418) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1419), .Y(n_1450) );
NAND2xp5_ASAP7_75t_L g1503 ( .A(n_1419), .B(n_1504), .Y(n_1503) );
OR2x2_ASAP7_75t_L g1515 ( .A(n_1419), .B(n_1459), .Y(n_1515) );
OAI21xp33_ASAP7_75t_L g1536 ( .A1(n_1419), .A2(n_1537), .B(n_1538), .Y(n_1536) );
OAI332xp33_ASAP7_75t_L g1581 ( .A1(n_1419), .A2(n_1522), .A3(n_1582), .B1(n_1584), .B2(n_1585), .B3(n_1586), .C1(n_1587), .C2(n_1588), .Y(n_1581) );
OR2x2_ASAP7_75t_L g1582 ( .A(n_1419), .B(n_1583), .Y(n_1582) );
CKINVDCx5p33_ASAP7_75t_R g1419 ( .A(n_1420), .Y(n_1419) );
NOR2xp33_ASAP7_75t_L g1480 ( .A(n_1420), .B(n_1481), .Y(n_1480) );
INVx3_ASAP7_75t_L g1485 ( .A(n_1420), .Y(n_1485) );
AND2x2_ASAP7_75t_L g1519 ( .A(n_1420), .B(n_1513), .Y(n_1519) );
NOR2xp33_ASAP7_75t_L g1545 ( .A(n_1420), .B(n_1488), .Y(n_1545) );
NAND2xp5_ASAP7_75t_L g1549 ( .A(n_1420), .B(n_1423), .Y(n_1549) );
OR2x2_ASAP7_75t_L g1603 ( .A(n_1420), .B(n_1604), .Y(n_1603) );
AND2x4_ASAP7_75t_SL g1420 ( .A(n_1421), .B(n_1422), .Y(n_1420) );
NAND2xp5_ASAP7_75t_L g1601 ( .A(n_1423), .B(n_1471), .Y(n_1601) );
AND2x2_ASAP7_75t_L g1423 ( .A(n_1424), .B(n_1429), .Y(n_1423) );
OR2x2_ASAP7_75t_L g1455 ( .A(n_1424), .B(n_1430), .Y(n_1455) );
AOI322xp5_ASAP7_75t_L g1518 ( .A1(n_1424), .A2(n_1504), .A3(n_1519), .B1(n_1520), .B2(n_1521), .C1(n_1523), .C2(n_1525), .Y(n_1518) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1425), .B(n_1430), .Y(n_1453) );
NOR2xp33_ASAP7_75t_L g1469 ( .A(n_1425), .B(n_1470), .Y(n_1469) );
OR2x2_ASAP7_75t_L g1488 ( .A(n_1425), .B(n_1489), .Y(n_1488) );
AND2x2_ASAP7_75t_L g1540 ( .A(n_1425), .B(n_1452), .Y(n_1540) );
NOR3xp33_ASAP7_75t_SL g1574 ( .A(n_1425), .B(n_1450), .C(n_1526), .Y(n_1574) );
AND2x2_ASAP7_75t_L g1425 ( .A(n_1426), .B(n_1427), .Y(n_1425) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1430), .Y(n_1483) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1430), .Y(n_1489) );
NAND2xp5_ASAP7_75t_L g1583 ( .A(n_1430), .B(n_1452), .Y(n_1583) );
NAND2x1_ASAP7_75t_L g1430 ( .A(n_1431), .B(n_1432), .Y(n_1430) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1433), .Y(n_1566) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1434), .B(n_1438), .Y(n_1433) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1435), .Y(n_1457) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1435), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1474 ( .A(n_1435), .B(n_1438), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_1435), .B(n_1439), .Y(n_1479) );
NAND2xp5_ASAP7_75t_L g1435 ( .A(n_1436), .B(n_1437), .Y(n_1435) );
OR2x2_ASAP7_75t_L g1492 ( .A(n_1438), .B(n_1444), .Y(n_1492) );
NAND2xp5_ASAP7_75t_L g1505 ( .A(n_1438), .B(n_1445), .Y(n_1505) );
HB1xp67_ASAP7_75t_SL g1554 ( .A(n_1438), .Y(n_1554) );
NAND2xp5_ASAP7_75t_L g1586 ( .A(n_1438), .B(n_1543), .Y(n_1586) );
CKINVDCx5p33_ASAP7_75t_R g1438 ( .A(n_1439), .Y(n_1438) );
NAND2xp5_ASAP7_75t_L g1459 ( .A(n_1439), .B(n_1460), .Y(n_1459) );
OR2x2_ASAP7_75t_L g1464 ( .A(n_1439), .B(n_1445), .Y(n_1464) );
HB1xp67_ASAP7_75t_SL g1490 ( .A(n_1439), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1525 ( .A(n_1439), .B(n_1457), .Y(n_1525) );
AND2x4_ASAP7_75t_L g1439 ( .A(n_1440), .B(n_1441), .Y(n_1439) );
NOR2xp33_ASAP7_75t_L g1442 ( .A(n_1443), .B(n_1448), .Y(n_1442) );
OAI32xp33_ASAP7_75t_L g1578 ( .A1(n_1443), .A2(n_1444), .A3(n_1508), .B1(n_1538), .B2(n_1579), .Y(n_1578) );
NAND2xp5_ASAP7_75t_L g1588 ( .A(n_1443), .B(n_1474), .Y(n_1588) );
INVx2_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1555 ( .A(n_1444), .B(n_1524), .Y(n_1555) );
NAND2xp5_ASAP7_75t_L g1594 ( .A(n_1444), .B(n_1561), .Y(n_1594) );
INVx2_ASAP7_75t_SL g1444 ( .A(n_1445), .Y(n_1444) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1445), .Y(n_1460) );
AND2x2_ASAP7_75t_L g1569 ( .A(n_1445), .B(n_1485), .Y(n_1569) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1446), .B(n_1447), .Y(n_1445) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
O2A1O1Ixp33_ASAP7_75t_L g1544 ( .A1(n_1449), .A2(n_1545), .B(n_1546), .C(n_1547), .Y(n_1544) );
AND2x2_ASAP7_75t_L g1449 ( .A(n_1450), .B(n_1451), .Y(n_1449) );
OR2x2_ASAP7_75t_L g1475 ( .A(n_1450), .B(n_1476), .Y(n_1475) );
AOI221xp5_ASAP7_75t_L g1461 ( .A1(n_1451), .A2(n_1462), .B1(n_1465), .B2(n_1469), .C(n_1472), .Y(n_1461) );
AND2x2_ASAP7_75t_L g1451 ( .A(n_1452), .B(n_1453), .Y(n_1451) );
OR2x2_ASAP7_75t_L g1476 ( .A(n_1452), .B(n_1455), .Y(n_1476) );
AND2x2_ASAP7_75t_L g1482 ( .A(n_1452), .B(n_1483), .Y(n_1482) );
OR2x2_ASAP7_75t_L g1487 ( .A(n_1452), .B(n_1488), .Y(n_1487) );
NAND2xp5_ASAP7_75t_L g1495 ( .A(n_1452), .B(n_1485), .Y(n_1495) );
OR2x2_ASAP7_75t_L g1533 ( .A(n_1452), .B(n_1534), .Y(n_1533) );
AND2x2_ASAP7_75t_L g1538 ( .A(n_1452), .B(n_1501), .Y(n_1538) );
OR2x2_ASAP7_75t_L g1597 ( .A(n_1452), .B(n_1494), .Y(n_1597) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1453), .Y(n_1494) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1453), .B(n_1471), .Y(n_1524) );
NAND2xp5_ASAP7_75t_L g1534 ( .A(n_1453), .B(n_1485), .Y(n_1534) );
NOR2xp33_ASAP7_75t_L g1454 ( .A(n_1455), .B(n_1456), .Y(n_1454) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1455), .Y(n_1500) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1456), .Y(n_1546) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_1457), .B(n_1458), .Y(n_1456) );
AND2x2_ASAP7_75t_L g1462 ( .A(n_1457), .B(n_1463), .Y(n_1462) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1457), .Y(n_1513) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1457), .Y(n_1552) );
AND2x2_ASAP7_75t_L g1610 ( .A(n_1457), .B(n_1512), .Y(n_1610) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1459), .Y(n_1537) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1459), .Y(n_1609) );
AND2x2_ASAP7_75t_L g1478 ( .A(n_1460), .B(n_1479), .Y(n_1478) );
INVx2_ASAP7_75t_L g1512 ( .A(n_1460), .Y(n_1512) );
NAND2xp5_ASAP7_75t_L g1466 ( .A(n_1463), .B(n_1467), .Y(n_1466) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_1463), .B(n_1485), .Y(n_1577) );
INVx2_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
NOR2xp33_ASAP7_75t_L g1612 ( .A(n_1464), .B(n_1485), .Y(n_1612) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
OAI332xp33_ASAP7_75t_L g1563 ( .A1(n_1468), .A2(n_1503), .A3(n_1549), .B1(n_1564), .B2(n_1565), .B3(n_1566), .C1(n_1567), .C2(n_1570), .Y(n_1563) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
AND2x2_ASAP7_75t_L g1508 ( .A(n_1471), .B(n_1501), .Y(n_1508) );
NOR2xp33_ASAP7_75t_L g1472 ( .A(n_1473), .B(n_1475), .Y(n_1472) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
AOI21xp33_ASAP7_75t_L g1514 ( .A1(n_1476), .A2(n_1515), .B(n_1516), .Y(n_1514) );
INVx2_ASAP7_75t_L g1559 ( .A(n_1476), .Y(n_1559) );
AOI221xp5_ASAP7_75t_L g1477 ( .A1(n_1478), .A2(n_1480), .B1(n_1484), .B2(n_1490), .C(n_1491), .Y(n_1477) );
OAI31xp33_ASAP7_75t_L g1590 ( .A1(n_1479), .A2(n_1532), .A3(n_1591), .B(n_1593), .Y(n_1590) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
A2O1A1Ixp33_ASAP7_75t_L g1611 ( .A1(n_1483), .A2(n_1571), .B(n_1612), .C(n_1613), .Y(n_1611) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1485), .B(n_1486), .Y(n_1484) );
NOR2xp33_ASAP7_75t_L g1541 ( .A(n_1485), .B(n_1492), .Y(n_1541) );
CKINVDCx14_ASAP7_75t_R g1558 ( .A(n_1485), .Y(n_1558) );
NAND2xp5_ASAP7_75t_L g1592 ( .A(n_1486), .B(n_1512), .Y(n_1592) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
INVx1_ASAP7_75t_L g1501 ( .A(n_1488), .Y(n_1501) );
A2O1A1Ixp33_ASAP7_75t_L g1531 ( .A1(n_1490), .A2(n_1532), .B(n_1535), .C(n_1543), .Y(n_1531) );
NOR2xp33_ASAP7_75t_L g1491 ( .A(n_1492), .B(n_1493), .Y(n_1491) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1492), .Y(n_1520) );
OAI22xp33_ASAP7_75t_L g1600 ( .A1(n_1492), .A2(n_1509), .B1(n_1516), .B2(n_1601), .Y(n_1600) );
OR2x2_ASAP7_75t_L g1493 ( .A(n_1494), .B(n_1495), .Y(n_1493) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1495), .Y(n_1510) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1499), .Y(n_1498) );
NOR2xp33_ASAP7_75t_L g1499 ( .A(n_1500), .B(n_1501), .Y(n_1499) );
NAND2xp5_ASAP7_75t_L g1509 ( .A(n_1500), .B(n_1510), .Y(n_1509) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1503), .Y(n_1502) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1504), .Y(n_1562) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
OR2x2_ASAP7_75t_L g1551 ( .A(n_1505), .B(n_1552), .Y(n_1551) );
AOI21xp5_ASAP7_75t_L g1506 ( .A1(n_1507), .A2(n_1509), .B(n_1511), .Y(n_1506) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1508), .Y(n_1507) );
OAI22xp5_ASAP7_75t_L g1547 ( .A1(n_1511), .A2(n_1548), .B1(n_1550), .B2(n_1551), .Y(n_1547) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1511), .Y(n_1598) );
OR2x2_ASAP7_75t_L g1511 ( .A(n_1512), .B(n_1513), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_1512), .B(n_1513), .Y(n_1517) );
AND2x2_ASAP7_75t_L g1523 ( .A(n_1512), .B(n_1524), .Y(n_1523) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1512), .Y(n_1585) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
NAND2xp5_ASAP7_75t_L g1542 ( .A(n_1520), .B(n_1521), .Y(n_1542) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
NOR2xp33_ASAP7_75t_SL g1570 ( .A(n_1525), .B(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1525), .Y(n_1605) );
INVx3_ASAP7_75t_L g1543 ( .A(n_1526), .Y(n_1543) );
NOR2xp33_ASAP7_75t_L g1571 ( .A(n_1526), .B(n_1552), .Y(n_1571) );
NOR3xp33_ASAP7_75t_L g1602 ( .A(n_1526), .B(n_1603), .C(n_1605), .Y(n_1602) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1527), .B(n_1529), .Y(n_1526) );
NAND4xp25_ASAP7_75t_L g1530 ( .A(n_1531), .B(n_1544), .C(n_1553), .D(n_1572), .Y(n_1530) );
AOI22xp5_ASAP7_75t_L g1606 ( .A1(n_1532), .A2(n_1561), .B1(n_1607), .B2(n_1610), .Y(n_1606) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1534), .Y(n_1579) );
NAND3xp33_ASAP7_75t_SL g1535 ( .A(n_1536), .B(n_1539), .C(n_1542), .Y(n_1535) );
INVx2_ASAP7_75t_L g1550 ( .A(n_1538), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1561 ( .A(n_1538), .B(n_1558), .Y(n_1561) );
NAND2xp5_ASAP7_75t_L g1539 ( .A(n_1540), .B(n_1541), .Y(n_1539) );
CKINVDCx14_ASAP7_75t_R g1564 ( .A(n_1540), .Y(n_1564) );
CKINVDCx14_ASAP7_75t_R g1565 ( .A(n_1543), .Y(n_1565) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1543), .B(n_1552), .Y(n_1580) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1551), .Y(n_1573) );
NAND2xp5_ASAP7_75t_L g1607 ( .A(n_1551), .B(n_1608), .Y(n_1607) );
AOI211xp5_ASAP7_75t_L g1553 ( .A1(n_1554), .A2(n_1555), .B(n_1556), .C(n_1563), .Y(n_1553) );
AOI21xp33_ASAP7_75t_L g1556 ( .A1(n_1557), .A2(n_1560), .B(n_1562), .Y(n_1556) );
NAND2xp5_ASAP7_75t_L g1557 ( .A(n_1558), .B(n_1559), .Y(n_1557) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
CKINVDCx14_ASAP7_75t_R g1599 ( .A(n_1565), .Y(n_1599) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_1568), .B(n_1569), .Y(n_1567) );
OAI21xp5_ASAP7_75t_L g1575 ( .A1(n_1568), .A2(n_1576), .B(n_1578), .Y(n_1575) );
INVxp67_ASAP7_75t_SL g1584 ( .A(n_1571), .Y(n_1584) );
AOI221xp5_ASAP7_75t_L g1572 ( .A1(n_1573), .A2(n_1574), .B1(n_1575), .B2(n_1580), .C(n_1581), .Y(n_1572) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1577), .Y(n_1576) );
NAND4xp25_ASAP7_75t_L g1589 ( .A(n_1590), .B(n_1595), .C(n_1606), .D(n_1611), .Y(n_1589) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1594), .Y(n_1593) );
AOI311xp33_ASAP7_75t_L g1595 ( .A1(n_1596), .A2(n_1598), .A3(n_1599), .B(n_1600), .C(n_1602), .Y(n_1595) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1601), .Y(n_1613) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1609), .Y(n_1608) );
CKINVDCx20_ASAP7_75t_R g1614 ( .A(n_1615), .Y(n_1614) );
CKINVDCx20_ASAP7_75t_R g1615 ( .A(n_1616), .Y(n_1615) );
INVx2_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
HB1xp67_ASAP7_75t_L g1672 ( .A(n_1619), .Y(n_1672) );
AOI21xp5_ASAP7_75t_L g1620 ( .A1(n_1621), .A2(n_1641), .B(n_1642), .Y(n_1620) );
NAND4xp25_ASAP7_75t_L g1621 ( .A(n_1622), .B(n_1624), .C(n_1633), .D(n_1637), .Y(n_1621) );
OAI22xp5_ASAP7_75t_SL g1646 ( .A1(n_1647), .A2(n_1648), .B1(n_1653), .B2(n_1654), .Y(n_1646) );
NAND2xp5_ASAP7_75t_L g1658 ( .A(n_1659), .B(n_1660), .Y(n_1658) );
INVx2_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
HB1xp67_ASAP7_75t_SL g1667 ( .A(n_1668), .Y(n_1667) );
BUFx3_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
INVxp33_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
HB1xp67_ASAP7_75t_L g1673 ( .A(n_1674), .Y(n_1673) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1677), .Y(n_1676) );
endmodule