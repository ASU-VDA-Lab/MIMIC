module fake_jpeg_183_n_704 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_704);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_704;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_61),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_62),
.Y(n_180)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_64),
.Y(n_162)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_67),
.Y(n_167)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_68),
.Y(n_144)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_70),
.B(n_74),
.Y(n_137)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_71),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_73),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_9),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_77),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_25),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_78),
.A2(n_114),
.B(n_16),
.Y(n_173)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_79),
.Y(n_184)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_81),
.Y(n_194)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_25),
.B(n_9),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_83),
.A2(n_101),
.B(n_109),
.C(n_112),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_38),
.B(n_9),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_84),
.B(n_100),
.Y(n_140)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

INVxp67_ASAP7_75t_SL g87 ( 
.A(n_47),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_89),
.Y(n_195)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_92),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_93),
.Y(n_212)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_94),
.Y(n_175)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_95),
.Y(n_166)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_96),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_98),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

NOR2xp67_ASAP7_75t_L g100 ( 
.A(n_35),
.B(n_8),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_35),
.B(n_8),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g155 ( 
.A(n_102),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_103),
.Y(n_200)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g186 ( 
.A(n_105),
.Y(n_186)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_108),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_35),
.B(n_10),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_34),
.B(n_53),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_21),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_113),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_34),
.B(n_10),
.Y(n_114)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_30),
.Y(n_115)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_45),
.Y(n_116)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_38),
.Y(n_117)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_118),
.Y(n_171)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_120),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_21),
.Y(n_121)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_121),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_37),
.Y(n_123)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_21),
.Y(n_124)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_124),
.Y(n_213)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_37),
.Y(n_125)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_125),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_28),
.Y(n_126)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_30),
.Y(n_127)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_127),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_30),
.Y(n_128)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_128),
.Y(n_226)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_37),
.Y(n_129)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_46),
.Y(n_130)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_130),
.Y(n_206)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_33),
.Y(n_131)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_131),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g132 ( 
.A(n_46),
.Y(n_132)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_132),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_78),
.A2(n_27),
.B1(n_36),
.B2(n_56),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_138),
.A2(n_141),
.B1(n_142),
.B2(n_149),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_72),
.A2(n_27),
.B1(n_36),
.B2(n_56),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_74),
.A2(n_84),
.B1(n_124),
.B2(n_121),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_49),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_146),
.B(n_172),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_49),
.B1(n_53),
.B2(n_50),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_83),
.A2(n_50),
.B1(n_43),
.B2(n_60),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_157),
.A2(n_160),
.B1(n_163),
.B2(n_208),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_L g160 ( 
.A1(n_68),
.A2(n_60),
.B1(n_43),
.B2(n_42),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_101),
.B(n_51),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_161),
.B(n_191),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_113),
.A2(n_42),
.B1(n_59),
.B2(n_44),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_109),
.B(n_51),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_173),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_51),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_183),
.B(n_187),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_88),
.B(n_44),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_87),
.B(n_39),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_190),
.B(n_0),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_65),
.B(n_44),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_94),
.A2(n_60),
.B1(n_43),
.B2(n_42),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g230 ( 
.A1(n_193),
.A2(n_222),
.B1(n_223),
.B2(n_62),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_127),
.B(n_39),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_201),
.B(n_203),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_128),
.B(n_59),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_89),
.B(n_59),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_204),
.B(n_207),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_96),
.B(n_52),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_102),
.A2(n_92),
.B1(n_111),
.B2(n_105),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_73),
.A2(n_52),
.B1(n_39),
.B2(n_29),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_209),
.A2(n_215),
.B1(n_0),
.B2(n_1),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_93),
.B(n_52),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_214),
.B(n_216),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_97),
.A2(n_54),
.B1(n_32),
.B2(n_31),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_98),
.B(n_32),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_99),
.A2(n_54),
.B1(n_32),
.B2(n_31),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_103),
.A2(n_54),
.B1(n_31),
.B2(n_29),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_132),
.B(n_29),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_0),
.Y(n_245)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_145),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_227),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_141),
.A2(n_28),
.B1(n_33),
.B2(n_46),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_228),
.A2(n_278),
.B1(n_279),
.B2(n_181),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_230),
.A2(n_271),
.B1(n_286),
.B2(n_289),
.Y(n_335)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

INVx4_ASAP7_75t_SL g308 ( 
.A(n_232),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_33),
.C(n_46),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_233),
.B(n_261),
.Y(n_311)
);

INVx11_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_234),
.Y(n_316)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

BUFx4f_ASAP7_75t_SL g329 ( 
.A(n_235),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_173),
.B(n_0),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_236),
.B(n_283),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_237),
.Y(n_312)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_176),
.Y(n_239)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_239),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_240),
.B(n_252),
.Y(n_309)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_180),
.Y(n_241)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_241),
.Y(n_330)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_165),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_242),
.Y(n_350)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_243),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_196),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_244),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_245),
.B(n_246),
.Y(n_334)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_168),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_247),
.B(n_258),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_145),
.Y(n_248)
);

INVx6_ASAP7_75t_L g331 ( 
.A(n_248),
.Y(n_331)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_185),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_250),
.Y(n_370)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_155),
.Y(n_251)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_251),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_140),
.B(n_7),
.Y(n_252)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_182),
.Y(n_253)
);

INVx5_ASAP7_75t_L g342 ( 
.A(n_253),
.Y(n_342)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_169),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_254),
.B(n_255),
.Y(n_340)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_162),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_155),
.Y(n_256)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_256),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_150),
.Y(n_258)
);

INVx11_ASAP7_75t_L g259 ( 
.A(n_180),
.Y(n_259)
);

INVx11_ASAP7_75t_L g359 ( 
.A(n_259),
.Y(n_359)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_219),
.Y(n_260)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_260),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_139),
.Y(n_261)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_199),
.Y(n_262)
);

INVx5_ASAP7_75t_L g349 ( 
.A(n_262),
.Y(n_349)
);

BUFx6f_ASAP7_75t_SL g264 ( 
.A(n_211),
.Y(n_264)
);

INVx13_ASAP7_75t_L g352 ( 
.A(n_264),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_182),
.Y(n_265)
);

INVx5_ASAP7_75t_L g367 ( 
.A(n_265),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_197),
.A2(n_46),
.B1(n_7),
.B2(n_11),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_266),
.A2(n_267),
.B1(n_285),
.B2(n_300),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_138),
.A2(n_6),
.B1(n_17),
.B2(n_14),
.Y(n_267)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_205),
.Y(n_268)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_178),
.Y(n_270)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_270),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_137),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_220),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_272),
.B(n_274),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_167),
.B(n_14),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_273),
.B(n_144),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_150),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_185),
.Y(n_275)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_275),
.Y(n_336)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_164),
.A2(n_18),
.B1(n_14),
.B2(n_13),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_276),
.A2(n_303),
.B1(n_212),
.B2(n_218),
.Y(n_362)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_154),
.Y(n_277)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_277),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_222),
.A2(n_18),
.B1(n_12),
.B2(n_7),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_158),
.Y(n_280)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_280),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_205),
.Y(n_281)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_281),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_139),
.B(n_12),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_282),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_133),
.B(n_1),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_186),
.Y(n_284)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_284),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_160),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_152),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_286)
);

HAxp5_ASAP7_75t_SL g287 ( 
.A(n_223),
.B(n_1),
.CON(n_287),
.SN(n_287)
);

NOR2x1_ASAP7_75t_L g320 ( 
.A(n_287),
.B(n_202),
.Y(n_320)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_226),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_298),
.Y(n_318)
);

INVx8_ASAP7_75t_L g289 ( 
.A(n_199),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_179),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_290),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_136),
.A2(n_2),
.B(n_4),
.C(n_5),
.Y(n_291)
);

A2O1A1Ixp33_ASAP7_75t_L g322 ( 
.A1(n_291),
.A2(n_156),
.B(n_199),
.C(n_170),
.Y(n_322)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_166),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_292),
.B(n_297),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_153),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_293),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_147),
.B(n_4),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_294),
.B(n_148),
.Y(n_333)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_177),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_194),
.Y(n_298)
);

BUFx4f_ASAP7_75t_L g299 ( 
.A(n_152),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_299),
.A2(n_301),
.B1(n_302),
.B2(n_159),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_188),
.A2(n_186),
.B1(n_210),
.B2(n_213),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_135),
.A2(n_4),
.B1(n_5),
.B2(n_151),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_143),
.A2(n_5),
.B1(n_217),
.B2(n_174),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_193),
.A2(n_134),
.B1(n_184),
.B2(n_171),
.Y(n_303)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_194),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_304),
.Y(n_360)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_192),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_156),
.Y(n_328)
);

INVx13_ASAP7_75t_L g306 ( 
.A(n_206),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_206),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_236),
.B(n_171),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_317),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_320),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_322),
.A2(n_323),
.B(n_291),
.Y(n_376)
);

NOR2x1_ASAP7_75t_L g323 ( 
.A(n_249),
.B(n_218),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_328),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_333),
.B(n_351),
.Y(n_373)
);

INVxp33_ASAP7_75t_L g401 ( 
.A(n_337),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_269),
.A2(n_134),
.B1(n_184),
.B2(n_212),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_338),
.A2(n_366),
.B1(n_308),
.B2(n_315),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_307),
.B(n_238),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_345),
.B(n_346),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_231),
.B(n_148),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_263),
.B(n_170),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_347),
.B(n_348),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_295),
.B(n_144),
.Y(n_348)
);

AO22x2_ASAP7_75t_L g353 ( 
.A1(n_228),
.A2(n_159),
.B1(n_181),
.B2(n_189),
.Y(n_353)
);

O2A1O1Ixp33_ASAP7_75t_SL g392 ( 
.A1(n_353),
.A2(n_227),
.B(n_281),
.C(n_265),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_296),
.B(n_195),
.Y(n_354)
);

BUFx24_ASAP7_75t_SL g407 ( 
.A(n_354),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_257),
.B(n_195),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_358),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_272),
.B(n_237),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_362),
.B(n_365),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_364),
.A2(n_259),
.B1(n_234),
.B2(n_235),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_261),
.B(n_189),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_368),
.B(n_284),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_323),
.A2(n_299),
.B1(n_230),
.B2(n_264),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_371),
.A2(n_379),
.B1(n_388),
.B2(n_396),
.Y(n_447)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_308),
.Y(n_372)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_372),
.Y(n_421)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_341),
.Y(n_374)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_341),
.Y(n_375)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_375),
.Y(n_422)
);

O2A1O1Ixp33_ASAP7_75t_L g430 ( 
.A1(n_376),
.A2(n_412),
.B(n_393),
.C(n_389),
.Y(n_430)
);

AO22x1_ASAP7_75t_L g377 ( 
.A1(n_322),
.A2(n_287),
.B1(n_230),
.B2(n_299),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_377),
.B(n_403),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_323),
.A2(n_230),
.B1(n_232),
.B2(n_270),
.Y(n_379)
);

NAND2x1_ASAP7_75t_L g380 ( 
.A(n_311),
.B(n_282),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_380),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_355),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_381),
.Y(n_453)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_356),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_382),
.B(n_383),
.Y(n_435)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_356),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_365),
.A2(n_294),
.B1(n_283),
.B2(n_200),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_384),
.A2(n_385),
.B1(n_411),
.B2(n_413),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_335),
.A2(n_200),
.B1(n_268),
.B2(n_253),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_321),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_387),
.B(n_390),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_343),
.A2(n_256),
.B1(n_251),
.B2(n_290),
.Y(n_388)
);

AND2x2_ASAP7_75t_SL g391 ( 
.A(n_311),
.B(n_233),
.Y(n_391)
);

MAJx2_ASAP7_75t_L g424 ( 
.A(n_391),
.B(n_337),
.C(n_318),
.Y(n_424)
);

AO21x2_ASAP7_75t_L g440 ( 
.A1(n_392),
.A2(n_336),
.B(n_363),
.Y(n_440)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_369),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_394),
.B(n_399),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_311),
.B(n_229),
.C(n_242),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_395),
.B(n_402),
.C(n_408),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_317),
.A2(n_357),
.B1(n_310),
.B2(n_313),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_397),
.A2(n_418),
.B(n_349),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_317),
.A2(n_248),
.B1(n_229),
.B2(n_260),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_398),
.A2(n_400),
.B1(n_404),
.B2(n_312),
.Y(n_454)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_310),
.A2(n_288),
.B1(n_275),
.B2(n_250),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_333),
.B(n_298),
.C(n_239),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_324),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_313),
.A2(n_304),
.B1(n_243),
.B2(n_262),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_324),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_405),
.B(n_416),
.Y(n_450)
);

BUFx8_ASAP7_75t_L g406 ( 
.A(n_359),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_406),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_320),
.B(n_334),
.C(n_340),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_320),
.B(n_241),
.Y(n_409)
);

XOR2x1_ASAP7_75t_L g455 ( 
.A(n_409),
.B(n_359),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_340),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_410),
.B(n_378),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_362),
.A2(n_289),
.B1(n_244),
.B2(n_306),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_353),
.A2(n_334),
.B1(n_351),
.B2(n_344),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_415),
.A2(n_326),
.B1(n_332),
.B2(n_350),
.Y(n_432)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_314),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_308),
.A2(n_360),
.B1(n_326),
.B2(n_318),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_325),
.B(n_344),
.C(n_361),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_419),
.B(n_387),
.C(n_395),
.Y(n_452)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_314),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_420),
.B(n_312),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_423),
.B(n_459),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_424),
.B(n_458),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_393),
.A2(n_316),
.B(n_360),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_425),
.A2(n_434),
.B(n_430),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_386),
.A2(n_353),
.B1(n_315),
.B2(n_366),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_426),
.A2(n_432),
.B1(n_433),
.B2(n_446),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_430),
.A2(n_455),
.B(n_383),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_391),
.B(n_361),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_431),
.B(n_436),
.C(n_457),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_386),
.A2(n_353),
.B1(n_342),
.B2(n_331),
.Y(n_433)
);

AOI211xp5_ASAP7_75t_SL g434 ( 
.A1(n_377),
.A2(n_353),
.B(n_318),
.C(n_309),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_391),
.B(n_419),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_412),
.A2(n_309),
.B(n_337),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_437),
.A2(n_449),
.B(n_451),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_438),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_386),
.A2(n_336),
.B1(n_342),
.B2(n_367),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_439),
.A2(n_444),
.B1(n_404),
.B2(n_372),
.Y(n_467)
);

OA22x2_ASAP7_75t_L g475 ( 
.A1(n_440),
.A2(n_442),
.B1(n_392),
.B2(n_398),
.Y(n_475)
);

OA22x2_ASAP7_75t_L g442 ( 
.A1(n_392),
.A2(n_332),
.B1(n_363),
.B2(n_367),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_413),
.A2(n_355),
.B1(n_350),
.B2(n_319),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_396),
.A2(n_331),
.B1(n_355),
.B2(n_350),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_409),
.A2(n_319),
.B(n_339),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_409),
.A2(n_312),
.B(n_330),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_452),
.B(n_374),
.Y(n_492)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_454),
.Y(n_465)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_456),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_408),
.B(n_339),
.C(n_330),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_380),
.B(n_329),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_410),
.B(n_370),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_373),
.B(n_329),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_461),
.B(n_390),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_376),
.A2(n_370),
.B1(n_349),
.B2(n_327),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_462),
.A2(n_385),
.B1(n_411),
.B2(n_389),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_460),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_463),
.B(n_494),
.Y(n_506)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_467),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_427),
.A2(n_373),
.B1(n_377),
.B2(n_414),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_469),
.A2(n_478),
.B1(n_482),
.B2(n_493),
.Y(n_510)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_470),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_428),
.B(n_384),
.Y(n_472)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_472),
.Y(n_507)
);

BUFx24_ASAP7_75t_SL g473 ( 
.A(n_423),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_473),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_428),
.B(n_407),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_474),
.B(n_476),
.Y(n_522)
);

OA21x2_ASAP7_75t_L g515 ( 
.A1(n_475),
.A2(n_442),
.B(n_426),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_417),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_462),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_477),
.Y(n_533)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_435),
.Y(n_480)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_480),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_447),
.A2(n_448),
.B1(n_429),
.B2(n_461),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_481),
.A2(n_484),
.B(n_487),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_427),
.A2(n_400),
.B1(n_417),
.B2(n_401),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_435),
.Y(n_483)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_483),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_447),
.A2(n_448),
.B1(n_429),
.B2(n_433),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_436),
.B(n_402),
.C(n_380),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_485),
.B(n_492),
.C(n_501),
.Y(n_509)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_460),
.Y(n_486)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_486),
.Y(n_523)
);

INVxp67_ASAP7_75t_R g488 ( 
.A(n_437),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_488),
.B(n_500),
.Y(n_531)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_450),
.Y(n_490)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_490),
.Y(n_537)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_450),
.Y(n_491)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_491),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_440),
.A2(n_415),
.B1(n_375),
.B2(n_382),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_422),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_422),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_495),
.B(n_499),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_440),
.A2(n_399),
.B1(n_394),
.B2(n_403),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_497),
.A2(n_454),
.B1(n_446),
.B2(n_445),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_498),
.A2(n_458),
.B(n_424),
.Y(n_526)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_445),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_459),
.B(n_327),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_431),
.B(n_405),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_480),
.Y(n_503)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_503),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_498),
.A2(n_425),
.B(n_451),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_504),
.A2(n_517),
.B(n_539),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_496),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_511),
.B(n_520),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_484),
.A2(n_440),
.B1(n_444),
.B2(n_434),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_513),
.A2(n_465),
.B1(n_477),
.B2(n_482),
.Y(n_541)
);

CKINVDCx14_ASAP7_75t_R g514 ( 
.A(n_470),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_514),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_515),
.A2(n_475),
.B1(n_488),
.B2(n_464),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_487),
.A2(n_438),
.B(n_449),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_479),
.A2(n_440),
.B(n_455),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_518),
.A2(n_526),
.B(n_535),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_466),
.B(n_441),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_519),
.B(n_524),
.C(n_525),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_497),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_493),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_521),
.B(n_534),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_466),
.B(n_441),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_492),
.B(n_424),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_485),
.B(n_457),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_527),
.B(n_475),
.C(n_416),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_529),
.A2(n_478),
.B1(n_468),
.B2(n_465),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_463),
.B(n_421),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_530),
.B(n_483),
.Y(n_547)
);

AO22x1_ASAP7_75t_L g534 ( 
.A1(n_469),
.A2(n_440),
.B1(n_442),
.B2(n_421),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_479),
.A2(n_439),
.B(n_442),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_499),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_536),
.B(n_471),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_489),
.A2(n_442),
.B(n_456),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_541),
.A2(n_543),
.B1(n_552),
.B2(n_554),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_542),
.A2(n_561),
.B1(n_515),
.B2(n_510),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_534),
.A2(n_491),
.B1(n_490),
.B2(n_468),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_506),
.Y(n_544)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_544),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_547),
.B(n_549),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_511),
.B(n_486),
.Y(n_549)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_551),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_508),
.B(n_474),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_506),
.Y(n_553)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_553),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_534),
.A2(n_471),
.B1(n_472),
.B2(n_467),
.Y(n_554)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_528),
.Y(n_556)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_556),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_521),
.A2(n_475),
.B1(n_481),
.B2(n_464),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_557),
.A2(n_567),
.B1(n_569),
.B2(n_535),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_528),
.B(n_495),
.Y(n_558)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_558),
.Y(n_586)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_530),
.Y(n_559)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_559),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_531),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_560),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_539),
.A2(n_489),
.B(n_501),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_562),
.A2(n_566),
.B(n_574),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_508),
.B(n_494),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_563),
.B(n_565),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_564),
.B(n_509),
.C(n_527),
.Y(n_589)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_512),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_539),
.A2(n_432),
.B(n_443),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_513),
.A2(n_443),
.B1(n_453),
.B2(n_406),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_533),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_568),
.B(n_571),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_515),
.A2(n_453),
.B1(n_381),
.B2(n_406),
.Y(n_569)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_512),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_523),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_572),
.B(n_573),
.Y(n_602)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_523),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_516),
.A2(n_504),
.B(n_518),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_575),
.A2(n_587),
.B1(n_594),
.B2(n_603),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_552),
.B(n_522),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_577),
.B(n_584),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_564),
.B(n_519),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_578),
.B(n_589),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_579),
.A2(n_583),
.B1(n_585),
.B2(n_588),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_SL g582 ( 
.A(n_555),
.B(n_525),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_582),
.B(n_526),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_543),
.A2(n_510),
.B1(n_507),
.B2(n_502),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_549),
.B(n_522),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_554),
.A2(n_507),
.B1(n_502),
.B2(n_520),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_542),
.A2(n_515),
.B1(n_537),
.B2(n_538),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_541),
.A2(n_505),
.B1(n_529),
.B2(n_538),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_540),
.A2(n_505),
.B1(n_537),
.B2(n_517),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_555),
.B(n_524),
.C(n_509),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_595),
.B(n_562),
.C(n_553),
.Y(n_614)
);

INVx6_ASAP7_75t_L g600 ( 
.A(n_568),
.Y(n_600)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_600),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_551),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_SL g604 ( 
.A(n_601),
.B(n_546),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_540),
.A2(n_533),
.B1(n_516),
.B2(n_536),
.Y(n_603)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_604),
.Y(n_633)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_597),
.Y(n_605)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_605),
.Y(n_639)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_589),
.B(n_561),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g637 ( 
.A(n_609),
.B(n_611),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_SL g610 ( 
.A(n_595),
.B(n_531),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_610),
.B(n_614),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_598),
.B(n_557),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_613),
.B(n_616),
.Y(n_640)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_597),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_578),
.B(n_548),
.C(n_574),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_617),
.B(n_618),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_580),
.B(n_532),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_580),
.B(n_603),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g638 ( 
.A(n_619),
.B(n_620),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_588),
.B(n_591),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_602),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_621),
.B(n_622),
.Y(n_632)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_602),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_591),
.B(n_548),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g643 ( 
.A(n_623),
.B(n_624),
.Y(n_643)
);

XOR2xp5_ASAP7_75t_L g624 ( 
.A(n_582),
.B(n_545),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_581),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_625),
.B(n_626),
.Y(n_641)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_581),
.Y(n_626)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_585),
.B(n_544),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_627),
.B(n_628),
.Y(n_644)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_583),
.B(n_545),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_614),
.B(n_575),
.C(n_579),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g650 ( 
.A(n_629),
.B(n_630),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_606),
.B(n_587),
.C(n_594),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_606),
.B(n_550),
.C(n_566),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g651 ( 
.A(n_631),
.B(n_635),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_623),
.A2(n_593),
.B(n_550),
.Y(n_634)
);

NOR3xp33_ASAP7_75t_L g660 ( 
.A(n_634),
.B(n_649),
.C(n_563),
.Y(n_660)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_609),
.B(n_590),
.C(n_576),
.Y(n_635)
);

FAx1_ASAP7_75t_SL g636 ( 
.A(n_617),
.B(n_546),
.CI(n_547),
.CON(n_636),
.SN(n_636)
);

AOI22xp5_ASAP7_75t_SL g665 ( 
.A1(n_636),
.A2(n_599),
.B1(n_570),
.B2(n_568),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_620),
.A2(n_586),
.B(n_590),
.Y(n_642)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_642),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_615),
.A2(n_596),
.B1(n_592),
.B2(n_569),
.Y(n_646)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_646),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_613),
.B(n_576),
.C(n_556),
.Y(n_648)
);

XNOR2xp5_ASAP7_75t_L g658 ( 
.A(n_648),
.B(n_619),
.Y(n_658)
);

OAI21xp5_ASAP7_75t_SL g649 ( 
.A1(n_607),
.A2(n_586),
.B(n_559),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_SL g652 ( 
.A(n_645),
.B(n_627),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_652),
.B(n_659),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_633),
.B(n_608),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_653),
.B(n_654),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_SL g654 ( 
.A1(n_639),
.A2(n_612),
.B1(n_567),
.B2(n_572),
.Y(n_654)
);

XNOR2xp5_ASAP7_75t_L g655 ( 
.A(n_647),
.B(n_612),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_655),
.B(n_656),
.Y(n_675)
);

XNOR2xp5_ASAP7_75t_L g656 ( 
.A(n_635),
.B(n_628),
.Y(n_656)
);

XOR2xp5_ASAP7_75t_SL g657 ( 
.A(n_643),
.B(n_624),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_657),
.B(n_637),
.Y(n_671)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_658),
.Y(n_669)
);

XOR2xp5_ASAP7_75t_L g659 ( 
.A(n_643),
.B(n_611),
.Y(n_659)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_660),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g661 ( 
.A(n_629),
.B(n_599),
.C(n_558),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g668 ( 
.A(n_661),
.B(n_666),
.C(n_631),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_SL g664 ( 
.A1(n_640),
.A2(n_573),
.B1(n_565),
.B2(n_571),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_664),
.A2(n_644),
.B1(n_420),
.B2(n_406),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_665),
.A2(n_644),
.B(n_638),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_630),
.B(n_570),
.C(n_600),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_SL g667 ( 
.A1(n_665),
.A2(n_634),
.B(n_641),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_667),
.B(n_676),
.Y(n_680)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_668),
.Y(n_685)
);

XNOR2xp5_ASAP7_75t_L g683 ( 
.A(n_671),
.B(n_678),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_672),
.A2(n_679),
.B1(n_659),
.B2(n_656),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_651),
.A2(n_632),
.B(n_637),
.Y(n_674)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_674),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_SL g676 ( 
.A1(n_663),
.A2(n_642),
.B1(n_636),
.B2(n_649),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_SL g678 ( 
.A1(n_662),
.A2(n_648),
.B1(n_636),
.B2(n_638),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_668),
.B(n_666),
.Y(n_681)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_681),
.Y(n_694)
);

INVx11_ASAP7_75t_L g682 ( 
.A(n_675),
.Y(n_682)
);

AOI21xp33_ASAP7_75t_L g691 ( 
.A1(n_682),
.A2(n_687),
.B(n_670),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_675),
.B(n_655),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_684),
.A2(n_686),
.B(n_672),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_669),
.B(n_661),
.Y(n_686)
);

AOI21x1_ASAP7_75t_L g696 ( 
.A1(n_689),
.A2(n_693),
.B(n_682),
.Y(n_696)
);

MAJIxp5_ASAP7_75t_L g690 ( 
.A(n_685),
.B(n_650),
.C(n_673),
.Y(n_690)
);

XOR2xp5_ASAP7_75t_L g695 ( 
.A(n_690),
.B(n_691),
.Y(n_695)
);

MAJIxp5_ASAP7_75t_L g692 ( 
.A(n_688),
.B(n_677),
.C(n_678),
.Y(n_692)
);

MAJIxp5_ASAP7_75t_L g697 ( 
.A(n_692),
.B(n_683),
.C(n_687),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_SL g693 ( 
.A1(n_680),
.A2(n_679),
.B(n_657),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_696),
.A2(n_695),
.B(n_683),
.Y(n_698)
);

MAJIxp5_ASAP7_75t_L g699 ( 
.A(n_697),
.B(n_694),
.C(n_690),
.Y(n_699)
);

MAJIxp5_ASAP7_75t_L g700 ( 
.A(n_698),
.B(n_699),
.C(n_381),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_700),
.B(n_329),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_701),
.A2(n_329),
.B(n_316),
.Y(n_702)
);

XOR2xp5_ASAP7_75t_L g703 ( 
.A(n_702),
.B(n_352),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_703),
.A2(n_352),
.B(n_653),
.Y(n_704)
);


endmodule