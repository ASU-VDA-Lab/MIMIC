module real_jpeg_10616_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_191;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx24_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_SL g71 ( 
.A(n_5),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_7),
.A2(n_27),
.B1(n_30),
.B2(n_48),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_8),
.A2(n_53),
.B1(n_62),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_8),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_103),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_8),
.A2(n_27),
.B1(n_30),
.B2(n_103),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_8),
.A2(n_38),
.B1(n_39),
.B2(n_103),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_9),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_9),
.A2(n_55),
.B(n_59),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_9),
.A2(n_53),
.B1(n_62),
.B2(n_126),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_9),
.B(n_66),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_9),
.A2(n_38),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_9),
.B(n_38),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_9),
.A2(n_83),
.B1(n_84),
.B2(n_202),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_10),
.A2(n_53),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_10),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_63),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_10),
.A2(n_27),
.B1(n_30),
.B2(n_63),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_63),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_12),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_12),
.A2(n_35),
.B1(n_53),
.B2(n_62),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_12),
.A2(n_35),
.B1(n_58),
.B2(n_59),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_12),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_13),
.A2(n_53),
.B1(n_62),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_13),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_122),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_122),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_13),
.A2(n_27),
.B1(n_30),
.B2(n_122),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_14),
.A2(n_41),
.B1(n_58),
.B2(n_59),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_14),
.A2(n_27),
.B1(n_30),
.B2(n_41),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_15),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_15),
.A2(n_29),
.B1(n_58),
.B2(n_59),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_15),
.A2(n_29),
.B1(n_38),
.B2(n_39),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_132),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_107),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_19),
.B(n_107),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_91),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_79),
.B2(n_80),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_49),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_24),
.B(n_36),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_25),
.A2(n_84),
.B(n_129),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_26),
.B(n_32),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_27),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_27),
.A2(n_30),
.B1(n_43),
.B2(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_27),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_193)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_30),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_30),
.B(n_46),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_30),
.B(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_31),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_31),
.A2(n_32),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_32),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_33),
.A2(n_83),
.B(n_186),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_34),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_37),
.A2(n_45),
.B(n_97),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_43),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_39),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_38),
.B(n_70),
.Y(n_230)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_39),
.A2(n_75),
.B1(n_225),
.B2(n_230),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_42),
.A2(n_47),
.B(n_87),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_42),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_42),
.A2(n_45),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_42),
.A2(n_45),
.B1(n_192),
.B2(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_42),
.A2(n_45),
.B1(n_215),
.B2(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_42),
.A2(n_223),
.B(n_246),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_44),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_45),
.B(n_126),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_45),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_67),
.B2(n_78),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_61),
.B(n_64),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_52),
.A2(n_57),
.B1(n_61),
.B2(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_52),
.A2(n_57),
.B1(n_102),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_52),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B(n_56),
.C(n_57),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_54),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_53),
.A2(n_54),
.B(n_126),
.C(n_127),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_69),
.B(n_70),
.C(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_70),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g225 ( 
.A(n_59),
.B(n_126),
.CON(n_225),
.SN(n_225)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_66),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_67),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B(n_73),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_77),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_68),
.A2(n_116),
.B1(n_117),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_68),
.A2(n_116),
.B1(n_146),
.B2(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_68),
.B(n_126),
.Y(n_213)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_105),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_69),
.A2(n_74),
.B1(n_170),
.B2(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_74),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_90),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B(n_85),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_83),
.A2(n_84),
.B1(n_94),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_83),
.A2(n_84),
.B1(n_184),
.B2(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_83),
.A2(n_85),
.B(n_95),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_84),
.B(n_126),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_88),
.A2(n_99),
.B(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_100),
.C(n_104),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_96),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_101),
.B1(n_104),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.C(n_112),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_108),
.B(n_111),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_112),
.A2(n_113),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.C(n_123),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_115),
.B1(n_119),
.B2(n_120),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_125),
.B1(n_128),
.B2(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_128),
.Y(n_164)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_175),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_156),
.B(n_174),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_176),
.C(n_257),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_153),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_153),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_142),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.C(n_151),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_145),
.B1(n_151),
.B2(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_151),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_152),
.B(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_157),
.B(n_159),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_165),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_160),
.B(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_163),
.A2(n_165),
.B1(n_166),
.B2(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_163),
.Y(n_255)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_171),
.C(n_172),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_167),
.A2(n_168),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_171),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_251),
.B(n_256),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_234),
.B(n_250),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_218),
.B(n_233),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_209),
.B(n_217),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_198),
.B(n_208),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_187),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_182),
.B(n_187),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_193),
.B2(n_197),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_188),
.B(n_197),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_191),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_193),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_203),
.B(n_207),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_200),
.B(n_201),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_210),
.B(n_211),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_219),
.Y(n_233)
);

FAx1_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.CI(n_216),
.CON(n_212),
.SN(n_212)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_228),
.B2(n_232),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_222),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_224),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_227),
.C(n_232),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_228),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_231),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_235),
.B(n_236),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_242),
.B2(n_243),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_245),
.C(n_248),
.Y(n_252)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_248),
.B2(n_249),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_244),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_245),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_252),
.B(n_253),
.Y(n_256)
);


endmodule