module fake_jpeg_3031_n_184 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_184);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_21),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_16),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_66),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_65),
.Y(n_70)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_51),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_68),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_38),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_68),
.B1(n_65),
.B2(n_64),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_66),
.B1(n_44),
.B2(n_45),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_54),
.B1(n_50),
.B2(n_56),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_44),
.B1(n_50),
.B2(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_92),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_45),
.B1(n_56),
.B2(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_89),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_79),
.B(n_73),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_91),
.B(n_44),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_61),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_1),
.Y(n_113)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_36),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_102),
.B1(n_94),
.B2(n_2),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_60),
.B1(n_61),
.B2(n_59),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_111),
.Y(n_117)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_59),
.B1(n_55),
.B2(n_53),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_112),
.B1(n_4),
.B2(n_5),
.Y(n_127)
);

OAI22x1_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_49),
.B1(n_55),
.B2(n_53),
.Y(n_108)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_47),
.C(n_57),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_81),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_47),
.B1(n_58),
.B2(n_49),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_4),
.C(n_5),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_111),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_127),
.Y(n_134)
);

AOI32xp33_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_96),
.A3(n_83),
.B1(n_91),
.B2(n_49),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_118),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_81),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_119),
.B(n_123),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_126),
.B1(n_98),
.B2(n_109),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_107),
.B(n_106),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_132),
.B(n_120),
.Y(n_149)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_129),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_98),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_24),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_37),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_131),
.B(n_32),
.Y(n_143)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_148),
.B1(n_10),
.B2(n_11),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_142),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_34),
.C(n_33),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_144),
.C(n_145),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_147),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_30),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_29),
.C(n_28),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_121),
.B(n_6),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_146),
.B(n_149),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_26),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_148)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_140),
.A2(n_133),
.B1(n_131),
.B2(n_125),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_155),
.B1(n_160),
.B2(n_163),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_23),
.Y(n_159)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_170),
.C(n_159),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_141),
.C(n_139),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_169),
.C(n_156),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_163),
.A2(n_144),
.B1(n_139),
.B2(n_147),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_173),
.A2(n_174),
.B(n_175),
.Y(n_178)
);

OAI322xp33_ASAP7_75t_L g174 ( 
.A1(n_164),
.A2(n_161),
.A3(n_152),
.B1(n_156),
.B2(n_155),
.C1(n_145),
.C2(n_22),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_12),
.C(n_13),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_164),
.B(n_169),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_166),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_177),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_178),
.C(n_165),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_167),
.A3(n_15),
.B1(n_17),
.B2(n_18),
.C1(n_19),
.C2(n_20),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_19),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_14),
.Y(n_184)
);


endmodule