module real_jpeg_27419_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_300;
wire n_221;
wire n_286;
wire n_288;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_299;
wire n_255;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_295;
wire n_167;
wire n_179;
wire n_216;
wire n_202;
wire n_133;
wire n_213;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_L g88 ( 
.A(n_0),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_0),
.B(n_232),
.Y(n_237)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_0),
.Y(n_248)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_2),
.A2(n_32),
.B1(n_46),
.B2(n_50),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_2),
.A2(n_32),
.B1(n_52),
.B2(n_54),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_4),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_137),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_4),
.A2(n_46),
.B1(n_50),
.B2(n_137),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_4),
.A2(n_52),
.B1(n_54),
.B2(n_137),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_6),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_6),
.A2(n_46),
.B1(n_50),
.B2(n_69),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_69),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_6),
.A2(n_52),
.B1(n_54),
.B2(n_69),
.Y(n_152)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_8),
.A2(n_30),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_8),
.B(n_30),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_8),
.A2(n_46),
.B1(n_50),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_8),
.A2(n_52),
.B1(n_54),
.B2(n_58),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_8),
.B(n_21),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_SL g198 ( 
.A1(n_8),
.A2(n_10),
.B(n_46),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_8),
.A2(n_49),
.B(n_52),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_8),
.B(n_65),
.Y(n_227)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_11),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_112),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_111),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_94),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_16),
.B(n_94),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_73),
.C(n_81),
.Y(n_16)
);

FAx1_ASAP7_75t_SL g143 ( 
.A(n_17),
.B(n_73),
.CI(n_81),
.CON(n_143),
.SN(n_143)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_39),
.B2(n_40),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_18),
.A2(n_19),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_19),
.B(n_41),
.C(n_60),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_33),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_20),
.B(n_133),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_28),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_21),
.B(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_22),
.A2(n_23),
.B(n_30),
.C(n_36),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_22),
.A2(n_35),
.B(n_37),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_22),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_22),
.B(n_136),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_22)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_24),
.B(n_27),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_25),
.A2(n_62),
.B(n_63),
.C(n_65),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_25),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_25),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_25),
.A2(n_58),
.B(n_197),
.C(n_198),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_29),
.B(n_35),
.Y(n_101)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_34),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_35),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_36),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_37),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_38),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_59),
.B2(n_60),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_41),
.B(n_157),
.C(n_159),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_41),
.A2(n_42),
.B1(n_159),
.B2(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_42),
.B(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_55),
.B(n_56),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_43),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_44),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_44),
.B(n_57),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_44),
.B(n_205),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_51),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_50),
.B1(n_64),
.B2(n_66),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_46),
.A2(n_48),
.B(n_58),
.C(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_49),
.B1(n_52),
.B2(n_54),
.Y(n_51)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_51),
.B(n_57),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_51),
.B(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_51),
.B(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_52),
.Y(n_54)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_54),
.B(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_55),
.A2(n_79),
.B(n_91),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_55),
.B(n_58),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_58),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_67),
.B(n_70),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_61),
.B(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_61),
.B(n_162),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_61),
.Y(n_279)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_65),
.B(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_66),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_75),
.B(n_76),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_71),
.B(n_170),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_73),
.A2(n_74),
.B(n_77),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_75),
.A2(n_106),
.B(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_76),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_76),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_78),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_79),
.B(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B(n_93),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_82),
.A2(n_83),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_90),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_84),
.A2(n_85),
.B1(n_93),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_84),
.A2(n_85),
.B1(n_196),
.B2(n_199),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_84),
.A2(n_85),
.B1(n_90),
.B2(n_293),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_85),
.B(n_196),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_89),
.Y(n_85)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_86),
.B(n_89),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_86),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_87),
.B(n_89),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_87),
.B(n_123),
.Y(n_153)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_87),
.Y(n_177)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_90),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_92),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_92),
.B(n_214),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_93),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_110),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_102),
.B1(n_103),
.B2(n_109),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_101),
.B(n_158),
.Y(n_276)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_105),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_144),
.B(n_302),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_143),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_114),
.B(n_143),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_138),
.C(n_139),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_115),
.A2(n_116),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_126),
.C(n_129),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_117),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_125),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_118),
.B(n_125),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_119),
.B(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_120),
.A2(n_152),
.B(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_121),
.B(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_126),
.A2(n_129),
.B1(n_130),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_126),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_128),
.B(n_161),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_138),
.B(n_139),
.Y(n_300)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_143),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_296),
.B(n_301),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_283),
.B(n_295),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_190),
.B(n_266),
.C(n_282),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_178),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_148),
.B(n_178),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_163),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_156),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_150),
.B(n_156),
.C(n_163),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_151),
.B(n_154),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_153),
.B(n_231),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_155),
.B(n_204),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_171),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_165),
.B(n_168),
.C(n_171),
.Y(n_280)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_176),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.C(n_184),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_179),
.A2(n_180),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_184),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.C(n_188),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_188),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_189),
.B(n_237),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_265),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_258),
.B(n_264),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_216),
.B(n_257),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_206),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_194),
.B(n_206),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_200),
.C(n_202),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_195),
.B(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_196),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_255)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_211),
.B2(n_212),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_207),
.B(n_213),
.C(n_215),
.Y(n_259)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_252),
.B(n_256),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_233),
.B(n_251),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_224),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_219),
.B(n_224),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_222),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_230),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_229),
.C(n_230),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_240),
.B(n_250),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_235),
.B(n_238),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_244),
.B(n_249),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_242),
.B(n_243),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_253),
.B(n_254),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_259),
.B(n_260),
.Y(n_264)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_267),
.B(n_268),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_280),
.B2(n_281),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_272),
.C(n_281),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_276),
.C(n_277),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_284),
.B(n_285),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_294),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_291),
.B2(n_292),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_292),
.C(n_294),
.Y(n_297)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_298),
.Y(n_301)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);


endmodule