module fake_netlist_1_8157_n_682 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_682);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_682;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_47), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_68), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_73), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_26), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_70), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_35), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_62), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_50), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_23), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_18), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_66), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_21), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_37), .Y(n_89) );
INVxp67_ASAP7_75t_L g90 ( .A(n_46), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_61), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_21), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_36), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_40), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_42), .Y(n_95) );
CKINVDCx16_ASAP7_75t_R g96 ( .A(n_6), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_56), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_20), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_22), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_6), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_10), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_65), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_18), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_30), .Y(n_104) );
BUFx2_ASAP7_75t_SL g105 ( .A(n_52), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_7), .Y(n_106) );
INVxp33_ASAP7_75t_SL g107 ( .A(n_67), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_14), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_23), .Y(n_109) );
INVxp33_ASAP7_75t_SL g110 ( .A(n_20), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_71), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_17), .Y(n_112) );
INVxp33_ASAP7_75t_L g113 ( .A(n_64), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_16), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_60), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_31), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_10), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_48), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_7), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_75), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_74), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_17), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_59), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_5), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_33), .Y(n_125) );
INVxp67_ASAP7_75t_L g126 ( .A(n_109), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_124), .Y(n_127) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_124), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_120), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_82), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_77), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_82), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_77), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_100), .B(n_0), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_120), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_89), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_96), .B(n_0), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_78), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_78), .Y(n_139) );
NOR2xp33_ASAP7_75t_R g140 ( .A(n_89), .B(n_32), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_79), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_96), .B(n_1), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_107), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_110), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_120), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_85), .B(n_1), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_80), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_100), .B(n_2), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_80), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_83), .Y(n_150) );
INVx1_ASAP7_75t_SL g151 ( .A(n_84), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_87), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_87), .Y(n_153) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_85), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_93), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_115), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_105), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_86), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_93), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_105), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_94), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_91), .B(n_2), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_103), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_90), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_94), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_95), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_95), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_103), .B(n_3), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_81), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_127), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_151), .B(n_113), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_147), .Y(n_172) );
BUFx2_ASAP7_75t_L g173 ( .A(n_151), .Y(n_173) );
INVxp67_ASAP7_75t_L g174 ( .A(n_128), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_137), .A2(n_108), .B1(n_88), .B2(n_122), .Y(n_176) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_126), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_147), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_149), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_135), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_128), .B(n_126), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_135), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_149), .Y(n_183) );
INVx5_ASAP7_75t_L g184 ( .A(n_135), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_135), .Y(n_185) );
INVx1_ASAP7_75t_SL g186 ( .A(n_130), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_149), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_153), .Y(n_188) );
BUFx2_ASAP7_75t_L g189 ( .A(n_132), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_135), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_135), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_153), .Y(n_192) );
NAND2x1p5_ASAP7_75t_L g193 ( .A(n_134), .B(n_125), .Y(n_193) );
NAND2x1p5_ASAP7_75t_L g194 ( .A(n_134), .B(n_125), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_154), .B(n_117), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_153), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_129), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_164), .B(n_123), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_155), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_155), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_129), .Y(n_202) );
NAND2x1p5_ASAP7_75t_L g203 ( .A(n_134), .B(n_123), .Y(n_203) );
OAI21xp33_ASAP7_75t_L g204 ( .A1(n_131), .A2(n_122), .B(n_86), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_159), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_157), .B(n_121), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_129), .Y(n_207) );
INVxp33_ASAP7_75t_L g208 ( .A(n_137), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_159), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_134), .B(n_117), .Y(n_210) );
NAND3xp33_ASAP7_75t_L g211 ( .A(n_154), .B(n_106), .C(n_119), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_145), .Y(n_212) );
AND2x2_ASAP7_75t_SL g213 ( .A(n_148), .B(n_121), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_145), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_148), .B(n_119), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_159), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_148), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_145), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_131), .B(n_118), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_127), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_127), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_133), .B(n_118), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_165), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_137), .B(n_88), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_163), .B(n_133), .Y(n_225) );
INVx4_ASAP7_75t_L g226 ( .A(n_148), .Y(n_226) );
NAND3x1_ASAP7_75t_L g227 ( .A(n_146), .B(n_92), .C(n_112), .Y(n_227) );
NAND2x1p5_ASAP7_75t_L g228 ( .A(n_168), .B(n_104), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_127), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_165), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_165), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_213), .A2(n_138), .B(n_161), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_226), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g234 ( .A1(n_181), .A2(n_142), .B(n_146), .C(n_167), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_224), .B(n_168), .Y(n_235) );
INVxp67_ASAP7_75t_L g236 ( .A(n_173), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_210), .Y(n_237) );
NOR2xp33_ASAP7_75t_R g238 ( .A(n_173), .B(n_141), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_217), .A2(n_139), .B(n_138), .C(n_167), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_177), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_171), .B(n_169), .Y(n_241) );
OR2x6_ASAP7_75t_SL g242 ( .A(n_208), .B(n_136), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_223), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_210), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_174), .B(n_144), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_223), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_189), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_223), .Y(n_248) );
INVx3_ASAP7_75t_L g249 ( .A(n_226), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_223), .Y(n_250) );
NOR3xp33_ASAP7_75t_SL g251 ( .A(n_211), .B(n_143), .C(n_160), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_210), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_189), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_186), .B(n_163), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_210), .Y(n_255) );
INVx1_ASAP7_75t_SL g256 ( .A(n_224), .Y(n_256) );
INVxp67_ASAP7_75t_SL g257 ( .A(n_193), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_215), .B(n_168), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_215), .B(n_168), .Y(n_259) );
INVx6_ASAP7_75t_L g260 ( .A(n_226), .Y(n_260) );
INVx3_ASAP7_75t_SL g261 ( .A(n_213), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_225), .B(n_150), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_193), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_170), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_223), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_193), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_194), .Y(n_267) );
AND3x2_ASAP7_75t_SL g268 ( .A(n_213), .B(n_158), .C(n_140), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_176), .B(n_161), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_225), .B(n_156), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_194), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_195), .B(n_152), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_170), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_176), .Y(n_274) );
OR2x2_ASAP7_75t_L g275 ( .A(n_195), .B(n_152), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_202), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_194), .B(n_139), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_203), .B(n_162), .Y(n_278) );
BUFx8_ASAP7_75t_SL g279 ( .A(n_215), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_203), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_203), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_215), .B(n_162), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_228), .B(n_166), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_228), .B(n_166), .Y(n_284) );
INVx2_ASAP7_75t_SL g285 ( .A(n_228), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_206), .B(n_166), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_172), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_199), .B(n_217), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_202), .Y(n_289) );
BUFx8_ASAP7_75t_L g290 ( .A(n_172), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_217), .B(n_116), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_227), .Y(n_292) );
AND2x2_ASAP7_75t_SL g293 ( .A(n_219), .B(n_102), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_222), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_220), .B(n_102), .Y(n_295) );
NOR2xp67_ASAP7_75t_L g296 ( .A(n_204), .B(n_3), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_202), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_175), .Y(n_298) );
AND2x6_ASAP7_75t_L g299 ( .A(n_263), .B(n_175), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_236), .B(n_178), .Y(n_300) );
INVx5_ASAP7_75t_L g301 ( .A(n_285), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_277), .A2(n_229), .B(n_221), .Y(n_302) );
INVx2_ASAP7_75t_SL g303 ( .A(n_285), .Y(n_303) );
INVx5_ASAP7_75t_L g304 ( .A(n_260), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_277), .A2(n_229), .B(n_221), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_261), .A2(n_220), .B1(n_196), .B2(n_231), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_273), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_261), .B(n_178), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_290), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_283), .A2(n_198), .B(n_212), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_239), .A2(n_231), .B(n_179), .C(n_183), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_257), .B(n_266), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_294), .B(n_179), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_237), .Y(n_314) );
OAI21x1_ASAP7_75t_SL g315 ( .A1(n_232), .A2(n_187), .B(n_183), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_244), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_267), .B(n_187), .Y(n_317) );
INVx2_ASAP7_75t_SL g318 ( .A(n_290), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_252), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_294), .B(n_92), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_290), .Y(n_321) );
INVx3_ASAP7_75t_SL g322 ( .A(n_247), .Y(n_322) );
INVx3_ASAP7_75t_SL g323 ( .A(n_247), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_255), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_254), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_264), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_258), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_273), .Y(n_328) );
INVx2_ASAP7_75t_SL g329 ( .A(n_271), .Y(n_329) );
OR2x6_ASAP7_75t_L g330 ( .A(n_280), .B(n_227), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_292), .A2(n_209), .B1(n_188), .B2(n_216), .Y(n_331) );
A2O1A1Ixp33_ASAP7_75t_L g332 ( .A1(n_239), .A2(n_200), .B(n_188), .C(n_216), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_281), .Y(n_333) );
INVx1_ASAP7_75t_SL g334 ( .A(n_254), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_283), .A2(n_198), .B(n_218), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_258), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_289), .Y(n_337) );
A2O1A1Ixp33_ASAP7_75t_L g338 ( .A1(n_288), .A2(n_201), .B(n_192), .C(n_196), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_258), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_235), .A2(n_200), .B1(n_192), .B2(n_197), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_240), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_284), .A2(n_218), .B(n_212), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_240), .B(n_197), .Y(n_343) );
OAI21x1_ASAP7_75t_SL g344 ( .A1(n_282), .A2(n_209), .B(n_205), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_259), .Y(n_345) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_289), .Y(n_346) );
INVx2_ASAP7_75t_SL g347 ( .A(n_260), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_273), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_264), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_238), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_235), .B(n_201), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_299), .Y(n_352) );
INVx3_ASAP7_75t_SL g353 ( .A(n_318), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_313), .B(n_256), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_325), .A2(n_274), .B1(n_279), .B2(n_278), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_313), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_322), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_334), .B(n_272), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_312), .B(n_235), .Y(n_359) );
A2O1A1Ixp33_ASAP7_75t_L g360 ( .A1(n_338), .A2(n_286), .B(n_234), .C(n_259), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_341), .A2(n_274), .B1(n_279), .B2(n_278), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_322), .Y(n_362) );
NAND2x1p5_ASAP7_75t_L g363 ( .A(n_312), .B(n_233), .Y(n_363) );
INVx2_ASAP7_75t_SL g364 ( .A(n_301), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_337), .Y(n_365) );
OA21x2_ASAP7_75t_L g366 ( .A1(n_338), .A2(n_185), .B(n_182), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_300), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_343), .Y(n_368) );
AOI22xp33_ASAP7_75t_SL g369 ( .A1(n_318), .A2(n_253), .B1(n_268), .B2(n_293), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_301), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_323), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_312), .B(n_259), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_299), .A2(n_245), .B1(n_270), .B2(n_262), .Y(n_373) );
AOI222xp33_ASAP7_75t_L g374 ( .A1(n_320), .A2(n_241), .B1(n_293), .B2(n_98), .C1(n_101), .C2(n_106), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_302), .A2(n_284), .B(n_291), .Y(n_375) );
AO221x2_ASAP7_75t_L g376 ( .A1(n_330), .A2(n_268), .B1(n_98), .B2(n_99), .C(n_114), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_321), .B(n_233), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_320), .A2(n_245), .B1(n_269), .B2(n_249), .Y(n_378) );
AOI222xp33_ASAP7_75t_L g379 ( .A1(n_323), .A2(n_108), .B1(n_99), .B2(n_114), .C1(n_112), .C2(n_101), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_317), .Y(n_380) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_299), .Y(n_381) );
CKINVDCx12_ASAP7_75t_R g382 ( .A(n_330), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_350), .Y(n_383) );
AOI21xp33_ASAP7_75t_L g384 ( .A1(n_330), .A2(n_275), .B(n_249), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_321), .B(n_233), .Y(n_385) );
NAND4xp25_ASAP7_75t_L g386 ( .A(n_379), .B(n_296), .C(n_340), .D(n_332), .Y(n_386) );
OAI22xp33_ASAP7_75t_L g387 ( .A1(n_373), .A2(n_309), .B1(n_330), .B2(n_242), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_376), .A2(n_351), .B1(n_344), .B2(n_308), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_365), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_354), .A2(n_331), .B1(n_332), .B2(n_311), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_378), .A2(n_356), .B1(n_354), .B2(n_367), .C(n_368), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_381), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_380), .Y(n_393) );
OAI33xp33_ASAP7_75t_L g394 ( .A1(n_358), .A2(n_295), .A3(n_97), .B1(n_111), .B2(n_104), .B3(n_205), .Y(n_394) );
OAI211xp5_ASAP7_75t_SL g395 ( .A1(n_374), .A2(n_251), .B(n_311), .C(n_316), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_363), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_365), .Y(n_397) );
INVx4_ASAP7_75t_L g398 ( .A(n_381), .Y(n_398) );
OAI22xp33_ASAP7_75t_SL g399 ( .A1(n_352), .A2(n_242), .B1(n_329), .B2(n_301), .Y(n_399) );
OAI21x1_ASAP7_75t_L g400 ( .A1(n_366), .A2(n_315), .B(n_335), .Y(n_400) );
AOI21x1_ASAP7_75t_L g401 ( .A1(n_366), .A2(n_310), .B(n_342), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_359), .B(n_308), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_363), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_376), .A2(n_299), .B1(n_351), .B2(n_317), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_381), .Y(n_405) );
A2O1A1Ixp33_ASAP7_75t_L g406 ( .A1(n_360), .A2(n_329), .B(n_317), .C(n_303), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_376), .A2(n_351), .B1(n_299), .B2(n_327), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_357), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_359), .B(n_333), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_369), .A2(n_299), .B1(n_336), .B2(n_339), .Y(n_410) );
INVx2_ASAP7_75t_SL g411 ( .A(n_381), .Y(n_411) );
OAI22xp33_ASAP7_75t_L g412 ( .A1(n_362), .A2(n_301), .B1(n_303), .B2(n_333), .Y(n_412) );
AND2x4_ASAP7_75t_L g413 ( .A(n_352), .B(n_301), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_366), .Y(n_414) );
NAND4xp25_ASAP7_75t_L g415 ( .A(n_391), .B(n_355), .C(n_361), .D(n_410), .Y(n_415) );
OA21x2_ASAP7_75t_L g416 ( .A1(n_400), .A2(n_375), .B(n_384), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_404), .A2(n_359), .B1(n_382), .B2(n_352), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_391), .A2(n_382), .B1(n_372), .B2(n_362), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_396), .B(n_364), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_399), .B(n_364), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_414), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_396), .Y(n_422) );
NOR2xp33_ASAP7_75t_R g423 ( .A(n_403), .B(n_357), .Y(n_423) );
OA21x2_ASAP7_75t_L g424 ( .A1(n_400), .A2(n_305), .B(n_111), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_414), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_393), .Y(n_426) );
AOI33xp33_ASAP7_75t_L g427 ( .A1(n_387), .A2(n_97), .A3(n_385), .B1(n_377), .B2(n_345), .B3(n_314), .Y(n_427) );
OAI321xp33_ASAP7_75t_L g428 ( .A1(n_395), .A2(n_370), .A3(n_324), .B1(n_319), .B2(n_306), .C(n_333), .Y(n_428) );
BUFx2_ASAP7_75t_L g429 ( .A(n_405), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_390), .B(n_372), .Y(n_430) );
BUFx2_ASAP7_75t_SL g431 ( .A(n_403), .Y(n_431) );
AOI222xp33_ASAP7_75t_L g432 ( .A1(n_395), .A2(n_353), .B1(n_372), .B2(n_383), .C1(n_371), .C2(n_385), .Y(n_432) );
NOR2xp33_ASAP7_75t_R g433 ( .A(n_408), .B(n_371), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_390), .B(n_333), .Y(n_434) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_404), .Y(n_435) );
OAI31xp33_ASAP7_75t_L g436 ( .A1(n_399), .A2(n_385), .A3(n_377), .B(n_370), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_414), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_402), .Y(n_438) );
OAI211xp5_ASAP7_75t_L g439 ( .A1(n_407), .A2(n_383), .B(n_298), .C(n_287), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_393), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_406), .A2(n_337), .B(n_346), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_402), .B(n_230), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_388), .B(n_377), .Y(n_443) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_401), .A2(n_182), .B(n_185), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_409), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_389), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_409), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_389), .Y(n_448) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_392), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_423), .B(n_436), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_441), .A2(n_394), .B(n_412), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_426), .Y(n_452) );
AOI211xp5_ASAP7_75t_L g453 ( .A1(n_415), .A2(n_353), .B(n_386), .C(n_394), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g454 ( .A(n_432), .B(n_386), .C(n_397), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_421), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_421), .Y(n_456) );
INVx2_ASAP7_75t_SL g457 ( .A(n_422), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_430), .B(n_389), .Y(n_458) );
CKINVDCx16_ASAP7_75t_R g459 ( .A(n_431), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_449), .Y(n_460) );
OAI33xp33_ASAP7_75t_L g461 ( .A1(n_426), .A2(n_4), .A3(n_5), .B1(n_8), .B2(n_9), .B3(n_11), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_440), .Y(n_462) );
OAI31xp33_ASAP7_75t_L g463 ( .A1(n_439), .A2(n_413), .A3(n_405), .B(n_411), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_421), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_440), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_425), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_425), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_446), .B(n_397), .Y(n_468) );
NOR2xp67_ASAP7_75t_L g469 ( .A(n_418), .B(n_398), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_438), .B(n_397), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_418), .A2(n_413), .B1(n_392), .B2(n_398), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_446), .B(n_400), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_430), .A2(n_413), .B1(n_348), .B2(n_307), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_433), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_448), .B(n_398), .Y(n_475) );
AOI31xp33_ASAP7_75t_L g476 ( .A1(n_417), .A2(n_4), .A3(n_8), .B(n_9), .Y(n_476) );
NAND4xp25_ASAP7_75t_L g477 ( .A(n_427), .B(n_11), .C(n_12), .D(n_13), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_445), .B(n_12), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_447), .B(n_13), .Y(n_479) );
OAI221xp5_ASAP7_75t_L g480 ( .A1(n_436), .A2(n_443), .B1(n_417), .B2(n_435), .C(n_419), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_447), .B(n_14), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_428), .A2(n_214), .B1(n_207), .B2(n_202), .C(n_347), .Y(n_482) );
NOR4xp25_ASAP7_75t_L g483 ( .A(n_428), .B(n_15), .C(n_16), .D(n_19), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_442), .B(n_15), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_425), .Y(n_485) );
NAND3xp33_ASAP7_75t_L g486 ( .A(n_420), .B(n_207), .C(n_214), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_437), .B(n_214), .Y(n_487) );
OAI21xp33_ASAP7_75t_L g488 ( .A1(n_434), .A2(n_207), .B(n_214), .Y(n_488) );
INVx1_ASAP7_75t_SL g489 ( .A(n_431), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_437), .B(n_19), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_422), .B(n_76), .Y(n_491) );
INVx2_ASAP7_75t_SL g492 ( .A(n_419), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_442), .B(n_22), .Y(n_493) );
AOI33xp33_ASAP7_75t_L g494 ( .A1(n_437), .A2(n_347), .A3(n_248), .B1(n_250), .B2(n_265), .B3(n_246), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_443), .B(n_207), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_492), .B(n_429), .Y(n_496) );
NAND2x1p5_ASAP7_75t_L g497 ( .A(n_491), .B(n_429), .Y(n_497) );
NOR2xp33_ASAP7_75t_R g498 ( .A(n_459), .B(n_449), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_455), .Y(n_499) );
NAND4xp75_ASAP7_75t_L g500 ( .A(n_450), .B(n_434), .C(n_416), .D(n_424), .Y(n_500) );
INVx4_ASAP7_75t_L g501 ( .A(n_459), .Y(n_501) );
AOI32xp33_ASAP7_75t_L g502 ( .A1(n_474), .A2(n_307), .A3(n_348), .B1(n_328), .B2(n_349), .Y(n_502) );
NAND2xp33_ASAP7_75t_R g503 ( .A(n_491), .B(n_424), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_477), .A2(n_416), .B1(n_424), .B2(n_449), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_455), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_452), .Y(n_506) );
NOR2xp33_ASAP7_75t_R g507 ( .A(n_489), .B(n_457), .Y(n_507) );
INVx3_ASAP7_75t_L g508 ( .A(n_456), .Y(n_508) );
NOR2xp33_ASAP7_75t_R g509 ( .A(n_457), .B(n_449), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_492), .B(n_452), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_472), .B(n_416), .Y(n_511) );
NOR2xp33_ASAP7_75t_R g512 ( .A(n_491), .B(n_449), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_462), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_478), .B(n_449), .Y(n_514) );
NOR3xp33_ASAP7_75t_SL g515 ( .A(n_461), .B(n_24), .C(n_25), .Y(n_515) );
INVx2_ASAP7_75t_SL g516 ( .A(n_475), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_481), .B(n_444), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_465), .B(n_444), .Y(n_518) );
INVxp67_ASAP7_75t_L g519 ( .A(n_481), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_465), .B(n_444), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_490), .B(n_444), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_476), .B(n_214), .Y(n_522) );
NOR4xp25_ASAP7_75t_SL g523 ( .A(n_480), .B(n_27), .C(n_28), .D(n_29), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_456), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_490), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_470), .B(n_326), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_468), .B(n_453), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_464), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_475), .Y(n_529) );
NAND2x1p5_ASAP7_75t_L g530 ( .A(n_469), .B(n_326), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_468), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_458), .Y(n_532) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_464), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_472), .B(n_180), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_466), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_458), .B(n_349), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_466), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_453), .B(n_348), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_454), .B(n_328), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_467), .B(n_349), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_454), .A2(n_328), .B1(n_307), .B2(n_180), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_467), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_485), .B(n_191), .Y(n_543) );
CKINVDCx16_ASAP7_75t_R g544 ( .A(n_484), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_479), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_460), .B(n_191), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_460), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_493), .B(n_191), .Y(n_548) );
INVxp67_ASAP7_75t_SL g549 ( .A(n_533), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_506), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_504), .A2(n_471), .B1(n_469), .B2(n_473), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_529), .B(n_460), .Y(n_552) );
NAND2xp33_ASAP7_75t_L g553 ( .A(n_498), .B(n_486), .Y(n_553) );
AOI221x1_ASAP7_75t_L g554 ( .A1(n_545), .A2(n_451), .B1(n_488), .B2(n_495), .C(n_487), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_516), .B(n_473), .Y(n_555) );
NOR3xp33_ASAP7_75t_L g556 ( .A(n_544), .B(n_482), .C(n_494), .Y(n_556) );
AOI322xp5_ASAP7_75t_L g557 ( .A1(n_519), .A2(n_483), .A3(n_487), .B1(n_463), .B2(n_180), .C1(n_190), .C2(n_191), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_531), .B(n_487), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_504), .A2(n_487), .B1(n_304), .B2(n_260), .Y(n_559) );
NAND3x1_ASAP7_75t_SL g560 ( .A(n_501), .B(n_34), .C(n_38), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_513), .Y(n_561) );
XOR2xp5_ASAP7_75t_L g562 ( .A(n_516), .B(n_39), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_510), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_532), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_527), .B(n_190), .Y(n_565) );
OAI221xp5_ASAP7_75t_L g566 ( .A1(n_502), .A2(n_180), .B1(n_190), .B2(n_184), .C(n_304), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_511), .B(n_190), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_535), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_496), .B(n_41), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_501), .B(n_43), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_514), .B(n_44), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_507), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_522), .A2(n_304), .B1(n_289), .B2(n_184), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_535), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_520), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_525), .B(n_45), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_517), .B(n_184), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_538), .B(n_49), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_497), .A2(n_304), .B1(n_249), .B2(n_346), .Y(n_579) );
A2O1A1Ixp33_ASAP7_75t_L g580 ( .A1(n_515), .A2(n_184), .B(n_337), .C(n_54), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_511), .B(n_184), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_520), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_520), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_508), .B(n_521), .Y(n_584) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_507), .Y(n_585) );
OAI22xp33_ASAP7_75t_SL g586 ( .A1(n_497), .A2(n_184), .B1(n_53), .B2(n_55), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_503), .A2(n_289), .B1(n_297), .B2(n_276), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_537), .Y(n_588) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_509), .Y(n_589) );
AOI22xp5_ASAP7_75t_SL g590 ( .A1(n_498), .A2(n_530), .B1(n_512), .B2(n_509), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_512), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_542), .Y(n_592) );
OAI31xp33_ASAP7_75t_L g593 ( .A1(n_530), .A2(n_297), .A3(n_276), .B(n_265), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_508), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_508), .Y(n_595) );
CKINVDCx14_ASAP7_75t_R g596 ( .A(n_526), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_584), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_563), .B(n_518), .Y(n_598) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_549), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_550), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_575), .Y(n_601) );
INVx4_ASAP7_75t_L g602 ( .A(n_570), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_561), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_572), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_564), .B(n_539), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_588), .Y(n_606) );
AND2x2_ASAP7_75t_SL g607 ( .A(n_585), .B(n_503), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_592), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_582), .B(n_534), .Y(n_609) );
NAND4xp25_ASAP7_75t_L g610 ( .A(n_556), .B(n_541), .C(n_536), .D(n_548), .Y(n_610) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_596), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_568), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_583), .B(n_499), .Y(n_613) );
INVxp67_ASAP7_75t_L g614 ( .A(n_572), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_589), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_555), .B(n_499), .Y(n_616) );
XOR2x2_ASAP7_75t_L g617 ( .A(n_562), .B(n_500), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_574), .B(n_547), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_567), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_567), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_565), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_558), .B(n_528), .Y(n_622) );
AOI21xp33_ASAP7_75t_L g623 ( .A1(n_578), .A2(n_540), .B(n_546), .Y(n_623) );
AOI21xp33_ASAP7_75t_L g624 ( .A1(n_586), .A2(n_546), .B(n_528), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_595), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_552), .B(n_524), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_590), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_581), .B(n_524), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_581), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_594), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_577), .B(n_505), .Y(n_631) );
INVx2_ASAP7_75t_SL g632 ( .A(n_611), .Y(n_632) );
INVx2_ASAP7_75t_SL g633 ( .A(n_599), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_598), .B(n_551), .Y(n_634) );
NAND4xp75_ASAP7_75t_L g635 ( .A(n_607), .B(n_554), .C(n_571), .D(n_587), .Y(n_635) );
OAI32xp33_ASAP7_75t_L g636 ( .A1(n_627), .A2(n_591), .A3(n_569), .B1(n_559), .B2(n_566), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_619), .B(n_557), .Y(n_637) );
AO22x2_ASAP7_75t_L g638 ( .A1(n_615), .A2(n_591), .B1(n_559), .B2(n_570), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_604), .B(n_573), .Y(n_639) );
OAI21xp5_ASAP7_75t_SL g640 ( .A1(n_624), .A2(n_580), .B(n_593), .Y(n_640) );
XNOR2x1_ASAP7_75t_L g641 ( .A(n_617), .B(n_576), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_603), .Y(n_642) );
NOR2xp67_ASAP7_75t_L g643 ( .A(n_602), .B(n_579), .Y(n_643) );
NOR3xp33_ASAP7_75t_L g644 ( .A(n_610), .B(n_560), .C(n_553), .Y(n_644) );
XOR2x2_ASAP7_75t_L g645 ( .A(n_617), .B(n_579), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_602), .A2(n_523), .B1(n_543), .B2(n_243), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_603), .Y(n_647) );
NAND4xp25_ASAP7_75t_SL g648 ( .A(n_607), .B(n_543), .C(n_57), .D(n_58), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_614), .B(n_51), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_600), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_645), .A2(n_602), .B1(n_629), .B2(n_597), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_634), .A2(n_608), .B1(n_606), .B2(n_605), .C(n_612), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_634), .B(n_622), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_637), .B(n_619), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_644), .A2(n_623), .B1(n_620), .B2(n_621), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_633), .B(n_620), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_638), .A2(n_616), .B1(n_601), .B2(n_625), .C(n_626), .Y(n_657) );
A2O1A1Ixp33_ASAP7_75t_SL g658 ( .A1(n_649), .A2(n_601), .B(n_630), .C(n_631), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_641), .A2(n_609), .B1(n_618), .B2(n_622), .Y(n_659) );
OAI211xp5_ASAP7_75t_L g660 ( .A1(n_636), .A2(n_628), .B(n_613), .C(n_618), .Y(n_660) );
INVx1_ASAP7_75t_SL g661 ( .A(n_632), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_642), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_643), .A2(n_243), .B1(n_248), .B2(n_246), .Y(n_663) );
OAI211xp5_ASAP7_75t_L g664 ( .A1(n_640), .A2(n_250), .B(n_69), .C(n_72), .Y(n_664) );
NOR4xp75_ASAP7_75t_L g665 ( .A(n_635), .B(n_63), .C(n_646), .D(n_638), .Y(n_665) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_647), .Y(n_666) );
AOI322xp5_ASAP7_75t_L g667 ( .A1(n_639), .A2(n_632), .A3(n_627), .B1(n_611), .B2(n_634), .C1(n_644), .C2(n_637), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_646), .B(n_650), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_653), .Y(n_669) );
NOR3xp33_ASAP7_75t_SL g670 ( .A(n_664), .B(n_660), .C(n_668), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_662), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_654), .B(n_662), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_651), .B(n_661), .Y(n_673) );
NOR2x1_ASAP7_75t_L g674 ( .A(n_673), .B(n_648), .Y(n_674) );
OR3x1_ASAP7_75t_L g675 ( .A(n_669), .B(n_667), .C(n_665), .Y(n_675) );
XNOR2xp5_ASAP7_75t_L g676 ( .A(n_670), .B(n_655), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_676), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_674), .B(n_671), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_678), .Y(n_679) );
NAND2x2_ASAP7_75t_L g680 ( .A(n_677), .B(n_675), .Y(n_680) );
AOI322xp5_ASAP7_75t_L g681 ( .A1(n_679), .A2(n_670), .A3(n_657), .B1(n_659), .B2(n_652), .C1(n_656), .C2(n_666), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_681), .A2(n_680), .B1(n_663), .B2(n_672), .C(n_658), .Y(n_682) );
endmodule