module fake_jpeg_1235_n_153 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_55),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_58),
.B(n_59),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_54),
.C(n_48),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_46),
.Y(n_75)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_49),
.B1(n_60),
.B2(n_59),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_70),
.B1(n_57),
.B2(n_50),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_51),
.B1(n_40),
.B2(n_50),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_39),
.C(n_42),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_67),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_79),
.Y(n_92)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_45),
.A3(n_47),
.B1(n_39),
.B2(n_38),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_42),
.B(n_2),
.Y(n_99)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_72),
.B(n_52),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_86),
.Y(n_90)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_13),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_56),
.B1(n_64),
.B2(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_63),
.B1(n_62),
.B2(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_53),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_87),
.A2(n_62),
.B1(n_63),
.B2(n_56),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_0),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_97),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_37),
.C(n_30),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_1),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_83),
.B1(n_78),
.B2(n_19),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_102),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_79),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_4),
.Y(n_118)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_95),
.B(n_1),
.CI(n_3),
.CON(n_106),
.SN(n_106)
);

AOI32xp33_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_108),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_127)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_109),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_21),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_117),
.C(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_115),
.B(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_14),
.C(n_34),
.Y(n_117)
);

NOR4xp25_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_7),
.C(n_9),
.D(n_10),
.Y(n_132)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_24),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_108),
.A2(n_100),
.B(n_5),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_127),
.B(n_133),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_131),
.B1(n_117),
.B2(n_12),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_25),
.B(n_26),
.C(n_27),
.D(n_28),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_10),
.B(n_11),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_140),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_137),
.A2(n_129),
.B(n_134),
.Y(n_141)
);

AOI31xp67_ASAP7_75t_L g146 ( 
.A1(n_141),
.A2(n_142),
.A3(n_143),
.B(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_136),
.B(n_131),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_124),
.C(n_130),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_145),
.A2(n_146),
.B(n_122),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_123),
.B(n_139),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_137),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_128),
.B1(n_111),
.B2(n_29),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g151 ( 
.A(n_150),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_111),
.Y(n_153)
);


endmodule