module real_aes_10848_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_1380;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_399;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_1404;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1620;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1638;
wire n_495;
wire n_1072;
wire n_1078;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_729;
wire n_1323;
wire n_1352;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AO221x1_ASAP7_75t_L g712 ( .A1(n_0), .A2(n_173), .B1(n_713), .B2(n_720), .C(n_723), .Y(n_712) );
OAI222xp33_ASAP7_75t_L g1238 ( .A1(n_1), .A2(n_42), .B1(n_176), .B2(n_1239), .C1(n_1241), .C2(n_1243), .Y(n_1238) );
AOI221xp5_ASAP7_75t_L g1269 ( .A1(n_1), .A2(n_176), .B1(n_1270), .B2(n_1271), .C(n_1273), .Y(n_1269) );
AOI22xp33_ASAP7_75t_L g1286 ( .A1(n_2), .A2(n_14), .B1(n_451), .B2(n_659), .Y(n_1286) );
OAI22xp5_ASAP7_75t_L g1320 ( .A1(n_2), .A2(n_14), .B1(n_593), .B2(n_698), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_3), .B(n_219), .Y(n_377) );
AND2x2_ASAP7_75t_L g394 ( .A(n_3), .B(n_395), .Y(n_394) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_3), .Y(n_431) );
INVx1_ASAP7_75t_L g464 ( .A(n_3), .Y(n_464) );
INVx1_ASAP7_75t_L g637 ( .A(n_4), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_4), .A2(n_212), .B1(n_675), .B2(n_676), .Y(n_674) );
INVx1_ASAP7_75t_L g1437 ( .A(n_5), .Y(n_1437) );
AOI22xp33_ASAP7_75t_L g1464 ( .A1(n_5), .A2(n_87), .B1(n_1465), .B2(n_1466), .Y(n_1464) );
AOI22xp33_ASAP7_75t_SL g662 ( .A1(n_6), .A2(n_54), .B1(n_658), .B2(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g702 ( .A(n_6), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_7), .A2(n_121), .B1(n_713), .B2(n_722), .Y(n_752) );
OAI21xp33_ASAP7_75t_SL g940 ( .A1(n_8), .A2(n_941), .B(n_944), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_8), .A2(n_130), .B1(n_1013), .B2(n_1014), .Y(n_1012) );
CKINVDCx5p33_ASAP7_75t_R g1499 ( .A(n_9), .Y(n_1499) );
OAI221xp5_ASAP7_75t_L g1433 ( .A1(n_10), .A2(n_240), .B1(n_422), .B2(n_1336), .C(n_1434), .Y(n_1433) );
OAI22xp33_ASAP7_75t_L g1456 ( .A1(n_10), .A2(n_240), .B1(n_675), .B2(n_676), .Y(n_1456) );
CKINVDCx5p33_ASAP7_75t_R g1395 ( .A(n_11), .Y(n_1395) );
AOI221xp5_ASAP7_75t_L g1052 ( .A1(n_12), .A2(n_108), .B1(n_496), .B2(n_1053), .C(n_1054), .Y(n_1052) );
AOI22xp33_ASAP7_75t_SL g1075 ( .A1(n_12), .A2(n_161), .B1(n_1076), .B2(n_1077), .Y(n_1075) );
INVx1_ASAP7_75t_L g1540 ( .A(n_13), .Y(n_1540) );
INVx1_ASAP7_75t_L g950 ( .A(n_15), .Y(n_950) );
OAI222xp33_ASAP7_75t_L g978 ( .A1(n_15), .A2(n_26), .B1(n_270), .B2(n_519), .C1(n_979), .C2(n_981), .Y(n_978) );
INVx1_ASAP7_75t_L g484 ( .A(n_16), .Y(n_484) );
INVx1_ASAP7_75t_L g1439 ( .A(n_17), .Y(n_1439) );
AOI221xp5_ASAP7_75t_L g1463 ( .A1(n_17), .A2(n_248), .B1(n_688), .B2(n_690), .C(n_1370), .Y(n_1463) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_18), .A2(n_110), .B1(n_348), .B2(n_350), .Y(n_347) );
INVxp67_ASAP7_75t_SL g449 ( .A(n_18), .Y(n_449) );
INVxp33_ASAP7_75t_L g1172 ( .A(n_19), .Y(n_1172) );
AOI221xp5_ASAP7_75t_L g1210 ( .A1(n_19), .A2(n_156), .B1(n_601), .B2(n_602), .C(n_1211), .Y(n_1210) );
INVx1_ASAP7_75t_L g358 ( .A(n_20), .Y(n_358) );
AO221x2_ASAP7_75t_L g806 ( .A1(n_21), .A2(n_192), .B1(n_720), .B2(n_807), .C(n_809), .Y(n_806) );
OAI221xp5_ASAP7_75t_L g1335 ( .A1(n_22), .A2(n_190), .B1(n_426), .B2(n_527), .C(n_1336), .Y(n_1335) );
OAI22xp5_ASAP7_75t_L g1364 ( .A1(n_22), .A2(n_190), .B1(n_1365), .B2(n_1366), .Y(n_1364) );
INVx1_ASAP7_75t_L g1396 ( .A(n_23), .Y(n_1396) );
CKINVDCx5p33_ASAP7_75t_R g1483 ( .A(n_24), .Y(n_1483) );
INVx1_ASAP7_75t_L g606 ( .A(n_25), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g1026 ( .A1(n_26), .A2(n_196), .B1(n_301), .B2(n_1021), .Y(n_1026) );
INVx2_ASAP7_75t_L g310 ( .A(n_27), .Y(n_310) );
OR2x2_ASAP7_75t_L g323 ( .A(n_27), .B(n_324), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_28), .A2(n_111), .B1(n_334), .B2(n_476), .Y(n_475) );
OAI221xp5_ASAP7_75t_L g526 ( .A1(n_28), .A2(n_111), .B1(n_415), .B2(n_426), .C(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g1218 ( .A(n_29), .Y(n_1218) );
AOI221xp5_ASAP7_75t_L g1125 ( .A1(n_30), .A2(n_47), .B1(n_1025), .B2(n_1126), .C(n_1127), .Y(n_1125) );
INVx1_ASAP7_75t_L g1158 ( .A(n_30), .Y(n_1158) );
INVx1_ASAP7_75t_L g1428 ( .A(n_31), .Y(n_1428) );
AOI221xp5_ASAP7_75t_L g1457 ( .A1(n_31), .A2(n_141), .B1(n_350), .B2(n_1458), .C(n_1460), .Y(n_1457) );
CKINVDCx5p33_ASAP7_75t_R g1503 ( .A(n_32), .Y(n_1503) );
INVx1_ASAP7_75t_L g353 ( .A(n_33), .Y(n_353) );
AOI22xp33_ASAP7_75t_SL g312 ( .A1(n_34), .A2(n_153), .B1(n_313), .B2(n_317), .Y(n_312) );
INVxp33_ASAP7_75t_SL g407 ( .A(n_34), .Y(n_407) );
BUFx2_ASAP7_75t_L g292 ( .A(n_35), .Y(n_292) );
OR2x2_ASAP7_75t_L g376 ( .A(n_35), .B(n_377), .Y(n_376) );
BUFx2_ASAP7_75t_L g380 ( .A(n_35), .Y(n_380) );
INVx1_ASAP7_75t_L g393 ( .A(n_35), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g1384 ( .A1(n_36), .A2(n_44), .B1(n_1211), .B2(n_1385), .C(n_1386), .Y(n_1384) );
INVx1_ASAP7_75t_L g1404 ( .A(n_36), .Y(n_1404) );
INVx1_ASAP7_75t_L g505 ( .A(n_37), .Y(n_505) );
INVx1_ASAP7_75t_L g1348 ( .A(n_38), .Y(n_1348) );
INVx1_ASAP7_75t_L g1490 ( .A(n_39), .Y(n_1490) );
AOI221xp5_ASAP7_75t_SL g1508 ( .A1(n_39), .A2(n_178), .B1(n_344), .B2(n_1509), .C(n_1511), .Y(n_1508) );
INVx1_ASAP7_75t_L g957 ( .A(n_40), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g973 ( .A1(n_40), .A2(n_196), .B1(n_974), .B2(n_976), .Y(n_973) );
AOI22xp33_ASAP7_75t_SL g1287 ( .A1(n_41), .A2(n_84), .B1(n_655), .B2(n_1283), .Y(n_1287) );
INVx1_ASAP7_75t_L g1319 ( .A(n_41), .Y(n_1319) );
INVx1_ASAP7_75t_L g1274 ( .A(n_42), .Y(n_1274) );
INVx1_ASAP7_75t_L g1484 ( .A(n_43), .Y(n_1484) );
AOI221xp5_ASAP7_75t_L g1522 ( .A1(n_43), .A2(n_170), .B1(n_1523), .B2(n_1525), .C(n_1528), .Y(n_1522) );
INVx1_ASAP7_75t_L g1402 ( .A(n_44), .Y(n_1402) );
INVx1_ASAP7_75t_L g1191 ( .A(n_45), .Y(n_1191) );
AOI22xp33_ASAP7_75t_SL g1282 ( .A1(n_46), .A2(n_229), .B1(n_655), .B2(n_1283), .Y(n_1282) );
AOI22xp33_ASAP7_75t_L g1307 ( .A1(n_46), .A2(n_189), .B1(n_1208), .B2(n_1308), .Y(n_1307) );
INVx1_ASAP7_75t_L g1161 ( .A(n_47), .Y(n_1161) );
INVx1_ASAP7_75t_L g1141 ( .A(n_48), .Y(n_1141) );
INVx1_ASAP7_75t_L g729 ( .A(n_49), .Y(n_729) );
INVx1_ASAP7_75t_L g364 ( .A(n_50), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g1481 ( .A(n_51), .Y(n_1481) );
INVx1_ASAP7_75t_L g1496 ( .A(n_52), .Y(n_1496) );
AOI22xp33_ASAP7_75t_L g1513 ( .A1(n_52), .A2(n_60), .B1(n_1514), .B2(n_1515), .Y(n_1513) );
INVxp67_ASAP7_75t_SL g1060 ( .A(n_53), .Y(n_1060) );
AOI221xp5_ASAP7_75t_L g1095 ( .A1(n_53), .A2(n_105), .B1(n_1096), .B2(n_1098), .C(n_1099), .Y(n_1095) );
INVx1_ASAP7_75t_L g673 ( .A(n_54), .Y(n_673) );
INVxp67_ASAP7_75t_L g1330 ( .A(n_55), .Y(n_1330) );
AOI221xp5_ASAP7_75t_L g1362 ( .A1(n_55), .A2(n_157), .B1(n_296), .B2(n_307), .C(n_1130), .Y(n_1362) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_56), .A2(n_215), .B1(n_498), .B2(n_501), .Y(n_497) );
INVxp67_ASAP7_75t_SL g513 ( .A(n_56), .Y(n_513) );
INVxp67_ASAP7_75t_SL g1064 ( .A(n_57), .Y(n_1064) );
OAI211xp5_ASAP7_75t_SL g1081 ( .A1(n_57), .A2(n_1082), .B(n_1085), .C(n_1089), .Y(n_1081) );
INVx1_ASAP7_75t_L g1067 ( .A(n_58), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1567 ( .A1(n_59), .A2(n_78), .B1(n_1526), .B2(n_1568), .Y(n_1567) );
INVxp67_ASAP7_75t_L g1616 ( .A(n_59), .Y(n_1616) );
INVx1_ASAP7_75t_L g1488 ( .A(n_60), .Y(n_1488) );
INVx1_ASAP7_75t_L g493 ( .A(n_61), .Y(n_493) );
XNOR2x2_ASAP7_75t_L g1275 ( .A(n_62), .B(n_1276), .Y(n_1275) );
INVxp33_ASAP7_75t_L g1339 ( .A(n_63), .Y(n_1339) );
AOI22xp33_ASAP7_75t_L g1371 ( .A1(n_63), .A2(n_233), .B1(n_580), .B2(n_601), .Y(n_1371) );
OAI222xp33_ASAP7_75t_L g1245 ( .A1(n_64), .A2(n_150), .B1(n_228), .B2(n_1066), .C1(n_1216), .C2(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1251 ( .A(n_64), .Y(n_1251) );
CKINVDCx5p33_ASAP7_75t_R g1296 ( .A(n_65), .Y(n_1296) );
CKINVDCx5p33_ASAP7_75t_R g1451 ( .A(n_66), .Y(n_1451) );
AOI221xp5_ASAP7_75t_L g477 ( .A1(n_67), .A2(n_238), .B1(n_350), .B2(n_478), .C(n_481), .Y(n_477) );
INVxp33_ASAP7_75t_L g533 ( .A(n_67), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g1284 ( .A1(n_68), .A2(n_189), .B1(n_1098), .B2(n_1285), .Y(n_1284) );
AOI21xp33_ASAP7_75t_L g1309 ( .A1(n_68), .A2(n_590), .B(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g471 ( .A(n_69), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_70), .A2(n_227), .B1(n_997), .B2(n_999), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_70), .A2(n_241), .B1(n_1020), .B2(n_1021), .Y(n_1019) );
INVxp33_ASAP7_75t_SL g543 ( .A(n_71), .Y(n_543) );
AOI221xp5_ASAP7_75t_L g591 ( .A1(n_71), .A2(n_265), .B1(n_580), .B2(n_592), .C(n_595), .Y(n_591) );
AOI22xp33_ASAP7_75t_SL g1049 ( .A1(n_72), .A2(n_161), .B1(n_301), .B2(n_1050), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_72), .A2(n_108), .B1(n_1009), .B2(n_1080), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_73), .A2(n_96), .B1(n_501), .B2(n_1056), .Y(n_1229) );
INVx1_ASAP7_75t_L g1256 ( .A(n_73), .Y(n_1256) );
INVx1_ASAP7_75t_L g730 ( .A(n_74), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_75), .A2(n_149), .B1(n_317), .B2(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1267 ( .A(n_75), .Y(n_1267) );
AOI22xp5_ASAP7_75t_L g1423 ( .A1(n_76), .A2(n_1424), .B1(n_1470), .B2(n_1471), .Y(n_1423) );
INVx1_ASAP7_75t_L g1470 ( .A(n_76), .Y(n_1470) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_77), .A2(n_232), .B1(n_654), .B2(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g686 ( .A(n_77), .Y(n_686) );
INVxp67_ASAP7_75t_L g1614 ( .A(n_78), .Y(n_1614) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_79), .A2(n_101), .B1(n_1050), .B2(n_1056), .Y(n_1055) );
INVxp67_ASAP7_75t_SL g1104 ( .A(n_79), .Y(n_1104) );
INVx1_ASAP7_75t_L g646 ( .A(n_80), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_80), .A2(n_104), .B1(n_313), .B2(n_580), .C(n_679), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g1057 ( .A1(n_81), .A2(n_163), .B1(n_301), .B2(n_307), .C(n_1021), .Y(n_1057) );
INVxp33_ASAP7_75t_SL g1092 ( .A(n_81), .Y(n_1092) );
CKINVDCx5p33_ASAP7_75t_R g645 ( .A(n_82), .Y(n_645) );
AO221x1_ASAP7_75t_L g760 ( .A1(n_83), .A2(n_126), .B1(n_713), .B2(n_722), .C(n_761), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g1302 ( .A(n_84), .B(n_360), .Y(n_1302) );
INVx1_ASAP7_75t_L g812 ( .A(n_85), .Y(n_812) );
INVx1_ASAP7_75t_L g1299 ( .A(n_86), .Y(n_1299) );
AOI22xp33_ASAP7_75t_L g1314 ( .A1(n_86), .A2(n_140), .B1(n_1308), .B2(n_1310), .Y(n_1314) );
INVx1_ASAP7_75t_L g1445 ( .A(n_87), .Y(n_1445) );
AO221x1_ASAP7_75t_L g755 ( .A1(n_88), .A2(n_185), .B1(n_713), .B2(n_722), .C(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g758 ( .A(n_89), .Y(n_758) );
INVx1_ASAP7_75t_L g311 ( .A(n_90), .Y(n_311) );
INVx1_ASAP7_75t_L g324 ( .A(n_90), .Y(n_324) );
INVx1_ASAP7_75t_L g465 ( .A(n_91), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g1500 ( .A(n_92), .Y(n_1500) );
INVx1_ASAP7_75t_L g1357 ( .A(n_93), .Y(n_1357) );
INVx1_ASAP7_75t_L g1291 ( .A(n_94), .Y(n_1291) );
AOI21xp5_ASAP7_75t_L g1315 ( .A1(n_94), .A2(n_489), .B(n_583), .Y(n_1315) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_95), .A2(n_276), .B1(n_327), .B2(n_676), .Y(n_1124) );
INVx1_ASAP7_75t_L g1145 ( .A(n_95), .Y(n_1145) );
INVx1_ASAP7_75t_L g1253 ( .A(n_96), .Y(n_1253) );
INVx1_ASAP7_75t_L g1556 ( .A(n_97), .Y(n_1556) );
INVxp67_ASAP7_75t_SL g1182 ( .A(n_98), .Y(n_1182) );
AOI221xp5_ASAP7_75t_L g1204 ( .A1(n_98), .A2(n_224), .B1(n_344), .B2(n_496), .C(n_1202), .Y(n_1204) );
CKINVDCx5p33_ASAP7_75t_R g1431 ( .A(n_99), .Y(n_1431) );
INVxp33_ASAP7_75t_SL g1169 ( .A(n_100), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g1212 ( .A1(n_100), .A2(n_122), .B1(n_495), .B2(n_613), .Y(n_1212) );
INVxp33_ASAP7_75t_L g1093 ( .A(n_101), .Y(n_1093) );
INVxp67_ASAP7_75t_L g1334 ( .A(n_102), .Y(n_1334) );
AOI22xp33_ASAP7_75t_L g1363 ( .A1(n_102), .A2(n_204), .B1(n_1025), .B2(n_1242), .Y(n_1363) );
AOI221xp5_ASAP7_75t_L g1391 ( .A1(n_103), .A2(n_168), .B1(n_344), .B2(n_602), .C(n_1392), .Y(n_1391) );
INVx1_ASAP7_75t_L g1413 ( .A(n_103), .Y(n_1413) );
INVx1_ASAP7_75t_L g641 ( .A(n_104), .Y(n_641) );
OAI211xp5_ASAP7_75t_SL g1047 ( .A1(n_105), .A2(n_366), .B(n_1048), .C(n_1058), .Y(n_1047) );
CKINVDCx5p33_ASAP7_75t_R g1429 ( .A(n_106), .Y(n_1429) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_107), .A2(n_236), .B1(n_713), .B2(n_722), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_109), .A2(n_137), .B1(n_965), .B2(n_967), .Y(n_964) );
AOI22xp33_ASAP7_75t_SL g1008 ( .A1(n_109), .A2(n_137), .B1(n_1009), .B2(n_1010), .Y(n_1008) );
INVxp33_ASAP7_75t_L g434 ( .A(n_110), .Y(n_434) );
OAI221xp5_ASAP7_75t_L g1485 ( .A1(n_112), .A2(n_147), .B1(n_415), .B2(n_426), .C(n_527), .Y(n_1485) );
OAI22xp5_ASAP7_75t_L g1518 ( .A1(n_112), .A2(n_147), .B1(n_1519), .B2(n_1520), .Y(n_1518) );
INVx1_ASAP7_75t_L g325 ( .A(n_113), .Y(n_325) );
INVx1_ASAP7_75t_L g1374 ( .A(n_114), .Y(n_1374) );
INVxp33_ASAP7_75t_SL g1548 ( .A(n_115), .Y(n_1548) );
AOI221xp5_ASAP7_75t_L g1601 ( .A1(n_115), .A2(n_274), .B1(n_665), .B2(n_1602), .C(n_1604), .Y(n_1601) );
INVx1_ASAP7_75t_L g763 ( .A(n_116), .Y(n_763) );
INVx1_ASAP7_75t_L g1188 ( .A(n_117), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g1205 ( .A1(n_117), .A2(n_188), .B1(n_317), .B2(n_1206), .Y(n_1205) );
CKINVDCx5p33_ASAP7_75t_R g1383 ( .A(n_118), .Y(n_1383) );
OAI22xp33_ASAP7_75t_L g1389 ( .A1(n_119), .A2(n_250), .B1(n_1216), .B2(n_1365), .Y(n_1389) );
OAI221xp5_ASAP7_75t_L g1407 ( .A1(n_119), .A2(n_250), .B1(n_527), .B2(n_1175), .C(n_1408), .Y(n_1407) );
INVx1_ASAP7_75t_L g718 ( .A(n_120), .Y(n_718) );
INVxp33_ASAP7_75t_SL g1173 ( .A(n_122), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1569 ( .A1(n_123), .A2(n_205), .B1(n_1465), .B2(n_1570), .Y(n_1569) );
INVxp67_ASAP7_75t_SL g1623 ( .A(n_123), .Y(n_1623) );
INVx1_ASAP7_75t_L g562 ( .A(n_124), .Y(n_562) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_124), .A2(n_223), .B1(n_580), .B2(n_581), .C(n_584), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_125), .A2(n_221), .B1(n_739), .B2(n_742), .Y(n_747) );
INVx1_ASAP7_75t_L g762 ( .A(n_127), .Y(n_762) );
INVx1_ASAP7_75t_L g1134 ( .A(n_128), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_128), .A2(n_180), .B1(n_665), .B2(n_1156), .Y(n_1155) );
AOI22xp5_ASAP7_75t_L g1044 ( .A1(n_129), .A2(n_1045), .B1(n_1105), .B2(n_1106), .Y(n_1044) );
CKINVDCx5p33_ASAP7_75t_R g1105 ( .A(n_129), .Y(n_1105) );
INVxp67_ASAP7_75t_SL g961 ( .A(n_130), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_131), .A2(n_159), .B1(n_658), .B2(n_660), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_131), .A2(n_220), .B1(n_590), .B2(n_688), .C(n_690), .Y(n_687) );
CKINVDCx5p33_ASAP7_75t_R g1447 ( .A(n_132), .Y(n_1447) );
INVx1_ASAP7_75t_L g607 ( .A(n_133), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_134), .A2(n_200), .B1(n_713), .B2(n_722), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_135), .A2(n_279), .B1(n_739), .B2(n_742), .Y(n_772) );
AOI221xp5_ASAP7_75t_L g1230 ( .A1(n_136), .A2(n_198), .B1(n_590), .B2(n_602), .C(n_1231), .Y(n_1230) );
AOI221xp5_ASAP7_75t_L g1263 ( .A1(n_136), .A2(n_149), .B1(n_1002), .B2(n_1264), .C(n_1266), .Y(n_1263) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_138), .A2(n_253), .B1(n_498), .B2(n_501), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1150 ( .A1(n_138), .A2(n_154), .B1(n_454), .B2(n_1076), .Y(n_1150) );
INVx1_ASAP7_75t_L g1162 ( .A(n_139), .Y(n_1162) );
INVx1_ASAP7_75t_L g1295 ( .A(n_140), .Y(n_1295) );
INVx1_ASAP7_75t_L g1432 ( .A(n_141), .Y(n_1432) );
XNOR2x1_ASAP7_75t_L g1475 ( .A(n_142), .B(n_1476), .Y(n_1475) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_143), .A2(n_206), .B1(n_327), .B2(n_334), .Y(n_326) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_143), .A2(n_206), .B1(n_415), .B2(n_422), .C(n_426), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g1450 ( .A(n_144), .Y(n_1450) );
CKINVDCx5p33_ASAP7_75t_R g1505 ( .A(n_145), .Y(n_1505) );
AOI221xp5_ASAP7_75t_L g1226 ( .A1(n_146), .A2(n_165), .B1(n_307), .B2(n_1227), .C(n_1228), .Y(n_1226) );
INVx1_ASAP7_75t_L g1254 ( .A(n_146), .Y(n_1254) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_148), .A2(n_220), .B1(n_654), .B2(n_655), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_148), .A2(n_159), .B1(n_695), .B2(n_697), .Y(n_694) );
INVx1_ASAP7_75t_L g1258 ( .A(n_150), .Y(n_1258) );
INVx1_ASAP7_75t_L g810 ( .A(n_151), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_152), .A2(n_241), .B1(n_1002), .B2(n_1004), .Y(n_1001) );
AOI22xp33_ASAP7_75t_SL g1023 ( .A1(n_152), .A2(n_227), .B1(n_1024), .B2(n_1025), .Y(n_1023) );
INVxp33_ASAP7_75t_L g385 ( .A(n_153), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g1135 ( .A1(n_154), .A2(n_162), .B1(n_590), .B2(n_1053), .C(n_1136), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_155), .A2(n_231), .B1(n_404), .B2(n_576), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_155), .A2(n_249), .B1(n_610), .B2(n_612), .Y(n_609) );
INVxp33_ASAP7_75t_L g1170 ( .A(n_156), .Y(n_1170) );
INVxp67_ASAP7_75t_L g1333 ( .A(n_157), .Y(n_1333) );
CKINVDCx5p33_ASAP7_75t_R g1502 ( .A(n_158), .Y(n_1502) );
CKINVDCx5p33_ASAP7_75t_R g1279 ( .A(n_160), .Y(n_1279) );
AOI22xp33_ASAP7_75t_SL g1147 ( .A1(n_162), .A2(n_253), .B1(n_1148), .B2(n_1149), .Y(n_1147) );
OAI21xp33_ASAP7_75t_SL g1072 ( .A1(n_163), .A2(n_1073), .B(n_1074), .Y(n_1072) );
INVx1_ASAP7_75t_L g1140 ( .A(n_164), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_164), .A2(n_197), .B1(n_1076), .B2(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1262 ( .A(n_165), .Y(n_1262) );
CKINVDCx5p33_ASAP7_75t_R g1237 ( .A(n_166), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g1387 ( .A1(n_167), .A2(n_202), .B1(n_1053), .B2(n_1388), .Y(n_1387) );
INVx1_ASAP7_75t_L g1401 ( .A(n_167), .Y(n_1401) );
INVx1_ASAP7_75t_L g1415 ( .A(n_168), .Y(n_1415) );
AOI22xp33_ASAP7_75t_L g1393 ( .A1(n_169), .A2(n_247), .B1(n_301), .B2(n_613), .Y(n_1393) );
INVx1_ASAP7_75t_L g1417 ( .A(n_169), .Y(n_1417) );
INVx1_ASAP7_75t_L g1480 ( .A(n_170), .Y(n_1480) );
INVx1_ASAP7_75t_L g1356 ( .A(n_171), .Y(n_1356) );
INVx1_ASAP7_75t_L g368 ( .A(n_172), .Y(n_368) );
XNOR2xp5_ASAP7_75t_L g1535 ( .A(n_173), .B(n_1536), .Y(n_1535) );
INVxp67_ASAP7_75t_L g1342 ( .A(n_174), .Y(n_1342) );
AOI221xp5_ASAP7_75t_L g1368 ( .A1(n_174), .A2(n_235), .B1(n_594), .B2(n_1369), .C(n_1370), .Y(n_1368) );
OAI221xp5_ASAP7_75t_L g1174 ( .A1(n_175), .A2(n_277), .B1(n_415), .B2(n_423), .C(n_1175), .Y(n_1174) );
OAI22xp33_ASAP7_75t_L g1213 ( .A1(n_175), .A2(n_277), .B1(n_1214), .B2(n_1216), .Y(n_1213) );
CKINVDCx5p33_ASAP7_75t_R g1380 ( .A(n_177), .Y(n_1380) );
INVx1_ASAP7_75t_L g1494 ( .A(n_178), .Y(n_1494) );
INVx1_ASAP7_75t_L g552 ( .A(n_179), .Y(n_552) );
INVx1_ASAP7_75t_L g1139 ( .A(n_180), .Y(n_1139) );
AOI22xp33_ASAP7_75t_SL g1572 ( .A1(n_181), .A2(n_243), .B1(n_1570), .B2(n_1573), .Y(n_1572) );
OAI221xp5_ASAP7_75t_L g1610 ( .A1(n_181), .A2(n_1611), .B1(n_1613), .B2(n_1621), .C(n_1626), .Y(n_1610) );
INVx1_ASAP7_75t_L g670 ( .A(n_182), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g1280 ( .A(n_183), .Y(n_1280) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_184), .A2(n_266), .B1(n_344), .B2(n_495), .C(n_496), .Y(n_494) );
INVxp33_ASAP7_75t_SL g516 ( .A(n_184), .Y(n_516) );
INVx1_ASAP7_75t_L g1164 ( .A(n_185), .Y(n_1164) );
INVx1_ASAP7_75t_L g474 ( .A(n_186), .Y(n_474) );
AND3x2_ASAP7_75t_L g717 ( .A(n_187), .B(n_718), .C(n_719), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_187), .B(n_718), .Y(n_726) );
HB1xp67_ASAP7_75t_L g1036 ( .A(n_187), .Y(n_1036) );
INVxp67_ASAP7_75t_SL g1181 ( .A(n_188), .Y(n_1181) );
INVx2_ASAP7_75t_L g375 ( .A(n_191), .Y(n_375) );
XOR2xp5_ASAP7_75t_L g468 ( .A(n_192), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g487 ( .A(n_193), .Y(n_487) );
XNOR2x2_ASAP7_75t_L g539 ( .A(n_194), .B(n_540), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g643 ( .A(n_195), .Y(n_643) );
INVx1_ASAP7_75t_L g1123 ( .A(n_197), .Y(n_1123) );
INVx1_ASAP7_75t_L g1268 ( .A(n_198), .Y(n_1268) );
AOI22xp5_ASAP7_75t_L g1575 ( .A1(n_199), .A2(n_244), .B1(n_1388), .B2(n_1576), .Y(n_1575) );
OAI22xp5_ASAP7_75t_L g1628 ( .A1(n_199), .A2(n_244), .B1(n_1629), .B2(n_1631), .Y(n_1628) );
INVxp67_ASAP7_75t_L g1324 ( .A(n_201), .Y(n_1324) );
INVx1_ASAP7_75t_L g1405 ( .A(n_202), .Y(n_1405) );
CKINVDCx5p33_ASAP7_75t_R g1453 ( .A(n_203), .Y(n_1453) );
INVxp67_ASAP7_75t_L g1329 ( .A(n_204), .Y(n_1329) );
INVxp67_ASAP7_75t_SL g1622 ( .A(n_205), .Y(n_1622) );
XNOR2xp5_ASAP7_75t_L g1375 ( .A(n_207), .B(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g719 ( .A(n_208), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g339 ( .A1(n_209), .A2(n_269), .B1(n_314), .B2(n_340), .C(n_344), .Y(n_339) );
INVxp67_ASAP7_75t_SL g443 ( .A(n_209), .Y(n_443) );
INVx1_ASAP7_75t_L g558 ( .A(n_210), .Y(n_558) );
INVx1_ASAP7_75t_L g545 ( .A(n_211), .Y(n_545) );
INVx1_ASAP7_75t_L g638 ( .A(n_212), .Y(n_638) );
OAI211xp5_ASAP7_75t_SL g1061 ( .A1(n_213), .A2(n_1062), .B(n_1063), .C(n_1069), .Y(n_1061) );
INVx1_ASAP7_75t_L g1102 ( .A(n_213), .Y(n_1102) );
INVxp33_ASAP7_75t_SL g988 ( .A(n_214), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_214), .A2(n_259), .B1(n_495), .B2(n_1025), .Y(n_1027) );
INVxp33_ASAP7_75t_L g515 ( .A(n_215), .Y(n_515) );
INVx1_ASAP7_75t_L g506 ( .A(n_216), .Y(n_506) );
INVx1_ASAP7_75t_L g1300 ( .A(n_217), .Y(n_1300) );
OAI211xp5_ASAP7_75t_L g1317 ( .A1(n_217), .A2(n_1066), .B(n_1318), .C(n_1321), .Y(n_1317) );
INVx1_ASAP7_75t_L g1194 ( .A(n_218), .Y(n_1194) );
INVx2_ASAP7_75t_L g395 ( .A(n_219), .Y(n_395) );
INVx1_ASAP7_75t_L g652 ( .A(n_219), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_222), .A2(n_239), .B1(n_739), .B2(n_742), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_223), .A2(n_225), .B1(n_564), .B2(n_567), .Y(n_563) );
INVxp67_ASAP7_75t_SL g1187 ( .A(n_224), .Y(n_1187) );
INVx1_ASAP7_75t_L g587 ( .A(n_225), .Y(n_587) );
INVx1_ASAP7_75t_L g757 ( .A(n_226), .Y(n_757) );
INVx1_ASAP7_75t_L g1250 ( .A(n_228), .Y(n_1250) );
INVx1_ASAP7_75t_L g1305 ( .A(n_229), .Y(n_1305) );
XOR2x1_ASAP7_75t_L g633 ( .A(n_230), .B(n_634), .Y(n_633) );
OAI22xp33_ASAP7_75t_L g614 ( .A1(n_231), .A2(n_258), .B1(n_615), .B2(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g701 ( .A(n_232), .Y(n_701) );
INVxp67_ASAP7_75t_L g1345 ( .A(n_233), .Y(n_1345) );
INVx1_ASAP7_75t_L g1192 ( .A(n_234), .Y(n_1192) );
INVxp33_ASAP7_75t_L g1340 ( .A(n_235), .Y(n_1340) );
INVx1_ASAP7_75t_L g1551 ( .A(n_237), .Y(n_1551) );
INVxp33_ASAP7_75t_L g530 ( .A(n_238), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g1448 ( .A(n_242), .Y(n_1448) );
OAI211xp5_ASAP7_75t_SL g1592 ( .A1(n_243), .A2(n_1593), .B(n_1597), .C(n_1605), .Y(n_1592) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_245), .A2(n_280), .B1(n_296), .B2(n_301), .C(n_307), .Y(n_295) );
INVxp33_ASAP7_75t_L g402 ( .A(n_245), .Y(n_402) );
INVx1_ASAP7_75t_L g716 ( .A(n_246), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_246), .B(n_728), .Y(n_733) );
INVx1_ASAP7_75t_L g1412 ( .A(n_247), .Y(n_1412) );
INVx1_ASAP7_75t_L g1441 ( .A(n_248), .Y(n_1441) );
INVxp67_ASAP7_75t_SL g574 ( .A(n_249), .Y(n_574) );
INVx1_ASAP7_75t_L g1068 ( .A(n_251), .Y(n_1068) );
INVx1_ASAP7_75t_L g1562 ( .A(n_252), .Y(n_1562) );
INVx1_ASAP7_75t_L g1350 ( .A(n_254), .Y(n_1350) );
AO22x1_ASAP7_75t_L g736 ( .A1(n_255), .A2(n_264), .B1(n_722), .B2(n_737), .Y(n_736) );
CKINVDCx5p33_ASAP7_75t_R g1381 ( .A(n_256), .Y(n_1381) );
AOI21xp5_ASAP7_75t_L g1129 ( .A1(n_257), .A2(n_682), .B(n_1130), .Y(n_1129) );
INVx1_ASAP7_75t_L g1160 ( .A(n_257), .Y(n_1160) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_258), .Y(n_573) );
INVxp33_ASAP7_75t_L g986 ( .A(n_259), .Y(n_986) );
INVx2_ASAP7_75t_L g374 ( .A(n_260), .Y(n_374) );
AO22x1_ASAP7_75t_L g738 ( .A1(n_261), .A2(n_268), .B1(n_739), .B2(n_742), .Y(n_738) );
XNOR2x1_ASAP7_75t_L g1222 ( .A(n_262), .B(n_1223), .Y(n_1222) );
CKINVDCx5p33_ASAP7_75t_R g1583 ( .A(n_263), .Y(n_1583) );
INVxp33_ASAP7_75t_SL g547 ( .A(n_265), .Y(n_547) );
INVxp67_ASAP7_75t_L g511 ( .A(n_266), .Y(n_511) );
INVx1_ASAP7_75t_L g549 ( .A(n_267), .Y(n_549) );
AOI222xp33_ASAP7_75t_L g933 ( .A1(n_268), .A2(n_934), .B1(n_1030), .B2(n_1039), .C1(n_1043), .C2(n_1107), .Y(n_933) );
XOR2xp5_ASAP7_75t_L g935 ( .A(n_268), .B(n_936), .Y(n_935) );
INVxp33_ASAP7_75t_SL g437 ( .A(n_269), .Y(n_437) );
INVx1_ASAP7_75t_L g945 ( .A(n_270), .Y(n_945) );
INVx1_ASAP7_75t_L g1195 ( .A(n_271), .Y(n_1195) );
BUFx3_ASAP7_75t_L g299 ( .A(n_272), .Y(n_299) );
INVx1_ASAP7_75t_L g320 ( .A(n_272), .Y(n_320) );
BUFx3_ASAP7_75t_L g300 ( .A(n_273), .Y(n_300) );
INVx1_ASAP7_75t_L g316 ( .A(n_273), .Y(n_316) );
INVxp33_ASAP7_75t_SL g1544 ( .A(n_274), .Y(n_1544) );
CKINVDCx5p33_ASAP7_75t_R g1128 ( .A(n_275), .Y(n_1128) );
INVx1_ASAP7_75t_L g1144 ( .A(n_276), .Y(n_1144) );
INVx1_ASAP7_75t_L g1059 ( .A(n_278), .Y(n_1059) );
INVxp33_ASAP7_75t_L g396 ( .A(n_280), .Y(n_396) );
OAI21xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_1111), .B(n_1635), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_705), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g1636 ( .A(n_283), .B(n_706), .Y(n_1636) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_536), .B1(n_537), .B2(n_704), .Y(n_283) );
INVx1_ASAP7_75t_L g704 ( .A(n_284), .Y(n_704) );
AO22x1_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_466), .B1(n_467), .B2(n_535), .Y(n_284) );
BUFx2_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g535 ( .A(n_286), .Y(n_535) );
XOR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_465), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_382), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_293), .B1(n_368), .B2(n_369), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g1377 ( .A1(n_289), .A2(n_1378), .B1(n_1396), .B2(n_1397), .Y(n_1377) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx8_ASAP7_75t_SL g507 ( .A(n_290), .Y(n_507) );
OAI31xp33_ASAP7_75t_L g1591 ( .A1(n_290), .A2(n_1592), .A3(n_1610), .B(n_1628), .Y(n_1591) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x4_ASAP7_75t_L g969 ( .A(n_291), .B(n_970), .Y(n_969) );
BUFx2_ASAP7_75t_L g1120 ( .A(n_291), .Y(n_1120) );
BUFx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x6_ASAP7_75t_L g429 ( .A(n_292), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g619 ( .A(n_292), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g293 ( .A(n_294), .B(n_338), .C(n_357), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_312), .B1(n_321), .B2(n_325), .C(n_326), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g1318 ( .A1(n_296), .A2(n_322), .B(n_1319), .C(n_1320), .Y(n_1318) );
BUFx4f_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g352 ( .A(n_297), .B(n_322), .Y(n_352) );
BUFx3_ASAP7_75t_L g496 ( .A(n_297), .Y(n_496) );
INVx2_ASAP7_75t_SL g1022 ( .A(n_297), .Y(n_1022) );
AND2x4_ASAP7_75t_L g1235 ( .A(n_297), .B(n_604), .Y(n_1235) );
BUFx6f_ASAP7_75t_L g1571 ( .A(n_297), .Y(n_1571) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_298), .Y(n_343) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx2_ASAP7_75t_L g305 ( .A(n_299), .Y(n_305) );
AND2x4_ASAP7_75t_L g315 ( .A(n_299), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g306 ( .A(n_300), .Y(n_306) );
AND2x4_ASAP7_75t_L g319 ( .A(n_300), .B(n_320), .Y(n_319) );
INVx4_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g1024 ( .A(n_302), .Y(n_1024) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g500 ( .A(n_303), .Y(n_500) );
INVx1_ASAP7_75t_L g583 ( .A(n_303), .Y(n_583) );
INVx2_ASAP7_75t_L g1130 ( .A(n_303), .Y(n_1130) );
INVx2_ASAP7_75t_SL g1208 ( .A(n_303), .Y(n_1208) );
HB1xp67_ASAP7_75t_L g1234 ( .A(n_303), .Y(n_1234) );
INVx1_ASAP7_75t_L g1574 ( .A(n_303), .Y(n_1574) );
INVx6_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g349 ( .A(n_304), .Y(n_349) );
AND2x2_ASAP7_75t_L g381 ( .A(n_304), .B(n_329), .Y(n_381) );
BUFx2_ASAP7_75t_L g601 ( .A(n_304), .Y(n_601) );
AND2x4_ASAP7_75t_L g958 ( .A(n_304), .B(n_959), .Y(n_958) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g337 ( .A(n_305), .Y(n_337) );
INVx1_ASAP7_75t_L g333 ( .A(n_306), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_SL g489 ( .A(n_308), .Y(n_489) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_308), .Y(n_598) );
INVx2_ASAP7_75t_L g682 ( .A(n_308), .Y(n_682) );
AND2x4_ASAP7_75t_L g1029 ( .A(n_308), .B(n_380), .Y(n_1029) );
INVx1_ASAP7_75t_L g1211 ( .A(n_308), .Y(n_1211) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
AND2x4_ASAP7_75t_L g329 ( .A(n_309), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g346 ( .A(n_310), .B(n_311), .Y(n_346) );
INVx1_ASAP7_75t_L g947 ( .A(n_310), .Y(n_947) );
INVx1_ASAP7_75t_L g952 ( .A(n_310), .Y(n_952) );
HB1xp67_ASAP7_75t_L g960 ( .A(n_310), .Y(n_960) );
INVx1_ASAP7_75t_L g970 ( .A(n_311), .Y(n_970) );
BUFx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g321 ( .A(n_314), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g1459 ( .A(n_314), .Y(n_1459) );
INVx2_ASAP7_75t_SL g1577 ( .A(n_314), .Y(n_1577) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_315), .Y(n_480) );
BUFx2_ASAP7_75t_L g495 ( .A(n_315), .Y(n_495) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_315), .Y(n_594) );
INVx2_ASAP7_75t_SL g689 ( .A(n_315), .Y(n_689) );
AND2x6_ASAP7_75t_L g968 ( .A(n_315), .B(n_955), .Y(n_968) );
BUFx6f_ASAP7_75t_L g1202 ( .A(n_315), .Y(n_1202) );
HB1xp67_ASAP7_75t_L g1231 ( .A(n_315), .Y(n_1231) );
BUFx2_ASAP7_75t_L g1242 ( .A(n_315), .Y(n_1242) );
BUFx3_ASAP7_75t_L g1310 ( .A(n_315), .Y(n_1310) );
INVx1_ASAP7_75t_L g363 ( .A(n_316), .Y(n_363) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g1051 ( .A(n_318), .Y(n_1051) );
BUFx3_ASAP7_75t_L g1388 ( .A(n_318), .Y(n_1388) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g351 ( .A(n_319), .Y(n_351) );
INVx2_ASAP7_75t_L g367 ( .A(n_319), .Y(n_367) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_319), .Y(n_503) );
INVx1_ASAP7_75t_L g1527 ( .A(n_319), .Y(n_1527) );
INVx1_ASAP7_75t_L g362 ( .A(n_320), .Y(n_362) );
AOI211xp5_ASAP7_75t_L g473 ( .A1(n_321), .A2(n_474), .B(n_475), .C(n_477), .Y(n_473) );
AOI211xp5_ASAP7_75t_L g672 ( .A1(n_321), .A2(n_673), .B(n_674), .C(n_678), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_321), .A2(n_359), .B1(n_1059), .B2(n_1060), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_321), .A2(n_359), .B1(n_1139), .B2(n_1140), .Y(n_1138) );
AOI211xp5_ASAP7_75t_L g1455 ( .A1(n_321), .A2(n_1448), .B(n_1456), .C(n_1457), .Y(n_1455) );
AOI211xp5_ASAP7_75t_L g1517 ( .A1(n_321), .A2(n_1499), .B(n_1518), .C(n_1522), .Y(n_1517) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_322), .A2(n_609), .B(n_614), .Y(n_608) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_322), .B(n_1202), .Y(n_1201) );
AOI221xp5_ASAP7_75t_L g1236 ( .A1(n_322), .A2(n_359), .B1(n_1237), .B2(n_1238), .C(n_1245), .Y(n_1236) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g360 ( .A(n_323), .B(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g366 ( .A(n_323), .B(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g1543 ( .A(n_323), .B(n_393), .Y(n_1543) );
INVx1_ASAP7_75t_L g330 ( .A(n_324), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_325), .A2(n_364), .B1(n_444), .B2(n_453), .Y(n_452) );
INVx2_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g476 ( .A(n_328), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_328), .A2(n_335), .B1(n_606), .B2(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g675 ( .A(n_328), .Y(n_675) );
AOI222xp33_ASAP7_75t_L g1063 ( .A1(n_328), .A2(n_677), .B1(n_1064), .B2(n_1065), .C1(n_1067), .C2(n_1068), .Y(n_1063) );
INVx2_ASAP7_75t_SL g1519 ( .A(n_328), .Y(n_1519) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
AND2x2_ASAP7_75t_L g335 ( .A(n_329), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g356 ( .A(n_329), .Y(n_356) );
BUFx2_ASAP7_75t_L g604 ( .A(n_329), .Y(n_604) );
AND2x2_ASAP7_75t_L g677 ( .A(n_329), .B(n_336), .Y(n_677) );
AND2x4_ASAP7_75t_L g1215 ( .A(n_329), .B(n_331), .Y(n_1215) );
AND2x4_ASAP7_75t_L g1217 ( .A(n_329), .B(n_336), .Y(n_1217) );
NAND2x1p5_ASAP7_75t_L g1561 ( .A(n_329), .B(n_461), .Y(n_1561) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g1559 ( .A(n_332), .Y(n_1559) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g949 ( .A(n_333), .Y(n_949) );
INVx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g1521 ( .A(n_336), .Y(n_1521) );
BUFx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x6_ASAP7_75t_L g951 ( .A(n_337), .B(n_952), .Y(n_951) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_347), .B1(n_352), .B2(n_353), .C(n_354), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g1136 ( .A(n_341), .Y(n_1136) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g354 ( .A(n_342), .B(n_355), .Y(n_354) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_342), .Y(n_602) );
INVx1_ASAP7_75t_L g1510 ( .A(n_342), .Y(n_1510) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g693 ( .A(n_343), .Y(n_693) );
AND2x4_ASAP7_75t_L g953 ( .A(n_343), .B(n_954), .Y(n_953) );
BUFx6f_ASAP7_75t_L g1369 ( .A(n_343), .Y(n_1369) );
INVx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g1054 ( .A(n_345), .Y(n_1054) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_SL g590 ( .A(n_346), .Y(n_590) );
INVx2_ASAP7_75t_L g1018 ( .A(n_346), .Y(n_1018) );
INVx1_ASAP7_75t_L g1370 ( .A(n_346), .Y(n_1370) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_SL g696 ( .A(n_349), .Y(n_696) );
INVx1_ASAP7_75t_L g1385 ( .A(n_349), .Y(n_1385) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g1025 ( .A(n_351), .Y(n_1025) );
INVx1_ASAP7_75t_L g492 ( .A(n_352), .Y(n_492) );
INVx1_ASAP7_75t_L g685 ( .A(n_352), .Y(n_685) );
INVx1_ASAP7_75t_L g1062 ( .A(n_352), .Y(n_1062) );
INVx2_ASAP7_75t_SL g1133 ( .A(n_352), .Y(n_1133) );
AOI221xp5_ASAP7_75t_L g1367 ( .A1(n_352), .A2(n_1235), .B1(n_1357), .B2(n_1368), .C(n_1371), .Y(n_1367) );
BUFx6f_ASAP7_75t_L g1516 ( .A(n_352), .Y(n_1516) );
OAI22xp33_ASAP7_75t_L g455 ( .A1(n_353), .A2(n_358), .B1(n_435), .B2(n_456), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g490 ( .A1(n_354), .A2(n_491), .B1(n_493), .B2(n_494), .C(n_497), .Y(n_490) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_354), .A2(n_684), .B1(n_686), .B2(n_687), .C(n_694), .Y(n_683) );
INVx1_ASAP7_75t_L g1069 ( .A(n_354), .Y(n_1069) );
AOI221xp5_ASAP7_75t_L g1131 ( .A1(n_354), .A2(n_1132), .B1(n_1134), .B2(n_1135), .C(n_1137), .Y(n_1131) );
AOI221xp5_ASAP7_75t_L g1203 ( .A1(n_354), .A2(n_1132), .B1(n_1195), .B2(n_1204), .C(n_1205), .Y(n_1203) );
AOI221xp5_ASAP7_75t_L g1462 ( .A1(n_354), .A2(n_684), .B1(n_1451), .B2(n_1463), .C(n_1464), .Y(n_1462) );
AOI221xp5_ASAP7_75t_L g1507 ( .A1(n_354), .A2(n_1503), .B1(n_1508), .B2(n_1513), .C(n_1516), .Y(n_1507) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g1520 ( .A(n_356), .B(n_1521), .Y(n_1520) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B1(n_364), .B2(n_365), .Y(n_357) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_359), .A2(n_365), .B1(n_505), .B2(n_506), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_359), .A2(n_365), .B1(n_701), .B2(n_702), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g1198 ( .A1(n_359), .A2(n_1191), .B1(n_1194), .B2(n_1199), .Y(n_1198) );
AOI22xp5_ASAP7_75t_L g1372 ( .A1(n_359), .A2(n_365), .B1(n_1350), .B2(n_1356), .Y(n_1372) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_359), .A2(n_1201), .B1(n_1380), .B2(n_1381), .Y(n_1379) );
AOI22xp33_ASAP7_75t_L g1468 ( .A1(n_359), .A2(n_365), .B1(n_1447), .B2(n_1450), .Y(n_1468) );
AOI22xp33_ASAP7_75t_SL g1532 ( .A1(n_359), .A2(n_365), .B1(n_1500), .B2(n_1502), .Y(n_1532) );
INVx6_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g486 ( .A(n_361), .Y(n_486) );
INVx2_ASAP7_75t_L g611 ( .A(n_361), .Y(n_611) );
OR2x2_ASAP7_75t_L g965 ( .A(n_361), .B(n_966), .Y(n_965) );
OR2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
AND2x2_ASAP7_75t_L g483 ( .A(n_362), .B(n_363), .Y(n_483) );
AOI211xp5_ASAP7_75t_L g1122 ( .A1(n_365), .A2(n_1123), .B(n_1124), .C(n_1125), .Y(n_1122) );
AOI221xp5_ASAP7_75t_L g1209 ( .A1(n_365), .A2(n_1192), .B1(n_1210), .B2(n_1212), .C(n_1213), .Y(n_1209) );
AOI221xp5_ASAP7_75t_L g1382 ( .A1(n_365), .A2(n_1383), .B1(n_1384), .B2(n_1387), .C(n_1389), .Y(n_1382) );
INVx4_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g613 ( .A(n_367), .Y(n_613) );
INVx2_ASAP7_75t_L g699 ( .A(n_367), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g470 ( .A1(n_369), .A2(n_471), .B(n_472), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g1119 ( .A1(n_369), .A2(n_1120), .B1(n_1121), .B2(n_1141), .Y(n_1119) );
INVx5_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g669 ( .A(n_370), .Y(n_669) );
INVx1_ASAP7_75t_L g1219 ( .A(n_370), .Y(n_1219) );
INVx2_ASAP7_75t_SL g1373 ( .A(n_370), .Y(n_1373) );
INVx2_ASAP7_75t_L g1397 ( .A(n_370), .Y(n_1397) );
AND2x4_ASAP7_75t_L g370 ( .A(n_371), .B(n_378), .Y(n_370) );
INVx2_ASAP7_75t_L g550 ( .A(n_371), .Y(n_550) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_376), .Y(n_371) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_372), .Y(n_436) );
INVx2_ASAP7_75t_SL g524 ( .A(n_372), .Y(n_524) );
OR2x6_ASAP7_75t_L g974 ( .A(n_372), .B(n_975), .Y(n_974) );
OR2x6_ASAP7_75t_L g976 ( .A(n_372), .B(n_977), .Y(n_976) );
BUFx2_ASAP7_75t_L g1084 ( .A(n_372), .Y(n_1084) );
INVx1_ASAP7_75t_L g1101 ( .A(n_372), .Y(n_1101) );
OAI22xp33_ASAP7_75t_L g1273 ( .A1(n_372), .A2(n_1087), .B1(n_1237), .B2(n_1274), .Y(n_1273) );
INVx2_ASAP7_75t_SL g1355 ( .A(n_372), .Y(n_1355) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
AND2x4_ASAP7_75t_L g390 ( .A(n_374), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g400 ( .A(n_374), .Y(n_400) );
AND2x2_ASAP7_75t_L g406 ( .A(n_374), .B(n_375), .Y(n_406) );
INVx2_ASAP7_75t_L g411 ( .A(n_374), .Y(n_411) );
INVx1_ASAP7_75t_L g441 ( .A(n_374), .Y(n_441) );
INVx2_ASAP7_75t_L g391 ( .A(n_375), .Y(n_391) );
INVx1_ASAP7_75t_L g413 ( .A(n_375), .Y(n_413) );
INVx1_ASAP7_75t_L g420 ( .A(n_375), .Y(n_420) );
INVx1_ASAP7_75t_L g440 ( .A(n_375), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_375), .B(n_411), .Y(n_448) );
INVx3_ASAP7_75t_L g421 ( .A(n_376), .Y(n_421) );
INVx1_ASAP7_75t_L g1590 ( .A(n_377), .Y(n_1590) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OR2x6_ASAP7_75t_L g1584 ( .A(n_379), .B(n_1585), .Y(n_1584) );
AND2x4_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
OR2x2_ASAP7_75t_L g992 ( .A(n_380), .B(n_993), .Y(n_992) );
INVx2_ASAP7_75t_L g1066 ( .A(n_381), .Y(n_1066) );
NOR3xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_414), .C(n_428), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_401), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B1(n_396), .B2(n_397), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g1094 ( .A1(n_386), .A2(n_667), .B1(n_1095), .B2(n_1104), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_386), .A2(n_397), .B1(n_1128), .B2(n_1158), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g1168 ( .A1(n_386), .A2(n_397), .B1(n_1169), .B2(n_1170), .Y(n_1168) );
BUFx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx2_ASAP7_75t_L g531 ( .A(n_387), .Y(n_531) );
BUFx2_ASAP7_75t_L g544 ( .A(n_387), .Y(n_544) );
BUFx2_ASAP7_75t_L g642 ( .A(n_387), .Y(n_642) );
BUFx2_ASAP7_75t_L g1257 ( .A(n_387), .Y(n_1257) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_392), .Y(n_387) );
BUFx3_ASAP7_75t_L g454 ( .A(n_388), .Y(n_454) );
INVx1_ASAP7_75t_L g521 ( .A(n_388), .Y(n_521) );
INVx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_389), .Y(n_561) );
INVx3_ASAP7_75t_L g1154 ( .A(n_389), .Y(n_1154) );
INVx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_390), .Y(n_451) );
INVx1_ASAP7_75t_L g991 ( .A(n_390), .Y(n_991) );
INVx1_ASAP7_75t_L g1007 ( .A(n_390), .Y(n_1007) );
AND2x4_ASAP7_75t_L g399 ( .A(n_391), .B(n_400), .Y(n_399) );
AND2x6_ASAP7_75t_L g397 ( .A(n_392), .B(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g403 ( .A(n_392), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g408 ( .A(n_392), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g534 ( .A(n_392), .B(n_409), .Y(n_534) );
AND2x2_ASAP7_75t_L g548 ( .A(n_392), .B(n_409), .Y(n_548) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_392), .B(n_1261), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_392), .B(n_409), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_392), .B(n_1154), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_392), .B(n_666), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_392), .B(n_409), .Y(n_1406) );
AND2x4_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g461 ( .A(n_393), .Y(n_461) );
INVx2_ASAP7_75t_L g1596 ( .A(n_394), .Y(n_1596) );
AND2x4_ASAP7_75t_L g1612 ( .A(n_394), .B(n_566), .Y(n_1612) );
AND2x2_ASAP7_75t_L g1630 ( .A(n_394), .B(n_410), .Y(n_1630) );
INVx1_ASAP7_75t_L g432 ( .A(n_395), .Y(n_432) );
INVx1_ASAP7_75t_L g463 ( .A(n_395), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_397), .A2(n_484), .B1(n_530), .B2(n_531), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_397), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_397), .A2(n_641), .B1(n_642), .B2(n_643), .Y(n_640) );
INVx1_ASAP7_75t_SL g1073 ( .A(n_397), .Y(n_1073) );
AOI22xp5_ASAP7_75t_L g1252 ( .A1(n_397), .A2(n_534), .B1(n_1253), .B2(n_1254), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g1293 ( .A1(n_397), .A2(n_1294), .B1(n_1295), .B2(n_1296), .Y(n_1293) );
AOI22xp33_ASAP7_75t_L g1400 ( .A1(n_397), .A2(n_531), .B1(n_1401), .B2(n_1402), .Y(n_1400) );
AOI22xp33_ASAP7_75t_L g1427 ( .A1(n_397), .A2(n_1257), .B1(n_1428), .B2(n_1429), .Y(n_1427) );
AOI22xp33_ASAP7_75t_L g1479 ( .A1(n_397), .A2(n_544), .B1(n_1480), .B2(n_1481), .Y(n_1479) );
NAND2x1p5_ASAP7_75t_L g427 ( .A(n_398), .B(n_421), .Y(n_427) );
BUFx2_ASAP7_75t_L g1080 ( .A(n_398), .Y(n_1080) );
BUFx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_399), .Y(n_569) );
BUFx3_ASAP7_75t_L g577 ( .A(n_399), .Y(n_577) );
BUFx2_ASAP7_75t_L g631 ( .A(n_399), .Y(n_631) );
INVx1_ASAP7_75t_L g656 ( .A(n_399), .Y(n_656) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_399), .Y(n_666) );
AND2x4_ASAP7_75t_L g982 ( .A(n_399), .B(n_983), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_407), .B2(n_408), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_403), .A2(n_487), .B1(n_533), .B2(n_534), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_403), .A2(n_552), .B(n_553), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_403), .A2(n_408), .B1(n_645), .B2(n_646), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_403), .A2(n_408), .B1(n_1092), .B2(n_1093), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_403), .A2(n_534), .B1(n_1160), .B2(n_1161), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_403), .A2(n_534), .B1(n_1172), .B2(n_1173), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_403), .B(n_1291), .Y(n_1290) );
AOI22xp33_ASAP7_75t_L g1403 ( .A1(n_403), .A2(n_1404), .B1(n_1405), .B2(n_1406), .Y(n_1403) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_403), .A2(n_548), .B1(n_1431), .B2(n_1432), .Y(n_1430) );
AOI22xp33_ASAP7_75t_L g1482 ( .A1(n_403), .A2(n_1406), .B1(n_1483), .B2(n_1484), .Y(n_1482) );
INVx1_ASAP7_75t_L g998 ( .A(n_404), .Y(n_998) );
INVx2_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g1009 ( .A(n_405), .Y(n_1009) );
INVx2_ASAP7_75t_SL g1261 ( .A(n_405), .Y(n_1261) );
INVx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_406), .Y(n_566) );
INVx2_ASAP7_75t_SL g1097 ( .A(n_409), .Y(n_1097) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_410), .Y(n_659) );
AND2x4_ASAP7_75t_L g987 ( .A(n_410), .B(n_977), .Y(n_987) );
INVx1_ASAP7_75t_L g1003 ( .A(n_410), .Y(n_1003) );
INVx1_ASAP7_75t_L g1011 ( .A(n_410), .Y(n_1011) );
BUFx2_ASAP7_75t_L g1076 ( .A(n_410), .Y(n_1076) );
BUFx6f_ASAP7_75t_L g1285 ( .A(n_410), .Y(n_1285) );
AND2x4_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx1_ASAP7_75t_L g425 ( .A(n_411), .Y(n_425) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g1336 ( .A(n_416), .Y(n_1336) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
HB1xp67_ASAP7_75t_L g1408 ( .A(n_417), .Y(n_1408) );
NAND2x1_ASAP7_75t_SL g417 ( .A(n_418), .B(n_421), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_418), .A2(n_424), .B1(n_1067), .B2(n_1068), .Y(n_1089) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_420), .Y(n_629) );
AND2x4_ASAP7_75t_L g980 ( .A(n_420), .B(n_975), .Y(n_980) );
NAND2x1p5_ASAP7_75t_L g423 ( .A(n_421), .B(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g623 ( .A(n_421), .B(n_624), .Y(n_623) );
AND2x4_ASAP7_75t_L g628 ( .A(n_421), .B(n_629), .Y(n_628) );
AND2x4_ASAP7_75t_L g630 ( .A(n_421), .B(n_631), .Y(n_630) );
AOI32xp33_ASAP7_75t_L g1074 ( .A1(n_421), .A2(n_649), .A3(n_1075), .B1(n_1079), .B2(n_1081), .Y(n_1074) );
BUFx4f_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx4f_ASAP7_75t_L g527 ( .A(n_423), .Y(n_527) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OR2x6_ASAP7_75t_L g1609 ( .A(n_425), .B(n_1589), .Y(n_1609) );
BUFx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g1175 ( .A(n_427), .Y(n_1175) );
BUFx2_ASAP7_75t_L g1434 ( .A(n_427), .Y(n_1434) );
OAI33xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_433), .A3(n_442), .B1(n_452), .B2(n_455), .B3(n_458), .Y(n_428) );
OAI33xp33_ASAP7_75t_L g509 ( .A1(n_429), .A2(n_458), .A3(n_510), .B1(n_514), .B2(n_520), .B3(n_522), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_429), .A2(n_458), .B1(n_554), .B2(n_570), .Y(n_553) );
HB1xp67_ASAP7_75t_L g1177 ( .A(n_429), .Y(n_1177) );
OAI33xp33_ASAP7_75t_L g1337 ( .A1(n_429), .A2(n_1338), .A3(n_1341), .B1(n_1347), .B2(n_1353), .B3(n_1358), .Y(n_1337) );
OAI33xp33_ASAP7_75t_L g1409 ( .A1(n_429), .A2(n_458), .A3(n_1410), .B1(n_1414), .B2(n_1419), .B3(n_1420), .Y(n_1409) );
OAI33xp33_ASAP7_75t_L g1435 ( .A1(n_429), .A2(n_458), .A3(n_1436), .B1(n_1440), .B2(n_1446), .B3(n_1449), .Y(n_1435) );
OAI33xp33_ASAP7_75t_L g1486 ( .A1(n_429), .A2(n_458), .A3(n_1487), .B1(n_1493), .B2(n_1497), .B3(n_1501), .Y(n_1486) );
OR2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g651 ( .A(n_431), .Y(n_651) );
INVx1_ASAP7_75t_L g977 ( .A(n_432), .Y(n_977) );
OAI22xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B1(n_437), .B2(n_438), .Y(n_433) );
OAI22xp33_ASAP7_75t_L g514 ( .A1(n_435), .A2(n_515), .B1(n_516), .B2(n_517), .Y(n_514) );
BUFx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g1180 ( .A(n_436), .Y(n_1180) );
OAI22xp33_ASAP7_75t_L g1446 ( .A1(n_436), .A2(n_1190), .B1(n_1447), .B2(n_1448), .Y(n_1446) );
OAI22xp33_ASAP7_75t_L g1338 ( .A1(n_438), .A2(n_1082), .B1(n_1339), .B2(n_1340), .Y(n_1338) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx2_ASAP7_75t_L g457 ( .A(n_439), .Y(n_457) );
INVx3_ASAP7_75t_L g519 ( .A(n_439), .Y(n_519) );
INVx2_ASAP7_75t_L g1627 ( .A(n_439), .Y(n_1627) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_440), .B(n_441), .Y(n_1088) );
INVx1_ASAP7_75t_L g625 ( .A(n_441), .Y(n_625) );
OAI22xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_444), .B1(n_449), .B2(n_450), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_444), .A2(n_474), .B1(n_506), .B2(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g512 ( .A(n_445), .Y(n_512) );
INVx2_ASAP7_75t_L g1416 ( .A(n_445), .Y(n_1416) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g1190 ( .A(n_446), .Y(n_1190) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g572 ( .A(n_447), .Y(n_572) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g557 ( .A(n_448), .Y(n_557) );
INVx1_ASAP7_75t_L g1186 ( .A(n_448), .Y(n_1186) );
OAI221xp5_ASAP7_75t_L g570 ( .A1(n_450), .A2(n_571), .B1(n_573), .B2(n_574), .C(n_575), .Y(n_570) );
OAI221xp5_ASAP7_75t_L g1597 ( .A1(n_450), .A2(n_1540), .B1(n_1551), .B2(n_1598), .C(n_1601), .Y(n_1597) );
INVx2_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_SL g661 ( .A(n_451), .Y(n_661) );
BUFx3_ASAP7_75t_L g663 ( .A(n_451), .Y(n_663) );
INVx4_ASAP7_75t_L g1078 ( .A(n_451), .Y(n_1078) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_453), .A2(n_511), .B1(n_512), .B2(n_513), .Y(n_510) );
OAI22xp33_ASAP7_75t_L g1449 ( .A1(n_453), .A2(n_1438), .B1(n_1450), .B2(n_1451), .Y(n_1449) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_454), .Y(n_453) );
OAI22xp33_ASAP7_75t_L g1410 ( .A1(n_456), .A2(n_1411), .B1(n_1412), .B2(n_1413), .Y(n_1410) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OAI33xp33_ASAP7_75t_L g1176 ( .A1(n_458), .A2(n_1177), .A3(n_1178), .B1(n_1183), .B2(n_1189), .B3(n_1193), .Y(n_1176) );
CKINVDCx8_ASAP7_75t_R g458 ( .A(n_459), .Y(n_458) );
INVx5_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx6_ASAP7_75t_L g667 ( .A(n_460), .Y(n_667) );
OR2x6_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx2_ASAP7_75t_L g1289 ( .A(n_462), .Y(n_1289) );
NAND2x1p5_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
INVx1_ASAP7_75t_L g984 ( .A(n_463), .Y(n_984) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_508), .Y(n_469) );
AOI31xp33_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_490), .A3(n_504), .B(n_507), .Y(n_472) );
INVx2_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_SL g588 ( .A(n_480), .Y(n_588) );
OAI221xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_484), .B1(n_485), .B2(n_487), .C(n_488), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_L g586 ( .A(n_483), .Y(n_586) );
BUFx4f_ASAP7_75t_L g597 ( .A(n_483), .Y(n_597) );
INVx1_ASAP7_75t_L g943 ( .A(n_483), .Y(n_943) );
INVx1_ASAP7_75t_L g1240 ( .A(n_483), .Y(n_1240) );
INVx2_ASAP7_75t_L g1313 ( .A(n_483), .Y(n_1313) );
OAI221xp5_ASAP7_75t_L g595 ( .A1(n_485), .A2(n_545), .B1(n_552), .B2(n_596), .C(n_598), .Y(n_595) );
OAI221xp5_ASAP7_75t_L g679 ( .A1(n_485), .A2(n_643), .B1(n_645), .B2(n_680), .C(n_681), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g1460 ( .A1(n_485), .A2(n_681), .B1(n_1429), .B2(n_1431), .C(n_1461), .Y(n_1460) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g1531 ( .A(n_489), .Y(n_1531) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
OAI22xp33_ASAP7_75t_L g522 ( .A1(n_493), .A2(n_505), .B1(n_523), .B2(n_525), .Y(n_522) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx6f_ASAP7_75t_L g1228 ( .A(n_500), .Y(n_1228) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_503), .Y(n_580) );
AND2x6_ASAP7_75t_L g962 ( .A(n_503), .B(n_963), .Y(n_962) );
BUFx6f_ASAP7_75t_L g1244 ( .A(n_503), .Y(n_1244) );
INVx1_ASAP7_75t_L g1467 ( .A(n_503), .Y(n_1467) );
INVx5_ASAP7_75t_L g1070 ( .A(n_507), .Y(n_1070) );
NOR3xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_526), .C(n_528), .Y(n_508) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g1438 ( .A(n_518), .Y(n_1438) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx2_ASAP7_75t_L g525 ( .A(n_519), .Y(n_525) );
OAI22xp33_ASAP7_75t_L g1436 ( .A1(n_523), .A2(n_1437), .B1(n_1438), .B2(n_1439), .Y(n_1436) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OAI22xp33_ASAP7_75t_L g1178 ( .A1(n_525), .A2(n_1179), .B1(n_1181), .B2(n_1182), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_532), .Y(n_528) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AO22x2_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_632), .B1(n_633), .B2(n_703), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g703 ( .A(n_539), .Y(n_703) );
NAND4xp25_ASAP7_75t_L g540 ( .A(n_541), .B(n_551), .C(n_578), .D(n_620), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .Y(n_541) );
AOI22xp33_ASAP7_75t_SL g546 ( .A1(n_547), .A2(n_548), .B1(n_549), .B2(n_550), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g600 ( .A1(n_549), .A2(n_601), .B(n_602), .C(n_603), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g1255 ( .A1(n_550), .A2(n_1256), .B1(n_1257), .B2(n_1258), .Y(n_1255) );
AOI22xp33_ASAP7_75t_L g1297 ( .A1(n_550), .A2(n_1298), .B1(n_1299), .B2(n_1300), .Y(n_1297) );
OAI221xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_558), .B1(n_559), .B2(n_562), .C(n_563), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g1440 ( .A1(n_555), .A2(n_1441), .B1(n_1442), .B2(n_1445), .Y(n_1440) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx2_ASAP7_75t_L g1498 ( .A(n_557), .Y(n_1498) );
OAI221xp5_ASAP7_75t_L g584 ( .A1(n_558), .A2(n_585), .B1(n_587), .B2(n_588), .C(n_589), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g1497 ( .A1(n_559), .A2(n_1498), .B1(n_1499), .B2(n_1500), .Y(n_1497) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g1013 ( .A(n_561), .Y(n_1013) );
INVx2_ASAP7_75t_L g1098 ( .A(n_561), .Y(n_1098) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g1283 ( .A(n_565), .Y(n_1283) );
INVx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
BUFx2_ASAP7_75t_L g654 ( .A(n_566), .Y(n_654) );
BUFx6f_ASAP7_75t_L g1148 ( .A(n_566), .Y(n_1148) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g1149 ( .A(n_568), .Y(n_1149) );
INVx2_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
BUFx2_ASAP7_75t_L g1014 ( .A(n_569), .Y(n_1014) );
BUFx2_ASAP7_75t_L g1615 ( .A(n_571), .Y(n_1615) );
INVx2_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g1349 ( .A(n_572), .Y(n_1349) );
INVx2_ASAP7_75t_L g1495 ( .A(n_572), .Y(n_1495) );
INVx2_ASAP7_75t_L g1600 ( .A(n_572), .Y(n_1600) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g1000 ( .A(n_577), .Y(n_1000) );
AND2x4_ASAP7_75t_L g1594 ( .A(n_577), .B(n_1595), .Y(n_1594) );
OAI31xp33_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_591), .A3(n_599), .B(n_617), .Y(n_578) );
HB1xp67_ASAP7_75t_L g1515 ( .A(n_580), .Y(n_1515) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
HB1xp67_ASAP7_75t_L g1465 ( .A(n_583), .Y(n_1465) );
OAI21xp5_ASAP7_75t_SL g1127 ( .A1(n_585), .A2(n_1128), .B(n_1129), .Y(n_1127) );
INVx2_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g1461 ( .A(n_586), .Y(n_1461) );
INVx1_ASAP7_75t_L g1529 ( .A(n_586), .Y(n_1529) );
INVx1_ASAP7_75t_L g1053 ( .A(n_588), .Y(n_1053) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g615 ( .A(n_594), .Y(n_615) );
BUFx3_ASAP7_75t_L g1056 ( .A(n_594), .Y(n_1056) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_SL g616 ( .A(n_597), .Y(n_616) );
INVx1_ASAP7_75t_L g680 ( .A(n_597), .Y(n_680) );
INVx1_ASAP7_75t_L g1306 ( .A(n_597), .Y(n_1306) );
NAND3xp33_ASAP7_75t_L g599 ( .A(n_600), .B(n_605), .C(n_608), .Y(n_599) );
BUFx3_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_606), .A2(n_607), .B1(n_621), .B2(n_626), .C(n_630), .Y(n_620) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g1530 ( .A(n_611), .Y(n_1530) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g1020 ( .A(n_615), .Y(n_1020) );
INVx1_ASAP7_75t_L g1126 ( .A(n_615), .Y(n_1126) );
AOI22xp5_ASAP7_75t_L g1359 ( .A1(n_617), .A2(n_1360), .B1(n_1373), .B2(n_1374), .Y(n_1359) );
INVx2_ASAP7_75t_L g1469 ( .A(n_617), .Y(n_1469) );
CKINVDCx8_ASAP7_75t_R g617 ( .A(n_618), .Y(n_617) );
AOI31xp33_ASAP7_75t_L g671 ( .A1(n_618), .A2(n_672), .A3(n_683), .B(n_700), .Y(n_671) );
BUFx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x4_ASAP7_75t_L g649 ( .A(n_619), .B(n_650), .Y(n_649) );
AND2x4_ASAP7_75t_L g995 ( .A(n_619), .B(n_650), .Y(n_995) );
OR2x6_ASAP7_75t_L g1017 ( .A(n_619), .B(n_1018), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_619), .B(n_1289), .Y(n_1288) );
INVx2_ASAP7_75t_L g1586 ( .A(n_619), .Y(n_1586) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_621), .A2(n_628), .B1(n_637), .B2(n_638), .C(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g1143 ( .A1(n_623), .A2(n_628), .B1(n_630), .B2(n_1144), .C(n_1145), .Y(n_1143) );
AOI221xp5_ASAP7_75t_L g1249 ( .A1(n_623), .A2(n_628), .B1(n_630), .B2(n_1250), .C(n_1251), .Y(n_1249) );
AOI221xp5_ASAP7_75t_L g1278 ( .A1(n_623), .A2(n_628), .B1(n_630), .B2(n_1279), .C(n_1280), .Y(n_1278) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g981 ( .A(n_625), .B(n_652), .Y(n_981) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_629), .B(n_1588), .Y(n_1607) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_630), .Y(n_639) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_668), .Y(n_634) );
AND4x1_ASAP7_75t_L g635 ( .A(n_636), .B(n_640), .C(n_644), .D(n_647), .Y(n_635) );
AOI33xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_653), .A3(n_657), .B1(n_662), .B2(n_664), .B3(n_667), .Y(n_647) );
BUFx3_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g1625 ( .A(n_650), .Y(n_1625) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
HB1xp67_ASAP7_75t_L g993 ( .A(n_651), .Y(n_993) );
INVx2_ASAP7_75t_SL g975 ( .A(n_652), .Y(n_975) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
BUFx3_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI33xp33_ASAP7_75t_L g994 ( .A1(n_667), .A2(n_995), .A3(n_996), .B1(n_1001), .B2(n_1008), .B3(n_1012), .Y(n_994) );
AOI33xp33_ASAP7_75t_L g1146 ( .A1(n_667), .A2(n_995), .A3(n_1147), .B1(n_1150), .B2(n_1151), .B3(n_1155), .Y(n_1146) );
AOI222xp33_ASAP7_75t_L g1259 ( .A1(n_667), .A2(n_995), .B1(n_1260), .B2(n_1262), .C1(n_1263), .C2(n_1269), .Y(n_1259) );
INVx1_ASAP7_75t_L g1358 ( .A(n_667), .Y(n_1358) );
AOI21xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B(n_671), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g1452 ( .A1(n_669), .A2(n_1453), .B(n_1454), .Y(n_1452) );
AOI21xp5_ASAP7_75t_L g1504 ( .A1(n_669), .A2(n_1505), .B(n_1506), .Y(n_1504) );
INVx2_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g1392 ( .A(n_689), .Y(n_1392) );
INVx2_ASAP7_75t_L g1553 ( .A(n_689), .Y(n_1553) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
BUFx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_696), .B(n_1550), .Y(n_1549) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
BUFx2_ASAP7_75t_L g1308 ( .A(n_699), .Y(n_1308) );
INVxp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g1637 ( .A(n_706), .B(n_1638), .Y(n_1637) );
OAI21xp5_ASAP7_75t_SL g706 ( .A1(n_707), .A2(n_931), .B(n_933), .Y(n_706) );
AND4x1_ASAP7_75t_L g707 ( .A(n_708), .B(n_844), .C(n_879), .D(n_909), .Y(n_707) );
A2O1A1Ixp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_796), .B(n_797), .C(n_828), .Y(n_708) );
OAI211xp5_ASAP7_75t_SL g709 ( .A1(n_710), .A2(n_744), .B(n_775), .C(n_778), .Y(n_709) );
OR2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_734), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_711), .B(n_793), .Y(n_820) );
AND2x2_ASAP7_75t_L g825 ( .A(n_711), .B(n_735), .Y(n_825) );
AND2x4_ASAP7_75t_SL g920 ( .A(n_711), .B(n_734), .Y(n_920) );
INVx2_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g791 ( .A(n_712), .B(n_734), .Y(n_791) );
INVx2_ASAP7_75t_L g796 ( .A(n_712), .Y(n_796) );
INVx1_ASAP7_75t_L g808 ( .A(n_713), .Y(n_808) );
AND2x4_ASAP7_75t_L g713 ( .A(n_714), .B(n_717), .Y(n_713) );
AND2x2_ASAP7_75t_L g737 ( .A(n_714), .B(n_717), .Y(n_737) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AND2x4_ASAP7_75t_L g722 ( .A(n_715), .B(n_717), .Y(n_722) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_716), .B(n_728), .Y(n_727) );
HB1xp67_ASAP7_75t_L g1034 ( .A(n_718), .Y(n_1034) );
INVx1_ASAP7_75t_L g728 ( .A(n_719), .Y(n_728) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI22xp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_723) );
OAI22xp33_ASAP7_75t_L g756 ( .A1(n_724), .A2(n_732), .B1(n_757), .B2(n_758), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_724), .A2(n_732), .B1(n_762), .B2(n_763), .Y(n_761) );
BUFx3_ASAP7_75t_L g811 ( .A(n_724), .Y(n_811) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
OR2x2_ASAP7_75t_L g732 ( .A(n_726), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g741 ( .A(n_726), .Y(n_741) );
INVx1_ASAP7_75t_L g740 ( .A(n_727), .Y(n_740) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g814 ( .A(n_732), .Y(n_814) );
INVx1_ASAP7_75t_L g743 ( .A(n_733), .Y(n_743) );
AND2x2_ASAP7_75t_L g781 ( .A(n_734), .B(n_770), .Y(n_781) );
AND2x2_ASAP7_75t_L g833 ( .A(n_734), .B(n_794), .Y(n_833) );
OAI221xp5_ASAP7_75t_L g880 ( .A1(n_734), .A2(n_862), .B1(n_881), .B2(n_883), .C(n_885), .Y(n_880) );
AND2x2_ASAP7_75t_L g888 ( .A(n_734), .B(n_846), .Y(n_888) );
CKINVDCx6p67_ASAP7_75t_R g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g803 ( .A(n_735), .B(n_804), .Y(n_803) );
AND2x2_ASAP7_75t_L g817 ( .A(n_735), .B(n_770), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_735), .B(n_850), .Y(n_849) );
AOI221xp5_ASAP7_75t_L g896 ( .A1(n_735), .A2(n_776), .B1(n_897), .B2(n_900), .C(n_902), .Y(n_896) );
A2O1A1Ixp33_ASAP7_75t_L g910 ( .A1(n_735), .A2(n_864), .B(n_911), .C(n_912), .Y(n_910) );
AOI221xp5_ASAP7_75t_L g912 ( .A1(n_735), .A2(n_803), .B1(n_856), .B2(n_913), .C(n_914), .Y(n_912) );
OR2x6_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
AND2x4_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
AND2x4_ASAP7_75t_L g742 ( .A(n_741), .B(n_743), .Y(n_742) );
HB1xp67_ASAP7_75t_L g1109 ( .A(n_743), .Y(n_1109) );
AOI211xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_753), .B(n_764), .C(n_768), .Y(n_744) );
AND2x2_ASAP7_75t_L g822 ( .A(n_745), .B(n_823), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_745), .B(n_766), .Y(n_865) );
AND2x2_ASAP7_75t_L g882 ( .A(n_745), .B(n_754), .Y(n_882) );
AND2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_749), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_746), .B(n_766), .Y(n_765) );
INVx4_ASAP7_75t_L g773 ( .A(n_746), .Y(n_773) );
INVx3_ASAP7_75t_L g786 ( .A(n_746), .Y(n_786) );
NOR2xp67_ASAP7_75t_SL g838 ( .A(n_746), .B(n_839), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g872 ( .A(n_746), .B(n_873), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_746), .B(n_754), .Y(n_894) );
OR2x2_ASAP7_75t_L g922 ( .A(n_746), .B(n_770), .Y(n_922) );
AND2x4_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
AND2x2_ASAP7_75t_L g776 ( .A(n_749), .B(n_777), .Y(n_776) );
OR2x2_ASAP7_75t_L g787 ( .A(n_749), .B(n_788), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_749), .B(n_759), .Y(n_839) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_749), .B(n_759), .Y(n_847) );
OR2x2_ASAP7_75t_L g893 ( .A(n_749), .B(n_894), .Y(n_893) );
BUFx3_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g802 ( .A(n_750), .Y(n_802) );
AND2x2_ASAP7_75t_L g818 ( .A(n_750), .B(n_788), .Y(n_818) );
AND2x2_ASAP7_75t_L g827 ( .A(n_750), .B(n_766), .Y(n_827) );
AND2x2_ASAP7_75t_L g837 ( .A(n_750), .B(n_754), .Y(n_837) );
AND2x2_ASAP7_75t_L g860 ( .A(n_750), .B(n_823), .Y(n_860) );
OR2x2_ASAP7_75t_L g908 ( .A(n_750), .B(n_877), .Y(n_908) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
AOI21xp33_ASAP7_75t_L g841 ( .A1(n_753), .A2(n_842), .B(n_843), .Y(n_841) );
AOI21xp5_ASAP7_75t_L g907 ( .A1(n_753), .A2(n_843), .B(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_754), .B(n_801), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_754), .B(n_786), .Y(n_899) );
AND2x2_ASAP7_75t_L g754 ( .A(n_755), .B(n_759), .Y(n_754) );
INVx1_ASAP7_75t_L g767 ( .A(n_755), .Y(n_767) );
INVx1_ASAP7_75t_L g788 ( .A(n_755), .Y(n_788) );
AND2x2_ASAP7_75t_L g823 ( .A(n_755), .B(n_760), .Y(n_823) );
AND2x2_ASAP7_75t_L g774 ( .A(n_759), .B(n_767), .Y(n_774) );
INVx2_ASAP7_75t_L g782 ( .A(n_759), .Y(n_782) );
AND2x2_ASAP7_75t_L g906 ( .A(n_759), .B(n_802), .Y(n_906) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
AND2x2_ASAP7_75t_L g766 ( .A(n_760), .B(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g777 ( .A(n_766), .B(n_773), .Y(n_777) );
INVx1_ASAP7_75t_L g877 ( .A(n_766), .Y(n_877) );
AND2x2_ASAP7_75t_L g884 ( .A(n_766), .B(n_801), .Y(n_884) );
AND2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_774), .Y(n_768) );
INVx1_ASAP7_75t_L g915 ( .A(n_769), .Y(n_915) );
AND2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_773), .Y(n_769) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_770), .Y(n_794) );
INVx1_ASAP7_75t_SL g804 ( .A(n_770), .Y(n_804) );
INVx1_ASAP7_75t_L g840 ( .A(n_770), .Y(n_840) );
INVx1_ASAP7_75t_L g869 ( .A(n_770), .Y(n_869) );
AND2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_773), .B(n_781), .Y(n_780) );
AND2x2_ASAP7_75t_L g801 ( .A(n_773), .B(n_802), .Y(n_801) );
AND2x2_ASAP7_75t_L g831 ( .A(n_773), .B(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g846 ( .A(n_773), .Y(n_846) );
AND2x2_ASAP7_75t_L g856 ( .A(n_773), .B(n_857), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_773), .B(n_803), .Y(n_878) );
AND2x2_ASAP7_75t_L g917 ( .A(n_773), .B(n_817), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_774), .B(n_802), .Y(n_863) );
INVx1_ASAP7_75t_L g923 ( .A(n_774), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_774), .B(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
AOI221xp5_ASAP7_75t_L g830 ( .A1(n_777), .A2(n_781), .B1(n_831), .B2(n_833), .C(n_834), .Y(n_830) );
A2O1A1Ixp33_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_782), .B(n_783), .C(n_789), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_781), .B(n_822), .Y(n_835) );
A2O1A1Ixp33_ASAP7_75t_L g903 ( .A1(n_781), .A2(n_805), .B(n_904), .C(n_907), .Y(n_903) );
INVxp67_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
OR2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_787), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_785), .B(n_833), .Y(n_843) );
A2O1A1Ixp33_ASAP7_75t_L g924 ( .A1(n_785), .A2(n_925), .B(n_926), .C(n_927), .Y(n_924) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_786), .B(n_854), .Y(n_853) );
OR2x2_ASAP7_75t_L g862 ( .A(n_786), .B(n_863), .Y(n_862) );
AND2x2_ASAP7_75t_L g867 ( .A(n_786), .B(n_847), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_786), .B(n_906), .Y(n_905) );
NOR2x1_ASAP7_75t_L g832 ( .A(n_788), .B(n_802), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_788), .B(n_802), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_792), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_795), .Y(n_792) );
AOI321xp33_ASAP7_75t_L g844 ( .A1(n_793), .A2(n_803), .A3(n_845), .B1(n_848), .B2(n_851), .C(n_861), .Y(n_844) );
OR2x2_ASAP7_75t_L g864 ( .A(n_793), .B(n_865), .Y(n_864) );
NOR2xp33_ASAP7_75t_L g883 ( .A(n_793), .B(n_884), .Y(n_883) );
INVx3_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g881 ( .A(n_794), .B(n_882), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_794), .B(n_920), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_795), .B(n_806), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_795), .B(n_806), .Y(n_829) );
AOI21xp5_ASAP7_75t_SL g909 ( .A1(n_795), .A2(n_910), .B(n_918), .Y(n_909) );
NOR3xp33_ASAP7_75t_L g921 ( .A(n_795), .B(n_922), .C(n_923), .Y(n_921) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AND2x2_ASAP7_75t_L g816 ( .A(n_796), .B(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g859 ( .A(n_796), .Y(n_859) );
INVxp67_ASAP7_75t_SL g797 ( .A(n_798), .Y(n_797) );
OAI211xp5_ASAP7_75t_L g828 ( .A1(n_798), .A2(n_829), .B(n_830), .C(n_836), .Y(n_828) );
AOI221xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_815), .B1(n_816), .B2(n_818), .C(n_819), .Y(n_798) );
OAI21xp33_ASAP7_75t_SL g799 ( .A1(n_800), .A2(n_803), .B(n_805), .Y(n_799) );
AND2x2_ASAP7_75t_L g857 ( .A(n_802), .B(n_823), .Y(n_857) );
OR2x2_ASAP7_75t_L g898 ( .A(n_802), .B(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g890 ( .A(n_803), .Y(n_890) );
A2O1A1Ixp33_ASAP7_75t_L g851 ( .A1(n_805), .A2(n_852), .B(n_855), .C(n_858), .Y(n_851) );
INVx2_ASAP7_75t_L g874 ( .A(n_805), .Y(n_874) );
BUFx3_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g850 ( .A(n_806), .Y(n_850) );
AOI21xp5_ASAP7_75t_L g866 ( .A1(n_806), .A2(n_867), .B(n_868), .Y(n_866) );
AOI31xp33_ASAP7_75t_L g918 ( .A1(n_806), .A2(n_919), .A3(n_924), .B(n_928), .Y(n_918) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
OAI22xp33_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_809) );
HB1xp67_ASAP7_75t_L g932 ( .A(n_813), .Y(n_932) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g891 ( .A(n_815), .Y(n_891) );
INVx1_ASAP7_75t_L g895 ( .A(n_816), .Y(n_895) );
AND2x2_ASAP7_75t_L g902 ( .A(n_816), .B(n_827), .Y(n_902) );
AOI21xp33_ASAP7_75t_L g871 ( .A1(n_817), .A2(n_872), .B(n_874), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_818), .B(n_917), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_821), .B1(n_824), .B2(n_826), .Y(n_819) );
INVx1_ASAP7_75t_L g927 ( .A(n_820), .Y(n_927) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g873 ( .A(n_823), .Y(n_873) );
NAND2xp5_ASAP7_75t_SL g900 ( .A(n_824), .B(n_901), .Y(n_900) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
AOI221xp5_ASAP7_75t_L g919 ( .A1(n_825), .A2(n_837), .B1(n_838), .B2(n_920), .C(n_921), .Y(n_919) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
OAI21xp5_ASAP7_75t_L g870 ( .A1(n_831), .A2(n_833), .B(n_838), .Y(n_870) );
INVx1_ASAP7_75t_L g854 ( .A(n_832), .Y(n_854) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
O2A1O1Ixp33_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_838), .B(n_840), .C(n_841), .Y(n_836) );
NAND2xp5_ASAP7_75t_SL g886 ( .A(n_839), .B(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g901 ( .A(n_840), .Y(n_901) );
INVx1_ASAP7_75t_L g925 ( .A(n_842), .Y(n_925) );
AND2x2_ASAP7_75t_L g845 ( .A(n_846), .B(n_847), .Y(n_845) );
AOI331xp33_ASAP7_75t_L g861 ( .A1(n_848), .A2(n_862), .A3(n_864), .B1(n_866), .B2(n_870), .B3(n_871), .C1(n_875), .Y(n_861) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVxp67_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g887 ( .A(n_857), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_863), .B(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g876 ( .A(n_877), .B(n_878), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_891), .B(n_892), .Y(n_879) );
INVx1_ASAP7_75t_L g911 ( .A(n_882), .Y(n_911) );
AOI21xp5_ASAP7_75t_SL g885 ( .A1(n_886), .A2(n_888), .B(n_889), .Y(n_885) );
OAI21xp33_ASAP7_75t_L g914 ( .A1(n_887), .A2(n_915), .B(n_916), .Y(n_914) );
OAI211xp5_ASAP7_75t_SL g892 ( .A1(n_893), .A2(n_895), .B(n_896), .C(n_903), .Y(n_892) );
INVx1_ASAP7_75t_L g913 ( .A(n_893), .Y(n_913) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g926 ( .A(n_908), .Y(n_926) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
BUFx2_ASAP7_75t_SL g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
NAND4xp25_ASAP7_75t_L g936 ( .A(n_937), .B(n_971), .C(n_994), .D(n_1015), .Y(n_936) );
OAI21xp5_ASAP7_75t_L g937 ( .A1(n_938), .A2(n_964), .B(n_969), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_939), .B(n_956), .Y(n_938) );
NOR2xp33_ASAP7_75t_SL g939 ( .A(n_940), .B(n_953), .Y(n_939) );
INVx2_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
AOI22xp5_ASAP7_75t_L g944 ( .A1(n_945), .A2(n_946), .B1(n_950), .B2(n_951), .Y(n_944) );
AND2x2_ASAP7_75t_L g946 ( .A(n_947), .B(n_948), .Y(n_946) );
INVx1_ASAP7_75t_SL g963 ( .A(n_947), .Y(n_963) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g955 ( .A(n_952), .Y(n_955) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g966 ( .A(n_955), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_957), .A2(n_958), .B1(n_961), .B2(n_962), .Y(n_956) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
CKINVDCx6p67_ASAP7_75t_R g967 ( .A(n_968), .Y(n_967) );
AO21x1_ASAP7_75t_SL g971 ( .A1(n_972), .A2(n_985), .B(n_992), .Y(n_971) );
NOR3xp33_ASAP7_75t_L g972 ( .A(n_973), .B(n_978), .C(n_982), .Y(n_972) );
NOR2xp33_ASAP7_75t_L g1037 ( .A(n_974), .B(n_1038), .Y(n_1037) );
AND2x4_ASAP7_75t_L g989 ( .A(n_977), .B(n_990), .Y(n_989) );
INVx2_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_986), .A2(n_987), .B1(n_988), .B2(n_989), .Y(n_985) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVxp67_ASAP7_75t_L g1038 ( .A(n_993), .Y(n_1038) );
AOI33xp33_ASAP7_75t_L g1281 ( .A1(n_995), .A2(n_1282), .A3(n_1284), .B1(n_1286), .B2(n_1287), .B3(n_1288), .Y(n_1281) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
INVx2_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
HB1xp67_ASAP7_75t_L g1352 ( .A(n_1006), .Y(n_1352) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
INVx2_ASAP7_75t_L g1620 ( .A(n_1007), .Y(n_1620) );
BUFx3_ASAP7_75t_L g1156 ( .A(n_1009), .Y(n_1156) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1011), .Y(n_1270) );
AOI33xp33_ASAP7_75t_L g1015 ( .A1(n_1016), .A2(n_1019), .A3(n_1023), .B1(n_1026), .B2(n_1027), .B3(n_1028), .Y(n_1015) );
INVx2_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
CKINVDCx5p33_ASAP7_75t_R g1566 ( .A(n_1017), .Y(n_1566) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1022), .Y(n_1227) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1022), .Y(n_1386) );
AOI33xp33_ASAP7_75t_L g1565 ( .A1(n_1028), .A2(n_1566), .A3(n_1567), .B1(n_1569), .B2(n_1572), .B3(n_1575), .Y(n_1565) );
BUFx4f_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
BUFx3_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
BUFx2_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
AND2x4_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1037), .Y(n_1032) );
AND2x4_ASAP7_75t_L g1639 ( .A(n_1033), .B(n_1640), .Y(n_1639) );
NOR2xp33_ASAP7_75t_SL g1033 ( .A(n_1034), .B(n_1035), .Y(n_1033) );
INVx1_ASAP7_75t_SL g1042 ( .A(n_1034), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1110 ( .A(n_1034), .B(n_1035), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_1035), .B(n_1042), .Y(n_1041) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1037), .Y(n_1640) );
INVx2_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
CKINVDCx5p33_ASAP7_75t_R g1040 ( .A(n_1041), .Y(n_1040) );
OAI21xp5_ASAP7_75t_L g1108 ( .A1(n_1042), .A2(n_1109), .B(n_1110), .Y(n_1108) );
INVxp33_ASAP7_75t_SL g1043 ( .A(n_1044), .Y(n_1043) );
INVx2_ASAP7_75t_SL g1106 ( .A(n_1045), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1071), .Y(n_1045) );
OAI21xp33_ASAP7_75t_L g1046 ( .A1(n_1047), .A2(n_1061), .B(n_1070), .Y(n_1046) );
AOI22xp5_ASAP7_75t_L g1048 ( .A1(n_1049), .A2(n_1052), .B1(n_1055), .B2(n_1057), .Y(n_1048) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
OAI22xp33_ASAP7_75t_L g1099 ( .A1(n_1059), .A2(n_1100), .B1(n_1102), .B2(n_1103), .Y(n_1099) );
INVx2_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
AOI22xp5_ASAP7_75t_L g1196 ( .A1(n_1070), .A2(n_1197), .B1(n_1218), .B2(n_1219), .Y(n_1196) );
NOR2xp33_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1090), .Y(n_1071) );
INVx2_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
OAI22xp5_ASAP7_75t_L g1183 ( .A1(n_1078), .A2(n_1184), .B1(n_1187), .B2(n_1188), .Y(n_1183) );
OAI22xp5_ASAP7_75t_L g1189 ( .A1(n_1078), .A2(n_1190), .B1(n_1191), .B2(n_1192), .Y(n_1189) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx2_ASAP7_75t_SL g1411 ( .A(n_1083), .Y(n_1411) );
INVx2_ASAP7_75t_SL g1083 ( .A(n_1084), .Y(n_1083) );
OAI22xp5_ASAP7_75t_L g1266 ( .A1(n_1084), .A2(n_1087), .B1(n_1267), .B2(n_1268), .Y(n_1266) );
OAI22xp33_ASAP7_75t_L g1193 ( .A1(n_1085), .A2(n_1179), .B1(n_1194), .B2(n_1195), .Y(n_1193) );
OAI22xp5_ASAP7_75t_SL g1353 ( .A1(n_1085), .A2(n_1354), .B1(n_1356), .B2(n_1357), .Y(n_1353) );
OAI22xp33_ASAP7_75t_L g1420 ( .A1(n_1085), .A2(n_1380), .B1(n_1395), .B2(n_1411), .Y(n_1420) );
INVx2_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
INVx2_ASAP7_75t_L g1103 ( .A(n_1086), .Y(n_1103) );
INVx2_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
BUFx3_ASAP7_75t_L g1492 ( .A(n_1087), .Y(n_1492) );
BUFx6f_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1094), .Y(n_1090) );
INVx3_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
OAI22xp33_ASAP7_75t_L g1501 ( .A1(n_1103), .A2(n_1489), .B1(n_1502), .B2(n_1503), .Y(n_1501) );
BUFx2_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
AOI21xp5_ASAP7_75t_L g1635 ( .A1(n_1111), .A2(n_1636), .B(n_1637), .Y(n_1635) );
AOI22xp33_ASAP7_75t_SL g1111 ( .A1(n_1112), .A2(n_1113), .B1(n_1473), .B2(n_1634), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
OAI21x1_ASAP7_75t_L g1113 ( .A1(n_1114), .A2(n_1421), .B(n_1472), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
OR2x2_ASAP7_75t_L g1472 ( .A(n_1115), .B(n_1422), .Y(n_1472) );
XNOR2xp5_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1220), .Y(n_1115) );
XOR2x2_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1163), .Y(n_1116) );
XNOR2xp5_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1162), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1142), .Y(n_1118) );
INVx2_ASAP7_75t_L g1247 ( .A(n_1120), .Y(n_1247) );
OAI31xp33_ASAP7_75t_L g1301 ( .A1(n_1120), .A2(n_1302), .A3(n_1303), .B(n_1317), .Y(n_1301) );
NAND3xp33_ASAP7_75t_SL g1121 ( .A(n_1122), .B(n_1131), .C(n_1138), .Y(n_1121) );
HB1xp67_ASAP7_75t_L g1514 ( .A(n_1130), .Y(n_1514) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1133), .Y(n_1394) );
AND4x1_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1146), .C(n_1157), .D(n_1159), .Y(n_1142) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1148), .Y(n_1603) );
INVx2_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
OAI22xp5_ASAP7_75t_L g1419 ( .A1(n_1153), .A2(n_1381), .B1(n_1383), .B2(n_1416), .Y(n_1419) );
INVx2_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx2_ASAP7_75t_L g1265 ( .A(n_1154), .Y(n_1265) );
INVx2_ASAP7_75t_L g1272 ( .A(n_1154), .Y(n_1272) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1154), .Y(n_1444) );
XNOR2x1_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1165), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1196), .Y(n_1165) );
NOR3xp33_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1174), .C(n_1176), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1171), .Y(n_1167) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
BUFx2_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
INVx2_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1186), .Y(n_1344) );
NAND3xp33_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1203), .C(n_1209), .Y(n_1197) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
AOI221xp5_ASAP7_75t_L g1361 ( .A1(n_1201), .A2(n_1348), .B1(n_1362), .B2(n_1363), .C(n_1364), .Y(n_1361) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1202), .Y(n_1524) );
INVx2_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
INVx2_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
INVx1_ASAP7_75t_SL g1246 ( .A(n_1215), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g1321 ( .A1(n_1215), .A2(n_1217), .B1(n_1279), .B2(n_1280), .Y(n_1321) );
INVx4_ASAP7_75t_L g1365 ( .A(n_1215), .Y(n_1365) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
INVx2_ASAP7_75t_SL g1366 ( .A(n_1217), .Y(n_1366) );
XOR2xp5_ASAP7_75t_L g1220 ( .A(n_1221), .B(n_1322), .Y(n_1220) );
XNOR2x1_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1275), .Y(n_1221) );
NOR2x1_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1248), .Y(n_1223) );
AOI21xp5_ASAP7_75t_L g1224 ( .A1(n_1225), .A2(n_1236), .B(n_1247), .Y(n_1224) );
AOI221xp5_ASAP7_75t_L g1225 ( .A1(n_1226), .A2(n_1229), .B1(n_1230), .B2(n_1232), .C(n_1235), .Y(n_1225) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1235), .Y(n_1316) );
AOI221xp5_ASAP7_75t_L g1390 ( .A1(n_1235), .A2(n_1391), .B1(n_1393), .B2(n_1394), .C(n_1395), .Y(n_1390) );
HB1xp67_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
INVx2_ASAP7_75t_SL g1243 ( .A(n_1244), .Y(n_1243) );
AOI31xp33_ASAP7_75t_L g1506 ( .A1(n_1247), .A2(n_1507), .A3(n_1517), .B(n_1532), .Y(n_1506) );
NAND4xp25_ASAP7_75t_L g1248 ( .A(n_1249), .B(n_1252), .C(n_1255), .D(n_1259), .Y(n_1248) );
AOI22xp5_ASAP7_75t_L g1332 ( .A1(n_1260), .A2(n_1294), .B1(n_1333), .B2(n_1334), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1587 ( .A(n_1261), .B(n_1588), .Y(n_1587) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1264), .Y(n_1418) );
INVx2_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1271), .Y(n_1346) );
INVx2_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
NAND3xp33_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1292), .C(n_1301), .Y(n_1276) );
AND3x1_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1281), .C(n_1290), .Y(n_1277) );
INVx2_ASAP7_75t_SL g1604 ( .A(n_1289), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1293), .B(n_1297), .Y(n_1292) );
OAI211xp5_ASAP7_75t_L g1311 ( .A1(n_1296), .A2(n_1312), .B(n_1314), .C(n_1315), .Y(n_1311) );
AOI22xp5_ASAP7_75t_L g1328 ( .A1(n_1298), .A2(n_1329), .B1(n_1330), .B2(n_1331), .Y(n_1328) );
NAND3xp33_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1311), .C(n_1316), .Y(n_1303) );
OAI211xp5_ASAP7_75t_L g1304 ( .A1(n_1305), .A2(n_1306), .B(n_1307), .C(n_1309), .Y(n_1304) );
INVx2_ASAP7_75t_SL g1512 ( .A(n_1310), .Y(n_1512) );
BUFx3_ASAP7_75t_L g1568 ( .A(n_1310), .Y(n_1568) );
BUFx3_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
OR2x6_ASAP7_75t_L g1546 ( .A(n_1313), .B(n_1543), .Y(n_1546) );
XNOR2xp5_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1375), .Y(n_1322) );
XNOR2x1_ASAP7_75t_L g1323 ( .A(n_1324), .B(n_1325), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1359), .Y(n_1325) );
NOR3xp33_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1335), .C(n_1337), .Y(n_1326) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1332), .Y(n_1327) );
OAI22xp5_ASAP7_75t_L g1341 ( .A1(n_1342), .A2(n_1343), .B1(n_1345), .B2(n_1346), .Y(n_1341) );
BUFx2_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
OAI22xp5_ASAP7_75t_SL g1347 ( .A1(n_1348), .A2(n_1349), .B1(n_1350), .B2(n_1351), .Y(n_1347) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
BUFx2_ASAP7_75t_L g1489 ( .A(n_1354), .Y(n_1489) );
OAI221xp5_ASAP7_75t_L g1621 ( .A1(n_1354), .A2(n_1491), .B1(n_1622), .B2(n_1623), .C(n_1624), .Y(n_1621) );
INVx2_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
NAND3xp33_ASAP7_75t_L g1360 ( .A(n_1361), .B(n_1367), .C(n_1372), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1376 ( .A(n_1377), .B(n_1398), .Y(n_1376) );
NAND3xp33_ASAP7_75t_SL g1378 ( .A(n_1379), .B(n_1382), .C(n_1390), .Y(n_1378) );
NOR3xp33_ASAP7_75t_L g1398 ( .A(n_1399), .B(n_1407), .C(n_1409), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1399 ( .A(n_1400), .B(n_1403), .Y(n_1399) );
OAI22xp5_ASAP7_75t_L g1414 ( .A1(n_1415), .A2(n_1416), .B1(n_1417), .B2(n_1418), .Y(n_1414) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1422), .Y(n_1421) );
HB1xp67_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1424), .Y(n_1471) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1425), .B(n_1452), .Y(n_1424) );
NOR3xp33_ASAP7_75t_L g1425 ( .A(n_1426), .B(n_1433), .C(n_1435), .Y(n_1425) );
NAND2xp5_ASAP7_75t_L g1426 ( .A(n_1427), .B(n_1430), .Y(n_1426) );
OAI22xp5_ASAP7_75t_L g1493 ( .A1(n_1442), .A2(n_1494), .B1(n_1495), .B2(n_1496), .Y(n_1493) );
INVx2_ASAP7_75t_SL g1442 ( .A(n_1443), .Y(n_1442) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
AOI31xp33_ASAP7_75t_L g1454 ( .A1(n_1455), .A2(n_1462), .A3(n_1468), .B(n_1469), .Y(n_1454) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1473), .Y(n_1634) );
AOI22xp5_ASAP7_75t_L g1473 ( .A1(n_1474), .A2(n_1533), .B1(n_1534), .B2(n_1633), .Y(n_1473) );
HB1xp67_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
INVx2_ASAP7_75t_L g1633 ( .A(n_1475), .Y(n_1633) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1504), .Y(n_1476) );
NOR3xp33_ASAP7_75t_SL g1477 ( .A(n_1478), .B(n_1485), .C(n_1486), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1478 ( .A(n_1479), .B(n_1482), .Y(n_1478) );
OAI221xp5_ASAP7_75t_L g1528 ( .A1(n_1481), .A2(n_1483), .B1(n_1529), .B2(n_1530), .C(n_1531), .Y(n_1528) );
OAI22xp33_ASAP7_75t_L g1487 ( .A1(n_1488), .A2(n_1489), .B1(n_1490), .B2(n_1491), .Y(n_1487) );
BUFx3_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1510), .Y(n_1509) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
OR2x6_ASAP7_75t_L g1564 ( .A(n_1521), .B(n_1561), .Y(n_1564) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
BUFx2_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
INVx2_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
OR2x6_ASAP7_75t_L g1542 ( .A(n_1527), .B(n_1543), .Y(n_1542) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
AND3x1_ASAP7_75t_L g1536 ( .A(n_1537), .B(n_1582), .C(n_1591), .Y(n_1536) );
NOR2xp33_ASAP7_75t_L g1537 ( .A(n_1538), .B(n_1554), .Y(n_1537) );
NAND2xp5_ASAP7_75t_L g1538 ( .A(n_1539), .B(n_1547), .Y(n_1538) );
AOI22xp33_ASAP7_75t_L g1539 ( .A1(n_1540), .A2(n_1541), .B1(n_1544), .B2(n_1545), .Y(n_1539) );
CKINVDCx6p67_ASAP7_75t_R g1541 ( .A(n_1542), .Y(n_1541) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1543), .Y(n_1550) );
CKINVDCx6p67_ASAP7_75t_R g1545 ( .A(n_1546), .Y(n_1545) );
AOI22xp33_ASAP7_75t_L g1547 ( .A1(n_1548), .A2(n_1549), .B1(n_1551), .B2(n_1552), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1552 ( .A(n_1550), .B(n_1553), .Y(n_1552) );
NAND3xp33_ASAP7_75t_SL g1554 ( .A(n_1555), .B(n_1565), .C(n_1578), .Y(n_1554) );
AOI22xp33_ASAP7_75t_L g1555 ( .A1(n_1556), .A2(n_1557), .B1(n_1562), .B2(n_1563), .Y(n_1555) );
AOI22xp33_ASAP7_75t_L g1605 ( .A1(n_1556), .A2(n_1562), .B1(n_1606), .B2(n_1608), .Y(n_1605) );
INVx2_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
NAND2x1p5_ASAP7_75t_L g1558 ( .A(n_1559), .B(n_1560), .Y(n_1558) );
INVx2_ASAP7_75t_SL g1560 ( .A(n_1561), .Y(n_1560) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1561), .Y(n_1581) );
INVx2_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
HB1xp67_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
NAND2xp5_ASAP7_75t_L g1580 ( .A(n_1571), .B(n_1581), .Y(n_1580) );
BUFx2_ASAP7_75t_L g1573 ( .A(n_1574), .Y(n_1573) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1577), .Y(n_1576) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
NAND2xp5_ASAP7_75t_L g1582 ( .A(n_1583), .B(n_1584), .Y(n_1582) );
NOR2xp67_ASAP7_75t_L g1585 ( .A(n_1586), .B(n_1587), .Y(n_1585) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
OR2x2_ASAP7_75t_L g1626 ( .A(n_1589), .B(n_1627), .Y(n_1626) );
INVx2_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
INVx8_ASAP7_75t_L g1593 ( .A(n_1594), .Y(n_1593) );
AND2x4_ASAP7_75t_L g1632 ( .A(n_1595), .B(n_1620), .Y(n_1632) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1596), .Y(n_1595) );
INVx2_ASAP7_75t_L g1598 ( .A(n_1599), .Y(n_1598) );
INVx2_ASAP7_75t_L g1599 ( .A(n_1600), .Y(n_1599) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
HB1xp67_ASAP7_75t_L g1606 ( .A(n_1607), .Y(n_1606) );
CKINVDCx11_ASAP7_75t_R g1608 ( .A(n_1609), .Y(n_1608) );
CKINVDCx6p67_ASAP7_75t_R g1611 ( .A(n_1612), .Y(n_1611) );
OAI22xp5_ASAP7_75t_SL g1613 ( .A1(n_1614), .A2(n_1615), .B1(n_1616), .B2(n_1617), .Y(n_1613) );
INVx1_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1619), .Y(n_1618) );
INVx1_ASAP7_75t_L g1619 ( .A(n_1620), .Y(n_1619) );
INVx2_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
INVx3_ASAP7_75t_L g1629 ( .A(n_1630), .Y(n_1629) );
INVx3_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
BUFx2_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
endmodule