module fake_aes_6658_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_3), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_1), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_1), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
INVx3_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_4), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_16), .B(n_0), .Y(n_18) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_16), .B(n_2), .Y(n_19) );
O2A1O1Ixp33_ASAP7_75t_SL g20 ( .A1(n_13), .A2(n_2), .B(n_3), .C(n_4), .Y(n_20) );
NAND2xp5_ASAP7_75t_SL g21 ( .A(n_16), .B(n_5), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_16), .Y(n_22) );
INVx6_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
NAND4xp25_ASAP7_75t_L g24 ( .A(n_20), .B(n_13), .C(n_16), .D(n_14), .Y(n_24) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
HB1xp67_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
AOI221xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_24), .B1(n_11), .B2(n_12), .C(n_17), .Y(n_28) );
AOI311xp33_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_18), .A3(n_15), .B(n_21), .C(n_27), .Y(n_29) );
NAND2xp5_ASAP7_75t_L g30 ( .A(n_29), .B(n_7), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_31), .B(n_7), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_30), .Y(n_33) );
AOI22xp5_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_9), .B1(n_10), .B2(n_32), .Y(n_34) );
endmodule