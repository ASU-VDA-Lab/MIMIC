module fake_aes_9396_n_652 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_652);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_652;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_613;
wire n_648;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_597;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_SL g75 ( .A(n_27), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_59), .Y(n_76) );
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_58), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_54), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_42), .Y(n_79) );
NOR2xp67_ASAP7_75t_L g80 ( .A(n_32), .B(n_45), .Y(n_80) );
NOR2xp67_ASAP7_75t_L g81 ( .A(n_35), .B(n_22), .Y(n_81) );
INVx1_ASAP7_75t_SL g82 ( .A(n_1), .Y(n_82) );
BUFx10_ASAP7_75t_L g83 ( .A(n_24), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_44), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_46), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_51), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_74), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_34), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_70), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_3), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_31), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_38), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_48), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_29), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_26), .Y(n_95) );
INVx2_ASAP7_75t_SL g96 ( .A(n_72), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_57), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_61), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_67), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_56), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_64), .Y(n_101) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_8), .Y(n_102) );
BUFx3_ASAP7_75t_L g103 ( .A(n_21), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_30), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_19), .Y(n_105) );
CKINVDCx14_ASAP7_75t_R g106 ( .A(n_37), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_53), .Y(n_107) );
INVx2_ASAP7_75t_SL g108 ( .A(n_40), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_50), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_52), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_4), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_65), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_73), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_15), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_9), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_71), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_20), .Y(n_117) );
NOR2xp67_ASAP7_75t_L g118 ( .A(n_6), .B(n_13), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_2), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_33), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_114), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_87), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_79), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_88), .B(n_0), .Y(n_124) );
XOR2xp5_ASAP7_75t_L g125 ( .A(n_115), .B(n_0), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_103), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_87), .Y(n_127) );
OAI21x1_ASAP7_75t_L g128 ( .A1(n_79), .A2(n_18), .B(n_68), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_111), .B(n_1), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_105), .B(n_2), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_90), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_131) );
OAI22xp5_ASAP7_75t_SL g132 ( .A1(n_90), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_113), .B(n_7), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_104), .Y(n_134) );
INVx6_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_111), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_106), .B(n_8), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_75), .B(n_108), .Y(n_138) );
OAI22xp5_ASAP7_75t_SL g139 ( .A1(n_119), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_139) );
OAI21x1_ASAP7_75t_L g140 ( .A1(n_110), .A2(n_36), .B(n_66), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_104), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_83), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_110), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_75), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_103), .Y(n_145) );
BUFx12f_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_120), .Y(n_147) );
INVxp67_ASAP7_75t_L g148 ( .A(n_119), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_109), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_102), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_120), .Y(n_151) );
INVxp67_ASAP7_75t_L g152 ( .A(n_102), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_96), .B(n_10), .Y(n_153) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_109), .A2(n_39), .B(n_63), .Y(n_154) );
AND2x6_ASAP7_75t_L g155 ( .A(n_116), .B(n_28), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_96), .B(n_11), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_116), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_108), .B(n_12), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_117), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_117), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_155), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_128), .Y(n_162) );
BUFx10_ASAP7_75t_L g163 ( .A(n_135), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_126), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_126), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_142), .B(n_85), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_123), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_129), .A2(n_102), .B1(n_118), .B2(n_82), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_126), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_126), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_142), .B(n_84), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_142), .B(n_77), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_138), .B(n_84), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_155), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_146), .B(n_98), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_126), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_129), .A2(n_158), .B1(n_155), .B2(n_159), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_155), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_138), .B(n_77), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_158), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_123), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_135), .B(n_112), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
INVx4_ASAP7_75t_SL g185 ( .A(n_155), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_135), .B(n_78), .Y(n_186) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_128), .A2(n_107), .B(n_101), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_143), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_121), .B(n_91), .Y(n_189) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_148), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_138), .B(n_94), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_143), .Y(n_192) );
OR2x6_ASAP7_75t_L g193 ( .A(n_131), .B(n_102), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_150), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_146), .B(n_85), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_135), .B(n_86), .Y(n_196) );
AND2x6_ASAP7_75t_L g197 ( .A(n_129), .B(n_93), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_144), .B(n_86), .Y(n_198) );
AND2x6_ASAP7_75t_L g199 ( .A(n_137), .B(n_76), .Y(n_199) );
BUFx2_ASAP7_75t_L g200 ( .A(n_137), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_155), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_144), .B(n_102), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_145), .Y(n_203) );
INVx1_ASAP7_75t_SL g204 ( .A(n_124), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_122), .B(n_94), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_150), .Y(n_206) );
NOR2xp33_ASAP7_75t_SL g207 ( .A(n_122), .B(n_98), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_150), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_145), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_151), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_145), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_151), .B(n_89), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_136), .B(n_100), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_145), .Y(n_214) );
NAND3xp33_ASAP7_75t_L g215 ( .A(n_127), .B(n_99), .C(n_97), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_204), .B(n_160), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_162), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_180), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_204), .B(n_160), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_162), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_162), .Y(n_221) );
BUFx3_ASAP7_75t_L g222 ( .A(n_178), .Y(n_222) );
NAND2xp33_ASAP7_75t_SL g223 ( .A(n_161), .B(n_153), .Y(n_223) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_189), .Y(n_224) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_189), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_196), .B(n_133), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_196), .B(n_159), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_199), .A2(n_157), .B1(n_141), .B2(n_127), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_173), .B(n_157), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_179), .B(n_134), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_162), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_180), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_191), .B(n_134), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_166), .B(n_141), .Y(n_234) );
OAI22xp5_ASAP7_75t_SL g235 ( .A1(n_193), .A2(n_125), .B1(n_132), .B2(n_139), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_199), .A2(n_149), .B1(n_156), .B2(n_130), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_200), .B(n_149), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_199), .A2(n_89), .B1(n_91), .B2(n_95), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_162), .Y(n_239) );
AND2x2_ASAP7_75t_SL g240 ( .A(n_161), .B(n_154), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_190), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_180), .Y(n_242) );
NAND2xp33_ASAP7_75t_L g243 ( .A(n_197), .B(n_92), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_178), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_180), .Y(n_245) );
BUFx2_ASAP7_75t_L g246 ( .A(n_199), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_199), .A2(n_152), .B1(n_147), .B2(n_81), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_171), .B(n_147), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_164), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_200), .Y(n_250) );
INVx2_ASAP7_75t_SL g251 ( .A(n_163), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_207), .B(n_147), .Y(n_252) );
NAND2x1p5_ASAP7_75t_L g253 ( .A(n_161), .B(n_140), .Y(n_253) );
AND2x6_ASAP7_75t_SL g254 ( .A(n_193), .B(n_125), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_172), .B(n_147), .Y(n_255) );
BUFx3_ASAP7_75t_L g256 ( .A(n_178), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_177), .A2(n_147), .B1(n_80), .B2(n_154), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_207), .B(n_140), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_164), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_161), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_184), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_174), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_199), .A2(n_154), .B1(n_13), .B2(n_14), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_199), .A2(n_154), .B1(n_14), .B2(n_15), .Y(n_264) );
INVxp67_ASAP7_75t_SL g265 ( .A(n_184), .Y(n_265) );
OR2x2_ASAP7_75t_L g266 ( .A(n_193), .B(n_12), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_174), .B(n_47), .Y(n_267) );
NOR2x1p5_ASAP7_75t_L g268 ( .A(n_193), .B(n_16), .Y(n_268) );
AO22x1_ASAP7_75t_L g269 ( .A1(n_197), .A2(n_16), .B1(n_17), .B2(n_23), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_212), .B(n_25), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_202), .Y(n_271) );
NOR2x2_ASAP7_75t_L g272 ( .A(n_193), .B(n_69), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_197), .A2(n_41), .B1(n_43), .B2(n_49), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_205), .B(n_62), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_216), .B(n_197), .Y(n_275) );
NOR2xp67_ASAP7_75t_SL g276 ( .A(n_260), .B(n_201), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_219), .A2(n_184), .B1(n_168), .B2(n_174), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_224), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_234), .A2(n_184), .B(n_213), .C(n_215), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_225), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_229), .A2(n_215), .B(n_186), .C(n_183), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_228), .A2(n_174), .B1(n_201), .B2(n_198), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g283 ( .A(n_241), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_241), .A2(n_197), .B1(n_175), .B2(n_195), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_218), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_222), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_268), .A2(n_197), .B1(n_202), .B2(n_192), .Y(n_287) );
INVx4_ASAP7_75t_L g288 ( .A(n_246), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_218), .Y(n_289) );
O2A1O1Ixp33_ASAP7_75t_L g290 ( .A1(n_227), .A2(n_188), .B(n_192), .C(n_181), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_246), .A2(n_201), .B1(n_210), .B2(n_181), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_250), .B(n_201), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_232), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_250), .B(n_226), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_251), .B(n_163), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_258), .A2(n_187), .B(n_210), .Y(n_296) );
OAI21xp33_ASAP7_75t_SL g297 ( .A1(n_232), .A2(n_188), .B(n_167), .Y(n_297) );
O2A1O1Ixp33_ASAP7_75t_L g298 ( .A1(n_230), .A2(n_167), .B(n_202), .C(n_210), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_226), .A2(n_197), .B1(n_163), .B2(n_210), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_226), .B(n_163), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_237), .B(n_202), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_251), .B(n_185), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_222), .B(n_185), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_237), .B(n_185), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_254), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_233), .B(n_185), .Y(n_306) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_257), .A2(n_208), .B(n_206), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_242), .Y(n_308) );
O2A1O1Ixp33_ASAP7_75t_L g309 ( .A1(n_266), .A2(n_187), .B(n_208), .C(n_206), .Y(n_309) );
OR2x6_ASAP7_75t_L g310 ( .A(n_266), .B(n_182), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_256), .B(n_194), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_271), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_272), .Y(n_313) );
A2O1A1Ixp33_ASAP7_75t_L g314 ( .A1(n_242), .A2(n_194), .B(n_211), .C(n_165), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_236), .B(n_187), .Y(n_315) );
A2O1A1Ixp33_ASAP7_75t_SL g316 ( .A1(n_255), .A2(n_176), .B(n_211), .C(n_165), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_256), .B(n_176), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_245), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_238), .B(n_182), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_245), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_283), .Y(n_321) );
O2A1O1Ixp33_ASAP7_75t_L g322 ( .A1(n_279), .A2(n_261), .B(n_243), .C(n_248), .Y(n_322) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_278), .A2(n_235), .B1(n_261), .B2(n_265), .C(n_264), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_294), .B(n_247), .Y(n_324) );
NAND3xp33_ASAP7_75t_SL g325 ( .A(n_313), .B(n_263), .C(n_274), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_280), .B(n_243), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_301), .Y(n_327) );
INVxp67_ASAP7_75t_L g328 ( .A(n_300), .Y(n_328) );
NOR4xp25_ASAP7_75t_L g329 ( .A(n_309), .B(n_272), .C(n_252), .D(n_273), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_286), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_310), .B(n_269), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_318), .Y(n_332) );
NAND2x1p5_ASAP7_75t_L g333 ( .A(n_288), .B(n_286), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g334 ( .A1(n_281), .A2(n_270), .B(n_267), .C(n_253), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_320), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_285), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_289), .Y(n_337) );
A2O1A1Ixp33_ASAP7_75t_L g338 ( .A1(n_290), .A2(n_223), .B(n_240), .C(n_262), .Y(n_338) );
OAI21xp5_ASAP7_75t_L g339 ( .A1(n_315), .A2(n_253), .B(n_223), .Y(n_339) );
INVx1_ASAP7_75t_SL g340 ( .A(n_310), .Y(n_340) );
INVx5_ASAP7_75t_L g341 ( .A(n_286), .Y(n_341) );
XOR2xp5_ASAP7_75t_L g342 ( .A(n_305), .B(n_269), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_310), .A2(n_221), .B1(n_239), .B2(n_231), .Y(n_343) );
OAI21xp5_ASAP7_75t_L g344 ( .A1(n_309), .A2(n_253), .B(n_240), .Y(n_344) );
O2A1O1Ixp33_ASAP7_75t_L g345 ( .A1(n_298), .A2(n_220), .B(n_239), .C(n_231), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_284), .B(n_260), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_287), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_287), .A2(n_217), .B1(n_221), .B2(n_220), .Y(n_348) );
O2A1O1Ixp33_ASAP7_75t_L g349 ( .A1(n_298), .A2(n_217), .B(n_262), .C(n_169), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_321), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_334), .A2(n_296), .B(n_316), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_321), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_328), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_344), .A2(n_297), .B(n_290), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_332), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_335), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_336), .Y(n_357) );
BUFx10_ASAP7_75t_L g358 ( .A(n_327), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_335), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_347), .A2(n_293), .B1(n_308), .B2(n_319), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_343), .A2(n_275), .B(n_306), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_339), .A2(n_307), .B(n_314), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_337), .Y(n_363) );
AOI22xp33_ASAP7_75t_SL g364 ( .A1(n_347), .A2(n_288), .B1(n_292), .B2(n_277), .Y(n_364) );
INVxp67_ASAP7_75t_L g365 ( .A(n_326), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_338), .A2(n_317), .B(n_303), .Y(n_366) );
AO31x2_ASAP7_75t_L g367 ( .A1(n_338), .A2(n_209), .A3(n_214), .B(n_169), .Y(n_367) );
OAI21x1_ASAP7_75t_SL g368 ( .A1(n_345), .A2(n_299), .B(n_304), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_340), .B(n_312), .Y(n_369) );
O2A1O1Ixp33_ASAP7_75t_L g370 ( .A1(n_324), .A2(n_282), .B(n_291), .C(n_311), .Y(n_370) );
AO21x2_ASAP7_75t_L g371 ( .A1(n_329), .A2(n_302), .B(n_214), .Y(n_371) );
OAI221xp5_ASAP7_75t_L g372 ( .A1(n_323), .A2(n_295), .B1(n_286), .B2(n_170), .C(n_203), .Y(n_372) );
A2O1A1Ixp33_ASAP7_75t_L g373 ( .A1(n_322), .A2(n_209), .B(n_203), .C(n_170), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_348), .A2(n_249), .B(n_259), .Y(n_374) );
AOI22xp33_ASAP7_75t_SL g375 ( .A1(n_331), .A2(n_346), .B1(n_342), .B2(n_333), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_356), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_356), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_359), .Y(n_378) );
AOI31xp33_ASAP7_75t_L g379 ( .A1(n_375), .A2(n_333), .A3(n_325), .B(n_346), .Y(n_379) );
OR2x6_ASAP7_75t_L g380 ( .A(n_354), .B(n_368), .Y(n_380) );
AO21x2_ASAP7_75t_L g381 ( .A1(n_351), .A2(n_349), .B(n_259), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_359), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g383 ( .A1(n_360), .A2(n_330), .B1(n_341), .B2(n_276), .C(n_249), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_367), .Y(n_384) );
OA21x2_ASAP7_75t_L g385 ( .A1(n_362), .A2(n_330), .B(n_341), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_355), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_357), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_358), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_367), .Y(n_389) );
BUFx2_ASAP7_75t_L g390 ( .A(n_369), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_367), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_363), .B(n_341), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_360), .B(n_330), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_371), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_352), .B(n_341), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_365), .A2(n_55), .B1(n_60), .B2(n_244), .C(n_353), .Y(n_396) );
INVxp67_ASAP7_75t_SL g397 ( .A(n_374), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_358), .B(n_244), .Y(n_398) );
OA21x2_ASAP7_75t_L g399 ( .A1(n_373), .A2(n_244), .B(n_366), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_358), .B(n_244), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_367), .Y(n_401) );
AO21x2_ASAP7_75t_L g402 ( .A1(n_373), .A2(n_244), .B(n_371), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_371), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_374), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_369), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_364), .A2(n_350), .B1(n_372), .B2(n_361), .Y(n_406) );
OA21x2_ASAP7_75t_L g407 ( .A1(n_370), .A2(n_351), .B(n_354), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_356), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_390), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_377), .Y(n_410) );
INVx2_ASAP7_75t_SL g411 ( .A(n_388), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_377), .Y(n_412) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_376), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_376), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_378), .Y(n_415) );
BUFx3_ASAP7_75t_L g416 ( .A(n_388), .Y(n_416) );
INVx3_ASAP7_75t_L g417 ( .A(n_385), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_395), .B(n_390), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_378), .Y(n_419) );
AO21x2_ASAP7_75t_L g420 ( .A1(n_404), .A2(n_397), .B(n_381), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_382), .B(n_408), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_382), .B(n_408), .Y(n_422) );
BUFx2_ASAP7_75t_L g423 ( .A(n_388), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_386), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_405), .B(n_386), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_405), .B(n_387), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_405), .B(n_387), .Y(n_427) );
INVx5_ASAP7_75t_SL g428 ( .A(n_380), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_385), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_380), .B(n_401), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_392), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_385), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_385), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_385), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_392), .B(n_379), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_384), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_384), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_384), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_380), .B(n_401), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_389), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_389), .Y(n_441) );
AO21x2_ASAP7_75t_L g442 ( .A1(n_404), .A2(n_397), .B(n_381), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_393), .B(n_380), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_389), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_391), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_380), .B(n_401), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_407), .B(n_380), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_379), .B(n_406), .Y(n_448) );
AO21x2_ASAP7_75t_L g449 ( .A1(n_381), .A2(n_391), .B(n_403), .Y(n_449) );
INVx4_ASAP7_75t_L g450 ( .A(n_398), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_391), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_403), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_403), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_407), .B(n_393), .Y(n_454) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_383), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_454), .B(n_394), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_415), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_418), .B(n_406), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_454), .B(n_394), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_415), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_447), .B(n_407), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_447), .B(n_407), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_412), .B(n_407), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_425), .B(n_396), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_452), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_412), .B(n_402), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_425), .B(n_402), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_419), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_416), .Y(n_469) );
OR2x6_ASAP7_75t_L g470 ( .A(n_423), .B(n_399), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_419), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_410), .B(n_402), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_424), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_426), .B(n_396), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_424), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_426), .B(n_402), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_452), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_421), .B(n_399), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_416), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_421), .B(n_399), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_410), .B(n_399), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_409), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_453), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_422), .B(n_399), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_422), .B(n_381), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_414), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_414), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_443), .B(n_398), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_413), .B(n_383), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_453), .Y(n_490) );
HB1xp67_ASAP7_75t_SL g491 ( .A(n_423), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_427), .B(n_400), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_443), .B(n_400), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_436), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_431), .B(n_448), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_430), .B(n_446), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_430), .B(n_446), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_436), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_431), .B(n_435), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_430), .B(n_439), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_437), .Y(n_501) );
INVx3_ASAP7_75t_L g502 ( .A(n_417), .Y(n_502) );
NAND4xp25_ASAP7_75t_L g503 ( .A(n_430), .B(n_439), .C(n_446), .D(n_417), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_437), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_438), .Y(n_505) );
INVxp67_ASAP7_75t_SL g506 ( .A(n_411), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_438), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_440), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_411), .B(n_450), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_439), .B(n_446), .Y(n_510) );
AND2x2_ASAP7_75t_SL g511 ( .A(n_489), .B(n_450), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_482), .B(n_450), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_499), .B(n_495), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_473), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_461), .B(n_439), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_473), .B(n_450), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_492), .B(n_440), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_475), .B(n_455), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_475), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_500), .B(n_417), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_457), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_465), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_458), .B(n_434), .C(n_432), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_465), .Y(n_524) );
INVx3_ASAP7_75t_L g525 ( .A(n_502), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_488), .B(n_451), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_457), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_460), .B(n_451), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_488), .B(n_441), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_461), .B(n_462), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_460), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_468), .B(n_445), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_462), .B(n_428), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_456), .B(n_428), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_468), .B(n_445), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_456), .B(n_428), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_471), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_471), .B(n_441), .Y(n_538) );
BUFx3_ASAP7_75t_L g539 ( .A(n_469), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_479), .B(n_444), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_491), .B(n_444), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_494), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_509), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_493), .B(n_428), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_494), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_459), .B(n_428), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_501), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_493), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_459), .B(n_429), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_506), .B(n_434), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_501), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_500), .B(n_417), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_496), .B(n_429), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_500), .B(n_432), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_464), .B(n_433), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_504), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_504), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_486), .B(n_433), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_485), .B(n_449), .Y(n_559) );
OAI31xp33_ASAP7_75t_L g560 ( .A1(n_503), .A2(n_420), .A3(n_442), .B(n_449), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_555), .B(n_485), .Y(n_561) );
NAND2x1p5_ASAP7_75t_L g562 ( .A(n_511), .B(n_489), .Y(n_562) );
AOI21xp33_ASAP7_75t_SL g563 ( .A1(n_511), .A2(n_474), .B(n_502), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_530), .B(n_510), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_555), .B(n_463), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_549), .B(n_463), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_548), .B(n_467), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_530), .B(n_510), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_549), .B(n_476), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_526), .B(n_476), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_523), .A2(n_541), .B(n_560), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_514), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_518), .B(n_467), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_513), .B(n_484), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_529), .B(n_497), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_559), .B(n_497), .Y(n_576) );
NOR2xp67_ASAP7_75t_SL g577 ( .A(n_539), .B(n_502), .Y(n_577) );
INVxp67_ASAP7_75t_L g578 ( .A(n_539), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_517), .B(n_496), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_519), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_521), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_527), .Y(n_582) );
OR2x6_ASAP7_75t_L g583 ( .A(n_541), .B(n_470), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_543), .B(n_484), .Y(n_584) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_550), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_531), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_553), .B(n_487), .Y(n_587) );
NOR2xp33_ASAP7_75t_SL g588 ( .A(n_512), .B(n_502), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g589 ( .A1(n_537), .A2(n_466), .B1(n_478), .B2(n_480), .C(n_507), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_542), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_545), .B(n_480), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_547), .B(n_505), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_558), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g594 ( .A(n_540), .B(n_507), .C(n_505), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_515), .B(n_487), .Y(n_595) );
AOI21xp33_ASAP7_75t_L g596 ( .A1(n_578), .A2(n_516), .B(n_525), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_585), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_572), .Y(n_598) );
AND2x2_ASAP7_75t_SL g599 ( .A(n_588), .B(n_520), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_571), .A2(n_515), .B1(n_554), .B2(n_552), .C(n_520), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_589), .B(n_554), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_587), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_593), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_580), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_595), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_561), .B(n_554), .Y(n_606) );
AOI322xp5_ASAP7_75t_L g607 ( .A1(n_565), .A2(n_533), .A3(n_546), .B1(n_534), .B2(n_536), .C1(n_520), .C2(n_552), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_562), .A2(n_533), .B1(n_552), .B2(n_536), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_581), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_582), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_574), .B(n_544), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_573), .B(n_557), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_579), .B(n_556), .Y(n_613) );
OAI21xp5_ASAP7_75t_SL g614 ( .A1(n_562), .A2(n_546), .B(n_534), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_563), .A2(n_538), .B(n_535), .Y(n_615) );
OAI211xp5_ASAP7_75t_SL g616 ( .A1(n_591), .A2(n_525), .B(n_551), .C(n_528), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g617 ( .A1(n_583), .A2(n_470), .B(n_525), .C(n_532), .Y(n_617) );
AOI222xp33_ASAP7_75t_L g618 ( .A1(n_600), .A2(n_594), .B1(n_584), .B2(n_590), .C1(n_586), .C2(n_566), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_615), .B(n_576), .Y(n_619) );
OAI211xp5_ASAP7_75t_SL g620 ( .A1(n_607), .A2(n_569), .B(n_567), .C(n_570), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_597), .Y(n_621) );
OAI21xp33_ASAP7_75t_L g622 ( .A1(n_601), .A2(n_588), .B(n_583), .Y(n_622) );
OAI22xp33_ASAP7_75t_L g623 ( .A1(n_614), .A2(n_583), .B1(n_594), .B2(n_575), .Y(n_623) );
INVxp67_ASAP7_75t_L g624 ( .A(n_598), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_599), .B(n_568), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_603), .B(n_564), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_602), .B(n_605), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_604), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_616), .A2(n_500), .B1(n_466), .B2(n_478), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_609), .Y(n_630) );
AOI321xp33_ASAP7_75t_L g631 ( .A1(n_623), .A2(n_617), .A3(n_608), .B1(n_596), .B2(n_613), .C(n_611), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_623), .A2(n_616), .B1(n_610), .B2(n_606), .Y(n_632) );
OAI221xp5_ASAP7_75t_L g633 ( .A1(n_622), .A2(n_617), .B1(n_612), .B2(n_577), .C(n_592), .Y(n_633) );
AOI221x1_ASAP7_75t_L g634 ( .A1(n_620), .A2(n_592), .B1(n_486), .B2(n_522), .C(n_524), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g635 ( .A1(n_619), .A2(n_481), .B(n_472), .C(n_524), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_618), .A2(n_522), .B(n_470), .Y(n_636) );
AOI211xp5_ASAP7_75t_L g637 ( .A1(n_627), .A2(n_481), .B(n_472), .C(n_483), .Y(n_637) );
INVx1_ASAP7_75t_SL g638 ( .A(n_632), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_634), .B(n_624), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_636), .B(n_625), .Y(n_640) );
OAI211xp5_ASAP7_75t_SL g641 ( .A1(n_631), .A2(n_629), .B(n_621), .C(n_628), .Y(n_641) );
NOR2xp67_ASAP7_75t_L g642 ( .A(n_639), .B(n_633), .Y(n_642) );
AND5x1_ASAP7_75t_L g643 ( .A(n_638), .B(n_635), .C(n_637), .D(n_629), .E(n_626), .Y(n_643) );
NAND4xp75_ASAP7_75t_L g644 ( .A(n_640), .B(n_626), .C(n_630), .D(n_483), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_642), .B(n_641), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_644), .A2(n_470), .B1(n_420), .B2(n_442), .Y(n_646) );
AOI22x1_ASAP7_75t_L g647 ( .A1(n_645), .A2(n_643), .B1(n_477), .B2(n_483), .Y(n_647) );
OAI22xp5_ASAP7_75t_SL g648 ( .A1(n_647), .A2(n_646), .B1(n_470), .B2(n_498), .Y(n_648) );
OAI22x1_ASAP7_75t_L g649 ( .A1(n_648), .A2(n_477), .B1(n_490), .B2(n_465), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_649), .A2(n_477), .B(n_490), .Y(n_650) );
AOI21xp33_ASAP7_75t_SL g651 ( .A1(n_650), .A2(n_420), .B(n_442), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_651), .A2(n_490), .B1(n_498), .B2(n_508), .C(n_449), .Y(n_652) );
endmodule