module fake_jpeg_5327_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_43),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_37),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_29),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_40),
.B(n_27),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_47),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_29),
.B(n_32),
.Y(n_71)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_18),
.Y(n_79)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_48),
.Y(n_57)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_53),
.Y(n_97)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_56),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_16),
.B1(n_25),
.B2(n_26),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_55),
.A2(n_74),
.B1(n_93),
.B2(n_28),
.Y(n_117)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_25),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_58),
.B(n_61),
.Y(n_107)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_59),
.B(n_60),
.Y(n_123)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_33),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_76),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_65),
.B(n_66),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

CKINVDCx12_ASAP7_75t_R g69 ( 
.A(n_36),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_69),
.B(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_28),
.B(n_21),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_19),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_78),
.Y(n_104)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_45),
.A2(n_26),
.B1(n_24),
.B2(n_22),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_38),
.A2(n_18),
.B1(n_32),
.B2(n_31),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_75),
.A2(n_85),
.B1(n_89),
.B2(n_92),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_38),
.B(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_39),
.B(n_17),
.Y(n_77)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_22),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_87),
.Y(n_111)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_41),
.B(n_23),
.Y(n_81)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g85 ( 
.A(n_37),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_37),
.B(n_34),
.Y(n_87)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_41),
.B(n_34),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_94),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_43),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_41),
.A2(n_31),
.B1(n_28),
.B2(n_21),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

AOI211xp5_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_30),
.B(n_4),
.C(n_5),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_96),
.A2(n_86),
.B1(n_49),
.B2(n_50),
.Y(n_146)
);

NOR3xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_95),
.C(n_94),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_95),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_21),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_121),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_120),
.A2(n_71),
.B1(n_60),
.B2(n_59),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_27),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_23),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_122),
.B(n_62),
.Y(n_140)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_129),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_67),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_126),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_127),
.A2(n_134),
.B1(n_142),
.B2(n_146),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_82),
.B(n_73),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_128),
.A2(n_150),
.B(n_156),
.Y(n_179)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_55),
.B1(n_76),
.B2(n_87),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_131),
.A2(n_138),
.B1(n_112),
.B2(n_98),
.Y(n_162)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_76),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_143),
.Y(n_183)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_135),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_109),
.Y(n_136)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_62),
.Y(n_137)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_90),
.B1(n_68),
.B2(n_64),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_89),
.Y(n_141)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_53),
.B1(n_52),
.B2(n_90),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_51),
.Y(n_147)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_80),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_120),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_86),
.B(n_49),
.C(n_63),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_115),
.B1(n_108),
.B2(n_102),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_99),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_152),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_8),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_153),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_9),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_155),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_104),
.B(n_10),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_134),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_98),
.C(n_105),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_175),
.C(n_176),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_174),
.Y(n_192)
);

AND2x6_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_108),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_SL g199 ( 
.A(n_164),
.B(n_152),
.C(n_139),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_108),
.B(n_106),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_173),
.A2(n_184),
.B(n_150),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_100),
.C(n_106),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_114),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_155),
.A2(n_102),
.B1(n_103),
.B2(n_100),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_150),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_114),
.B(n_101),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_129),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_186),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_173),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_161),
.A2(n_135),
.B1(n_101),
.B2(n_125),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_189),
.A2(n_193),
.B(n_201),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_134),
.B1(n_138),
.B2(n_148),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_191),
.B1(n_206),
.B2(n_162),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_164),
.A2(n_146),
.B1(n_127),
.B2(n_144),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_185),
.A2(n_103),
.B1(n_132),
.B2(n_136),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_194),
.B(n_203),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_139),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_202),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_199),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_163),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_140),
.C(n_137),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_167),
.C(n_158),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_172),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_204),
.B(n_195),
.Y(n_212)
);

NOR3xp33_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_126),
.C(n_153),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_160),
.A2(n_179),
.B1(n_171),
.B2(n_181),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_179),
.B(n_183),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_208),
.A2(n_211),
.B(n_224),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_217),
.C(n_187),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_172),
.B(n_185),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_204),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_171),
.B1(n_165),
.B2(n_180),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_222),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_197),
.B(n_170),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_194),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_190),
.A2(n_180),
.B1(n_170),
.B2(n_165),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_221),
.B(n_196),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_199),
.A2(n_184),
.B(n_169),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_229),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_227),
.B(n_228),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_216),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_232),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_234),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_187),
.C(n_191),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_224),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_211),
.Y(n_242)
);

OA21x2_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_192),
.B(n_206),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_237),
.A2(n_219),
.B1(n_218),
.B2(n_168),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_214),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_230),
.C(n_236),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_246),
.B(n_247),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_225),
.A2(n_207),
.B1(n_208),
.B2(n_219),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_237),
.Y(n_253)
);

OA22x2_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_223),
.B1(n_222),
.B2(n_207),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_245),
.A2(n_237),
.B1(n_217),
.B2(n_200),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_248),
.A2(n_249),
.B(n_252),
.Y(n_256)
);

XNOR2x1_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_236),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_218),
.Y(n_250)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_231),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_253),
.B(n_241),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_214),
.C(n_209),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_244),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_255),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_261),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_254),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_249),
.A2(n_245),
.B(n_247),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_263),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_259),
.A2(n_248),
.B1(n_251),
.B2(n_186),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_256),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_264),
.B(n_257),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_267),
.A2(n_266),
.B(n_166),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_262),
.A2(n_166),
.B(n_169),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_268),
.B(n_177),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_270),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_154),
.Y(n_272)
);


endmodule