module real_jpeg_12158_n_12 (n_5, n_4, n_8, n_0, n_256, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_256;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_3),
.A2(n_53),
.B1(n_55),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_3),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_65),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_65),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_65),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_42),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_6),
.A2(n_42),
.B1(n_59),
.B2(n_60),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_9),
.A2(n_31),
.B1(n_39),
.B2(n_40),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_9),
.A2(n_31),
.B1(n_59),
.B2(n_60),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_9),
.A2(n_31),
.B1(n_53),
.B2(n_55),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_10),
.A2(n_26),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_10),
.A2(n_26),
.B1(n_59),
.B2(n_60),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_10),
.A2(n_26),
.B1(n_39),
.B2(n_40),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_10),
.B(n_97),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_10),
.B(n_25),
.C(n_36),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_10),
.B(n_27),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_10),
.B(n_35),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_10),
.A2(n_60),
.B(n_70),
.C(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_10),
.B(n_56),
.Y(n_192)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_123),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_122),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_103),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_16),
.B(n_103),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_79),
.C(n_86),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_17),
.A2(n_18),
.B1(n_79),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_47),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_19),
.B(n_48),
.C(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_33),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_20),
.B(n_33),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_29),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_21),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_23),
.A2(n_28),
.B(n_32),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_23),
.B(n_32),
.Y(n_157)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

AO22x1_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_25),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_28),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_25),
.B(n_154),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_26),
.A2(n_39),
.B(n_71),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_26),
.B(n_57),
.C(n_60),
.Y(n_207)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_28),
.B(n_30),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_28),
.B(n_134),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_28),
.A2(n_29),
.B(n_89),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_29),
.B(n_166),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_32),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_32),
.B(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_38),
.B(n_43),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_34),
.A2(n_83),
.B(n_95),
.Y(n_220)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_35),
.B(n_46),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_35),
.B(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_35),
.B(n_139),
.Y(n_149)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_38),
.A2(n_83),
.B(n_84),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_39),
.A2(n_40),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_40),
.B(n_147),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_43),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_43),
.B(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_44),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_44),
.B(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_66),
.B2(n_67),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_61),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_56),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_52),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_52),
.B(n_112),
.Y(n_214)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_53),
.B(n_207),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_64),
.Y(n_100)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_56),
.B(n_102),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_60),
.B1(n_70),
.B2(n_71),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_61),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_62),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_68),
.B(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_72),
.B(n_76),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_74),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_78),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_76),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_78),
.B(n_97),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_79),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_85),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_81),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_80),
.A2(n_81),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_81),
.B(n_178),
.Y(n_186)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_84),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_84),
.B(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_86),
.B(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_96),
.C(n_98),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_87),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_88),
.B(n_92),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_91),
.B(n_133),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_91),
.B(n_157),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_93),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_96),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_97),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_100),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_114),
.B2(n_115),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_118),
.B(n_121),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_117),
.B(n_138),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_120),
.B(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_249),
.B(n_254),
.Y(n_123)
);

AOI321xp33_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_222),
.A3(n_242),
.B1(n_247),
.B2(n_248),
.C(n_256),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_199),
.B(n_221),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_182),
.B(n_198),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_169),
.B(n_181),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_150),
.B(n_168),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_144),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_144),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_135),
.B1(n_136),
.B2(n_143),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_131),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_141),
.C(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_145),
.A2(n_146),
.B1(n_148),
.B2(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_162),
.B(n_167),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_158),
.B(n_161),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_160),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_165),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_171),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_177),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_176),
.C(n_177),
.Y(n_197)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_197),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_197),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_189),
.B1(n_190),
.B2(n_196),
.Y(n_183)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_186),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_187),
.C(n_189),
.Y(n_200)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_190),
.B(n_204),
.C(n_210),
.Y(n_246)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_192),
.CI(n_193),
.CON(n_190),
.SN(n_190)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_201),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_210),
.B2(n_211),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_208),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_217),
.C(n_219),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_236),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_236),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_231),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_232),
.C(n_235),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.C(n_230),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_227),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_230),
.B(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_240),
.C(n_241),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_237),
.A2(n_238),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_241),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_246),
.Y(n_247)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_251),
.Y(n_254)
);


endmodule