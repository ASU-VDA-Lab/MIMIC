module real_aes_13308_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_884;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_931;
wire n_683;
wire n_904;
wire n_174;
wire n_780;
wire n_570;
wire n_675;
wire n_840;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_917;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_922;
wire n_520;
wire n_482;
wire n_633;
wire n_926;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx2_ASAP7_75t_SL g173 ( .A(n_0), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_1), .Y(n_335) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_2), .A2(n_48), .B(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g181 ( .A(n_2), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_3), .B(n_168), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_4), .B(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_5), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_6), .B(n_200), .Y(n_640) );
AND2x2_ASAP7_75t_L g274 ( .A(n_7), .B(n_191), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_8), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_9), .B(n_222), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_10), .B(n_222), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_11), .B(n_612), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_12), .B(n_154), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_13), .B(n_286), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_14), .B(n_171), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g659 ( .A(n_15), .Y(n_659) );
BUFx3_ASAP7_75t_L g150 ( .A(n_16), .Y(n_150) );
INVx1_ASAP7_75t_L g156 ( .A(n_16), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_17), .B(n_190), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_18), .B(n_262), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_19), .Y(n_637) );
BUFx10_ASAP7_75t_L g924 ( .A(n_20), .Y(n_924) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_21), .B(n_230), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_22), .Y(n_652) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_23), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_24), .B(n_600), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g250 ( .A(n_25), .B(n_248), .C(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_26), .B(n_230), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_27), .B(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_28), .B(n_262), .Y(n_692) );
NAND2xp33_ASAP7_75t_L g603 ( .A(n_29), .B(n_149), .Y(n_603) );
INVx1_ASAP7_75t_L g185 ( .A(n_30), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g650 ( .A1(n_31), .A2(n_264), .B(n_340), .C(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_32), .B(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_33), .B(n_337), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_34), .B(n_168), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_35), .B(n_313), .Y(n_630) );
INVx1_ASAP7_75t_L g112 ( .A(n_36), .Y(n_112) );
AND3x2_ASAP7_75t_L g939 ( .A(n_36), .B(n_921), .C(n_922), .Y(n_939) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_37), .B(n_224), .Y(n_223) );
AO221x1_ASAP7_75t_L g609 ( .A1(n_38), .A2(n_81), .B1(n_148), .B2(n_230), .C(n_312), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_39), .B(n_627), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_40), .B(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g184 ( .A(n_41), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_42), .B(n_190), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_43), .B(n_163), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g925 ( .A1(n_44), .A2(n_926), .B1(n_933), .B2(n_934), .Y(n_925) );
NAND3xp33_ASAP7_75t_L g695 ( .A(n_45), .B(n_339), .C(n_340), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_46), .B(n_190), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_47), .Y(n_127) );
INVx1_ASAP7_75t_L g180 ( .A(n_48), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_49), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g166 ( .A1(n_50), .A2(n_167), .B(n_170), .C(n_174), .Y(n_166) );
INVx1_ASAP7_75t_L g165 ( .A(n_51), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g656 ( .A(n_52), .Y(n_656) );
A2O1A1Ixp33_ASAP7_75t_L g663 ( .A1(n_53), .A2(n_664), .B(n_665), .C(n_667), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_54), .B(n_190), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g129 ( .A1(n_55), .A2(n_130), .B1(n_131), .B2(n_917), .Y(n_129) );
INVx1_ASAP7_75t_L g917 ( .A(n_55), .Y(n_917) );
INVx1_ASAP7_75t_L g941 ( .A(n_56), .Y(n_941) );
INVx2_ASAP7_75t_L g666 ( .A(n_57), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_58), .B(n_163), .Y(n_642) );
AND2x4_ASAP7_75t_L g109 ( .A(n_59), .B(n_110), .Y(n_109) );
INVx3_ASAP7_75t_L g296 ( .A(n_60), .Y(n_296) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_61), .Y(n_116) );
NOR2xp67_ASAP7_75t_L g126 ( .A(n_61), .B(n_73), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_62), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g110 ( .A(n_63), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_64), .B(n_196), .Y(n_205) );
INVx1_ASAP7_75t_L g311 ( .A(n_65), .Y(n_311) );
AND2x2_ASAP7_75t_L g632 ( .A(n_66), .B(n_163), .Y(n_632) );
INVx1_ASAP7_75t_L g615 ( .A(n_67), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_68), .B(n_108), .C(n_111), .Y(n_107) );
INVx2_ASAP7_75t_L g124 ( .A(n_68), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_69), .B(n_243), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_70), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_71), .B(n_251), .Y(n_332) );
OAI22xp33_ASAP7_75t_L g611 ( .A1(n_72), .A2(n_75), .B1(n_600), .B2(n_612), .Y(n_611) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_73), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_74), .B(n_340), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_76), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g151 ( .A(n_77), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_78), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_79), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_80), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g673 ( .A(n_82), .B(n_191), .Y(n_673) );
INVx1_ASAP7_75t_L g160 ( .A(n_83), .Y(n_160) );
INVx1_ASAP7_75t_L g176 ( .A(n_83), .Y(n_176) );
BUFx3_ASAP7_75t_L g286 ( .A(n_83), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_84), .B(n_243), .Y(n_333) );
INVx1_ASAP7_75t_L g294 ( .A(n_85), .Y(n_294) );
XNOR2xp5_ASAP7_75t_L g930 ( .A(n_86), .B(n_931), .Y(n_930) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_87), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_88), .B(n_178), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_89), .B(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_90), .B(n_191), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_91), .B(n_627), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_92), .B(n_163), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_93), .B(n_203), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_94), .Y(n_289) );
INVx1_ASAP7_75t_L g284 ( .A(n_95), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g697 ( .A(n_96), .Y(n_697) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_97), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_98), .B(n_196), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_117), .B(n_940), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
CKINVDCx14_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
NOR2xp33_ASAP7_75t_L g940 ( .A(n_102), .B(n_941), .Y(n_940) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx2_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
NAND2x1p5_ASAP7_75t_L g104 ( .A(n_105), .B(n_113), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g134 ( .A(n_111), .Y(n_134) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_112), .B(n_126), .Y(n_125) );
INVxp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
OR2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_128), .Y(n_117) );
INVxp67_ASAP7_75t_L g932 ( .A(n_118), .Y(n_932) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_127), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVxp67_ASAP7_75t_L g929 ( .A(n_121), .Y(n_929) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NOR2x1p5_ASAP7_75t_L g122 ( .A(n_123), .B(n_125), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx2_ASAP7_75t_L g922 ( .A(n_124), .Y(n_922) );
HB1xp67_ASAP7_75t_L g921 ( .A(n_126), .Y(n_921) );
OAI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_918), .B(n_925), .Y(n_128) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AO21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_135), .B(n_570), .Y(n_131) );
AOI31xp33_ASAP7_75t_L g570 ( .A1(n_132), .A2(n_571), .A3(n_805), .B(n_880), .Y(n_570) );
INVxp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_SL g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g931 ( .A(n_136), .Y(n_931) );
AND3x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_474), .C(n_520), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_418), .Y(n_137) );
NAND3xp33_ASAP7_75t_SL g138 ( .A(n_139), .B(n_355), .C(n_390), .Y(n_138) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_213), .B1(n_342), .B2(n_349), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_186), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g470 ( .A(n_143), .B(n_216), .Y(n_470) );
AND2x4_ASAP7_75t_L g483 ( .A(n_143), .B(n_378), .Y(n_483) );
AND2x2_ASAP7_75t_L g514 ( .A(n_143), .B(n_399), .Y(n_514) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_143), .Y(n_547) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OR2x6_ASAP7_75t_L g367 ( .A(n_144), .B(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_SL g379 ( .A(n_144), .B(n_346), .Y(n_379) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g345 ( .A(n_145), .Y(n_345) );
OAI21x1_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_161), .B(n_177), .Y(n_145) );
AOI21x1_ASAP7_75t_SL g146 ( .A1(n_147), .A2(n_152), .B(n_157), .Y(n_146) );
OR2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_151), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g222 ( .A(n_149), .Y(n_222) );
INVx2_ASAP7_75t_L g243 ( .A(n_149), .Y(n_243) );
INVx3_ASAP7_75t_L g262 ( .A(n_149), .Y(n_262) );
INVx2_ASAP7_75t_L g268 ( .A(n_149), .Y(n_268) );
INVx2_ASAP7_75t_L g337 ( .A(n_149), .Y(n_337) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_150), .Y(n_172) );
INVx2_ASAP7_75t_L g252 ( .A(n_150), .Y(n_252) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g224 ( .A(n_154), .Y(n_224) );
INVx2_ASAP7_75t_L g227 ( .A(n_154), .Y(n_227) );
INVx2_ASAP7_75t_L g245 ( .A(n_154), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_154), .B(n_659), .Y(n_658) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_155), .Y(n_230) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_156), .Y(n_169) );
AOI22x1_ASAP7_75t_L g259 ( .A1(n_157), .A2(n_175), .B1(n_260), .B2(n_266), .Y(n_259) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_158), .A2(n_195), .B(n_198), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_158), .B(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g291 ( .A(n_159), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_159), .A2(n_598), .B(n_599), .Y(n_597) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx3_ASAP7_75t_L g207 ( .A(n_160), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_166), .Y(n_161) );
OAI21xp33_ASAP7_75t_L g177 ( .A1(n_162), .A2(n_178), .B(n_183), .Y(n_177) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_163), .Y(n_209) );
INVx1_ASAP7_75t_L g348 ( .A(n_163), .Y(n_348) );
INVxp67_ASAP7_75t_SL g583 ( .A(n_163), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_163), .B(n_287), .Y(n_593) );
INVx2_ASAP7_75t_L g622 ( .A(n_163), .Y(n_622) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g192 ( .A(n_164), .Y(n_192) );
BUFx2_ASAP7_75t_L g304 ( .A(n_164), .Y(n_304) );
INVx1_ASAP7_75t_L g182 ( .A(n_165), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_167), .A2(n_267), .B1(n_269), .B2(n_270), .Y(n_266) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g200 ( .A(n_169), .Y(n_200) );
INVx1_ASAP7_75t_L g204 ( .A(n_169), .Y(n_204) );
INVx2_ASAP7_75t_L g339 ( .A(n_169), .Y(n_339) );
INVx1_ASAP7_75t_L g657 ( .A(n_169), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_171), .B(n_173), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g197 ( .A(n_172), .Y(n_197) );
INVx1_ASAP7_75t_L g317 ( .A(n_172), .Y(n_317) );
INVx2_ASAP7_75t_L g612 ( .A(n_172), .Y(n_612) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AOI21x1_ASAP7_75t_L g241 ( .A1(n_175), .A2(n_242), .B(n_244), .Y(n_241) );
AOI21xp5_ASAP7_75t_SL g623 ( .A1(n_175), .A2(n_624), .B(n_625), .Y(n_623) );
BUFx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g232 ( .A(n_176), .Y(n_232) );
INVxp67_ASAP7_75t_L g271 ( .A(n_178), .Y(n_271) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_179), .B(n_211), .Y(n_648) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_182), .Y(n_179) );
AOI21x1_ASAP7_75t_L g280 ( .A1(n_180), .A2(n_181), .B(n_182), .Y(n_280) );
INVx1_ASAP7_75t_L g273 ( .A(n_183), .Y(n_273) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g212 ( .A(n_184), .Y(n_212) );
BUFx6f_ASAP7_75t_SL g233 ( .A(n_184), .Y(n_233) );
INVx3_ASAP7_75t_L g287 ( .A(n_184), .Y(n_287) );
OR2x2_ASAP7_75t_L g459 ( .A(n_186), .B(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g480 ( .A(n_186), .B(n_367), .Y(n_480) );
BUFx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g387 ( .A(n_187), .Y(n_387) );
AND2x2_ASAP7_75t_L g394 ( .A(n_187), .B(n_346), .Y(n_394) );
INVx2_ASAP7_75t_L g399 ( .A(n_187), .Y(n_399) );
AND2x2_ASAP7_75t_L g414 ( .A(n_187), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g424 ( .A(n_187), .B(n_236), .Y(n_424) );
OR2x2_ASAP7_75t_L g440 ( .A(n_187), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g469 ( .A(n_187), .Y(n_469) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2x1_ASAP7_75t_L g188 ( .A(n_189), .B(n_193), .Y(n_188) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_190), .Y(n_239) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
OAI21x1_ASAP7_75t_SL g193 ( .A1(n_194), .A2(n_201), .B(n_208), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_196), .A2(n_293), .B1(n_295), .B2(n_297), .Y(n_292) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_197), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_205), .B(n_206), .Y(n_201) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_207), .A2(n_221), .B(n_223), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_207), .A2(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g667 ( .A(n_207), .Y(n_667) );
NOR2x1_ASAP7_75t_SL g208 ( .A(n_209), .B(n_210), .Y(n_208) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_209), .Y(n_218) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_SL g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g253 ( .A(n_212), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_255), .B1(n_319), .B2(n_323), .Y(n_213) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
OR2x2_ASAP7_75t_L g507 ( .A(n_215), .B(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_235), .Y(n_215) );
BUFx3_ASAP7_75t_L g321 ( .A(n_216), .Y(n_321) );
AND2x2_ASAP7_75t_L g412 ( .A(n_216), .B(n_387), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_216), .Y(n_415) );
AND2x2_ASAP7_75t_L g529 ( .A(n_216), .B(n_345), .Y(n_529) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_217), .Y(n_451) );
OAI21x1_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_234), .Y(n_217) );
OAI21x1_ASAP7_75t_L g352 ( .A1(n_218), .A2(n_259), .B(n_353), .Y(n_352) );
OAI21x1_ASAP7_75t_L g378 ( .A1(n_218), .A2(n_219), .B(n_234), .Y(n_378) );
OAI21x1_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_225), .B(n_233), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_228), .B(n_231), .Y(n_225) );
INVx2_ASAP7_75t_L g264 ( .A(n_227), .Y(n_264) );
INVxp67_ASAP7_75t_L g249 ( .A(n_229), .Y(n_249) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_230), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g297 ( .A(n_230), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_231), .A2(n_315), .B(n_316), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_231), .A2(n_332), .B(n_333), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_231), .A2(n_630), .B(n_631), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_231), .A2(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g672 ( .A(n_231), .Y(n_672) );
BUFx10_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g248 ( .A(n_232), .Y(n_248) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_233), .A2(n_306), .B(n_314), .Y(n_305) );
OAI21x1_ASAP7_75t_L g635 ( .A1(n_233), .A2(n_636), .B(n_639), .Y(n_635) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_235), .Y(n_427) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_236), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_236), .B(n_345), .Y(n_460) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g368 ( .A(n_237), .Y(n_368) );
INVxp67_ASAP7_75t_SL g441 ( .A(n_237), .Y(n_441) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OAI21x1_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_254), .Y(n_238) );
OA21x2_ASAP7_75t_L g346 ( .A1(n_240), .A2(n_254), .B(n_347), .Y(n_346) );
OAI21x1_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_246), .B(n_253), .Y(n_240) );
O2A1O1Ixp5_ASAP7_75t_L g636 ( .A1(n_245), .A2(n_592), .B(n_637), .C(n_638), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_249), .B(n_250), .Y(n_246) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g313 ( .A(n_252), .Y(n_313) );
INVx2_ASAP7_75t_L g600 ( .A(n_252), .Y(n_600) );
INVx2_ASAP7_75t_L g627 ( .A(n_252), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g330 ( .A1(n_253), .A2(n_331), .B(n_334), .Y(n_330) );
INVx2_ASAP7_75t_L g420 ( .A(n_255), .Y(n_420) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_275), .Y(n_255) );
INVx1_ASAP7_75t_L g385 ( .A(n_256), .Y(n_385) );
INVx1_ASAP7_75t_L g417 ( .A(n_256), .Y(n_417) );
BUFx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g403 ( .A(n_257), .Y(n_403) );
AO31x2_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_271), .A3(n_272), .B(n_274), .Y(n_257) );
AO31x2_ASAP7_75t_L g435 ( .A1(n_258), .A2(n_271), .A3(n_272), .B(n_274), .Y(n_435) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OAI22x1_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_263), .B1(n_264), .B2(n_265), .Y(n_260) );
INVxp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVxp67_ASAP7_75t_L g307 ( .A(n_268), .Y(n_307) );
BUFx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g353 ( .A(n_274), .Y(n_353) );
INVx1_ASAP7_75t_L g553 ( .A(n_275), .Y(n_553) );
INVxp67_ASAP7_75t_SL g564 ( .A(n_275), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_300), .Y(n_275) );
NOR2x1_ASAP7_75t_L g326 ( .A(n_276), .B(n_327), .Y(n_326) );
BUFx2_ASAP7_75t_L g389 ( .A(n_276), .Y(n_389) );
INVx1_ASAP7_75t_L g431 ( .A(n_276), .Y(n_431) );
AND2x2_ASAP7_75t_L g490 ( .A(n_276), .B(n_301), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_276), .B(n_354), .Y(n_512) );
INVx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g350 ( .A(n_277), .B(n_301), .Y(n_350) );
AO21x2_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_281), .B(n_298), .Y(n_277) );
AO21x1_ASAP7_75t_L g363 ( .A1(n_278), .A2(n_281), .B(n_298), .Y(n_363) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NOR2xp33_ASAP7_75t_SL g298 ( .A(n_279), .B(n_299), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_279), .B(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_R g613 ( .A(n_280), .B(n_287), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_292), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_285), .B1(n_288), .B2(n_290), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
NOR3xp33_ASAP7_75t_L g293 ( .A(n_286), .B(n_287), .C(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g312 ( .A(n_286), .Y(n_312) );
INVx2_ASAP7_75t_L g340 ( .A(n_286), .Y(n_340) );
INVx1_ASAP7_75t_L g592 ( .A(n_286), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_287), .B(n_291), .Y(n_290) );
NOR3xp33_ASAP7_75t_L g295 ( .A(n_287), .B(n_291), .C(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g604 ( .A(n_287), .Y(n_604) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_301), .Y(n_325) );
INVx3_ASAP7_75t_L g359 ( .A(n_301), .Y(n_359) );
INVx2_ASAP7_75t_L g372 ( .A(n_301), .Y(n_372) );
AND2x2_ASAP7_75t_L g376 ( .A(n_301), .B(n_352), .Y(n_376) );
INVx1_ASAP7_75t_L g400 ( .A(n_301), .Y(n_400) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI21x1_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_305), .B(n_318), .Y(n_302) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_303), .A2(n_330), .B(n_341), .Y(n_329) );
OAI21x1_ASAP7_75t_L g634 ( .A1(n_303), .A2(n_635), .B(n_642), .Y(n_634) );
BUFx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVxp67_ASAP7_75t_L g675 ( .A(n_304), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .B(n_309), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_L g588 ( .A(n_312), .Y(n_588) );
INVxp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_321), .B(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g438 ( .A(n_321), .Y(n_438) );
OR2x2_ASAP7_75t_L g479 ( .A(n_321), .B(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
OR2x2_ASAP7_75t_L g559 ( .A(n_324), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g375 ( .A(n_327), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_327), .B(n_359), .Y(n_408) );
NOR2xp67_ASAP7_75t_L g518 ( .A(n_327), .B(n_358), .Y(n_518) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx3_ASAP7_75t_L g354 ( .A(n_328), .Y(n_354) );
AND2x2_ASAP7_75t_L g361 ( .A(n_328), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g473 ( .A(n_328), .B(n_352), .Y(n_473) );
INVx1_ASAP7_75t_L g496 ( .A(n_328), .Y(n_496) );
INVx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
O2A1O1Ixp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B(n_338), .C(n_340), .Y(n_334) );
OAI21xp5_ASAP7_75t_L g693 ( .A1(n_336), .A2(n_694), .B(n_695), .Y(n_693) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AOI211xp5_ASAP7_75t_L g355 ( .A1(n_344), .A2(n_356), .B(n_364), .C(n_380), .Y(n_355) );
AND2x2_ASAP7_75t_L g504 ( .A(n_344), .B(n_468), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_344), .B(n_399), .Y(n_557) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_L g383 ( .A(n_345), .Y(n_383) );
AND2x4_ASAP7_75t_L g393 ( .A(n_345), .B(n_378), .Y(n_393) );
OA21x2_ASAP7_75t_L g595 ( .A1(n_347), .A2(n_596), .B(n_605), .Y(n_595) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
AOI32xp33_ASAP7_75t_L g481 ( .A1(n_349), .A2(n_423), .A3(n_482), .B1(n_484), .B2(n_486), .Y(n_481) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
AND2x2_ASAP7_75t_L g472 ( .A(n_350), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g373 ( .A(n_351), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_351), .B(n_431), .Y(n_447) );
AND2x2_ASAP7_75t_L g500 ( .A(n_351), .B(n_389), .Y(n_500) );
AND2x2_ASAP7_75t_L g563 ( .A(n_351), .B(n_564), .Y(n_563) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g410 ( .A(n_352), .Y(n_410) );
OR2x2_ASAP7_75t_L g434 ( .A(n_354), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
AOI21xp33_ASAP7_75t_SL g453 ( .A1(n_357), .A2(n_411), .B(n_452), .Y(n_453) );
OR2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
BUFx2_ASAP7_75t_L g498 ( .A(n_358), .Y(n_498) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_359), .B(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g463 ( .A(n_359), .B(n_435), .Y(n_463) );
INVx1_ASAP7_75t_L g397 ( .A(n_360), .Y(n_397) );
OR2x2_ASAP7_75t_L g443 ( .A(n_360), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g402 ( .A(n_361), .Y(n_402) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_361), .Y(n_464) );
AND2x2_ASAP7_75t_L g505 ( .A(n_361), .B(n_403), .Y(n_505) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g371 ( .A(n_363), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_363), .B(n_410), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_369), .B1(n_374), .B2(n_377), .Y(n_364) );
INVxp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2x1p5_ASAP7_75t_L g413 ( .A(n_366), .B(n_414), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_366), .A2(n_536), .B1(n_538), .B2(n_540), .Y(n_535) );
INVx2_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g456 ( .A(n_367), .B(n_399), .Y(n_456) );
AND2x2_ASAP7_75t_L g384 ( .A(n_368), .B(n_378), .Y(n_384) );
INVx2_ASAP7_75t_L g569 ( .A(n_369), .Y(n_569) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_373), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g477 ( .A(n_371), .B(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g486 ( .A(n_371), .B(n_473), .Y(n_486) );
AND2x2_ASAP7_75t_L g525 ( .A(n_371), .B(n_417), .Y(n_525) );
AND2x2_ASAP7_75t_L g544 ( .A(n_371), .B(n_508), .Y(n_544) );
INVx1_ASAP7_75t_L g391 ( .A(n_373), .Y(n_391) );
OAI321xp33_ASAP7_75t_L g561 ( .A1(n_374), .A2(n_450), .A3(n_484), .B1(n_562), .B2(n_565), .C(n_568), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_375), .B(n_376), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_375), .B(n_517), .Y(n_560) );
INVx1_ASAP7_75t_L g444 ( .A(n_376), .Y(n_444) );
AND2x4_ASAP7_75t_L g510 ( .A(n_376), .B(n_511), .Y(n_510) );
INVx3_ASAP7_75t_L g531 ( .A(n_377), .Y(n_531) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
AND2x4_ASAP7_75t_L g423 ( .A(n_378), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g405 ( .A(n_379), .Y(n_405) );
NOR4xp25_ASAP7_75t_L g380 ( .A(n_381), .B(n_385), .C(n_386), .D(n_388), .Y(n_380) );
NAND2x1_ASAP7_75t_L g421 ( .A(n_381), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_382), .A2(n_457), .B1(n_504), .B2(n_505), .Y(n_503) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
OAI322xp33_ASAP7_75t_L g542 ( .A1(n_385), .A2(n_543), .A3(n_545), .B1(n_551), .B2(n_554), .C1(n_555), .C2(n_559), .Y(n_542) );
AND2x2_ASAP7_75t_L g502 ( .A(n_386), .B(n_470), .Y(n_502) );
BUFx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g485 ( .A(n_387), .B(n_441), .Y(n_485) );
INVx1_ASAP7_75t_L g508 ( .A(n_387), .Y(n_508) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_389), .B(n_434), .Y(n_457) );
AOI211xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B(n_395), .C(n_406), .Y(n_390) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g466 ( .A(n_393), .Y(n_466) );
NOR2x1_ASAP7_75t_L g566 ( .A(n_393), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g452 ( .A(n_394), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_398), .B(n_401), .C(n_404), .Y(n_395) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
AND2x2_ASAP7_75t_L g558 ( .A(n_399), .B(n_529), .Y(n_558) );
INVx2_ASAP7_75t_L g433 ( .A(n_400), .Y(n_433) );
OR2x6_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx2_ASAP7_75t_L g478 ( .A(n_403), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_403), .B(n_490), .Y(n_489) );
NAND2xp33_ASAP7_75t_SL g540 ( .A(n_404), .B(n_541), .Y(n_540) );
INVx2_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
OAI32xp33_ASAP7_75t_L g406 ( .A1(n_405), .A2(n_407), .A3(n_411), .B1(n_413), .B2(n_416), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_405), .B(n_508), .Y(n_554) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx2_ASAP7_75t_L g517 ( .A(n_409), .Y(n_517) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g488 ( .A(n_415), .B(n_460), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g418 ( .A(n_419), .B(n_436), .C(n_454), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_425), .B2(n_428), .Y(n_419) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
O2A1O1Ixp5_ASAP7_75t_L g465 ( .A1(n_424), .A2(n_466), .B(n_467), .C(n_471), .Y(n_465) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_424), .Y(n_523) );
INVx1_ASAP7_75t_L g567 ( .A(n_424), .Y(n_567) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g534 ( .A(n_430), .Y(n_534) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g539 ( .A(n_431), .B(n_496), .Y(n_539) );
INVx1_ASAP7_75t_L g446 ( .A(n_432), .Y(n_446) );
NOR2x1p5_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g497 ( .A(n_435), .Y(n_497) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_442), .B1(n_445), .B2(n_448), .C(n_453), .Y(n_436) );
INVx1_ASAP7_75t_L g492 ( .A(n_437), .Y(n_492) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g527 ( .A(n_440), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_442), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g519 ( .A(n_451), .B(n_485), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_457), .B1(n_458), .B2(n_461), .C(n_465), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
AND2x4_ASAP7_75t_L g538 ( .A(n_462), .B(n_539), .Y(n_538) );
INVx2_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g537 ( .A(n_463), .B(n_512), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_470), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx3_ASAP7_75t_R g541 ( .A(n_470), .Y(n_541) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NOR4xp25_ASAP7_75t_L g474 ( .A(n_475), .B(n_487), .C(n_491), .D(n_506), .Y(n_474) );
OAI21xp33_ASAP7_75t_SL g475 ( .A1(n_476), .A2(n_479), .B(n_481), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AOI21xp33_ASAP7_75t_SL g487 ( .A1(n_479), .A2(n_488), .B(n_489), .Y(n_487) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_483), .A2(n_519), .B(n_569), .Y(n_568) );
BUFx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI221xp5_ASAP7_75t_SL g491 ( .A1(n_492), .A2(n_493), .B1(n_499), .B2(n_501), .C(n_503), .Y(n_491) );
OAI221xp5_ASAP7_75t_L g506 ( .A1(n_493), .A2(n_507), .B1(n_509), .B2(n_513), .C(n_515), .Y(n_506) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_498), .Y(n_494) );
INVx1_ASAP7_75t_L g533 ( .A(n_495), .Y(n_533) );
AND2x4_ASAP7_75t_L g552 ( .A(n_495), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g549 ( .A(n_496), .Y(n_549) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVxp67_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND4xp25_ASAP7_75t_L g530 ( .A(n_508), .B(n_531), .C(n_532), .D(n_534), .Y(n_530) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVxp67_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_519), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
NOR3xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_542), .C(n_561), .Y(n_520) );
NAND4xp25_ASAP7_75t_L g521 ( .A(n_522), .B(n_524), .C(n_530), .D(n_535), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_529), .Y(n_550) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NOR2xp33_ASAP7_75t_SL g545 ( .A(n_546), .B(n_550), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NOR2x1_ASAP7_75t_L g571 ( .A(n_572), .B(n_752), .Y(n_571) );
NAND3xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_722), .C(n_742), .Y(n_572) );
AOI221xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_616), .B1(n_676), .B2(n_685), .C(n_700), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_606), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_594), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g775 ( .A(n_578), .Y(n_775) );
AND2x2_ASAP7_75t_L g829 ( .A(n_578), .B(n_821), .Y(n_829) );
AND2x2_ASAP7_75t_L g910 ( .A(n_578), .B(n_608), .Y(n_910) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_579), .B(n_687), .Y(n_718) );
AND2x2_ASAP7_75t_L g852 ( .A(n_579), .B(n_608), .Y(n_852) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g699 ( .A(n_580), .B(n_595), .Y(n_699) );
AND2x2_ASAP7_75t_L g703 ( .A(n_580), .B(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g731 ( .A(n_580), .B(n_608), .Y(n_731) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_580), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_580), .B(n_595), .Y(n_786) );
AND2x4_ASAP7_75t_L g580 ( .A(n_581), .B(n_584), .Y(n_580) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OAI21xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_589), .B(n_593), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B(n_588), .Y(n_585) );
OAI21xp5_ASAP7_75t_L g654 ( .A1(n_588), .A2(n_655), .B(n_658), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B(n_592), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_592), .A2(n_691), .B(n_692), .Y(n_690) );
OR2x2_ASAP7_75t_L g751 ( .A(n_594), .B(n_706), .Y(n_751) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g704 ( .A(n_595), .Y(n_704) );
INVx1_ASAP7_75t_L g716 ( .A(n_595), .Y(n_716) );
INVx1_ASAP7_75t_L g741 ( .A(n_595), .Y(n_741) );
AND2x2_ASAP7_75t_L g799 ( .A(n_595), .B(n_688), .Y(n_799) );
OAI21xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_601), .B(n_604), .Y(n_596) );
AND2x4_ASAP7_75t_L g621 ( .A(n_604), .B(n_622), .Y(n_621) );
AOI21xp33_ASAP7_75t_L g674 ( .A1(n_604), .A2(n_673), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g760 ( .A(n_606), .Y(n_760) );
OR2x2_ASAP7_75t_L g789 ( .A(n_606), .B(n_751), .Y(n_789) );
OR2x2_ASAP7_75t_L g808 ( .A(n_606), .B(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g770 ( .A(n_607), .Y(n_770) );
AND2x2_ASAP7_75t_L g817 ( .A(n_607), .B(n_708), .Y(n_817) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_607), .Y(n_887) );
BUFx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g686 ( .A(n_608), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g705 ( .A(n_608), .B(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g773 ( .A(n_608), .B(n_704), .Y(n_773) );
INVx2_ASAP7_75t_SL g821 ( .A(n_608), .Y(n_821) );
AO31x2_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .A3(n_613), .B(n_614), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_612), .B(n_652), .Y(n_651) );
INVxp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_643), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_618), .B(n_757), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_618), .A2(n_792), .B1(n_799), .B2(n_800), .Y(n_798) );
AND2x2_ASAP7_75t_L g883 ( .A(n_618), .B(n_884), .Y(n_883) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_633), .Y(n_618) );
INVx2_ASAP7_75t_L g680 ( .A(n_619), .Y(n_680) );
INVx1_ASAP7_75t_L g735 ( .A(n_619), .Y(n_735) );
OR2x2_ASAP7_75t_L g746 ( .A(n_619), .B(n_662), .Y(n_746) );
AND2x2_ASAP7_75t_L g841 ( .A(n_619), .B(n_634), .Y(n_841) );
NAND2x1p5_ASAP7_75t_L g619 ( .A(n_620), .B(n_628), .Y(n_619) );
NAND2x1_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
AOI21x1_ASAP7_75t_L g628 ( .A1(n_621), .A2(n_629), .B(n_632), .Y(n_628) );
O2A1O1Ixp5_ASAP7_75t_L g689 ( .A1(n_621), .A2(n_690), .B(n_693), .C(n_696), .Y(n_689) );
INVx2_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g712 ( .A(n_633), .Y(n_712) );
INVx1_ASAP7_75t_L g726 ( .A(n_633), .Y(n_726) );
INVx1_ASAP7_75t_L g736 ( .A(n_633), .Y(n_736) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVxp33_ASAP7_75t_L g824 ( .A(n_634), .Y(n_824) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_643), .Y(n_754) );
INVx1_ASAP7_75t_L g853 ( .A(n_643), .Y(n_853) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_645), .B(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g867 ( .A(n_645), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_661), .Y(n_645) );
INVx3_ASAP7_75t_L g684 ( .A(n_646), .Y(n_684) );
AND2x2_ASAP7_75t_L g766 ( .A(n_646), .B(n_712), .Y(n_766) );
AO21x2_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B(n_653), .Y(n_646) );
AO21x1_ASAP7_75t_SL g709 ( .A1(n_647), .A2(n_649), .B(n_653), .Y(n_709) );
INVxp67_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
OAI21x1_ASAP7_75t_SL g653 ( .A1(n_648), .A2(n_654), .B(n_660), .Y(n_653) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g664 ( .A(n_657), .Y(n_664) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g681 ( .A(n_662), .Y(n_681) );
INVx2_ASAP7_75t_L g711 ( .A(n_662), .Y(n_711) );
AND2x2_ASAP7_75t_L g721 ( .A(n_662), .B(n_680), .Y(n_721) );
AND2x2_ASAP7_75t_L g757 ( .A(n_662), .B(n_684), .Y(n_757) );
AND2x2_ASAP7_75t_L g837 ( .A(n_662), .B(n_679), .Y(n_837) );
AO21x2_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_668), .B(n_674), .Y(n_662) );
NOR2xp67_ASAP7_75t_L g665 ( .A(n_664), .B(n_666), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_672), .B(n_673), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_675), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_682), .Y(n_677) );
OR2x2_ASAP7_75t_L g905 ( .A(n_678), .B(n_726), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
OR2x2_ASAP7_75t_L g783 ( .A(n_679), .B(n_712), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_679), .B(n_683), .Y(n_914) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g790 ( .A(n_682), .Y(n_790) );
BUFx2_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g728 ( .A(n_683), .Y(n_728) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g823 ( .A(n_684), .B(n_824), .Y(n_823) );
AND2x2_ASAP7_75t_L g830 ( .A(n_684), .B(n_711), .Y(n_830) );
OR2x2_ASAP7_75t_L g846 ( .A(n_684), .B(n_711), .Y(n_846) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_698), .Y(n_685) );
AND2x4_ASAP7_75t_L g785 ( .A(n_686), .B(n_786), .Y(n_785) );
AND2x4_ASAP7_75t_L g804 ( .A(n_686), .B(n_703), .Y(n_804) );
INVx2_ASAP7_75t_L g706 ( .A(n_687), .Y(n_706) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g730 ( .A(n_688), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_688), .B(n_741), .Y(n_740) );
BUFx2_ASAP7_75t_SL g762 ( .A(n_688), .Y(n_762) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g818 ( .A(n_698), .Y(n_818) );
BUFx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g761 ( .A(n_699), .B(n_762), .Y(n_761) );
AND2x4_ASAP7_75t_SL g835 ( .A(n_699), .B(n_821), .Y(n_835) );
AND2x2_ASAP7_75t_L g896 ( .A(n_699), .B(n_730), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_707), .B1(n_713), .B2(n_719), .Y(n_700) );
INVx3_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x4_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
NAND3xp33_ASAP7_75t_L g875 ( .A(n_706), .B(n_876), .C(n_877), .Y(n_875) );
INVx1_ASAP7_75t_L g909 ( .A(n_706), .Y(n_909) );
OR2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .Y(n_707) );
AND2x2_ASAP7_75t_L g720 ( .A(n_708), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g743 ( .A(n_708), .B(n_744), .Y(n_743) );
AND2x4_ASAP7_75t_SL g802 ( .A(n_708), .B(n_794), .Y(n_802) );
INVx5_ASAP7_75t_L g856 ( .A(n_708), .Y(n_856) );
AND2x4_ASAP7_75t_L g895 ( .A(n_708), .B(n_837), .Y(n_895) );
AND2x2_ASAP7_75t_L g899 ( .A(n_708), .B(n_782), .Y(n_899) );
BUFx6f_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_L g884 ( .A(n_709), .Y(n_884) );
NOR2x1_ASAP7_75t_L g913 ( .A(n_710), .B(n_914), .Y(n_913) );
OR2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g778 ( .A(n_711), .Y(n_778) );
NAND2xp5_ASAP7_75t_SL g874 ( .A(n_713), .B(n_875), .Y(n_874) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AND2x4_ASAP7_75t_L g886 ( .A(n_714), .B(n_887), .Y(n_886) );
AND2x4_ASAP7_75t_L g714 ( .A(n_715), .B(n_717), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_716), .B(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OR2x2_ASAP7_75t_L g819 ( .A(n_718), .B(n_820), .Y(n_819) );
OR2x2_ASAP7_75t_L g861 ( .A(n_718), .B(n_773), .Y(n_861) );
INVx2_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
AND2x4_ASAP7_75t_L g727 ( .A(n_721), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g738 ( .A(n_721), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_721), .B(n_766), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_729), .B(n_732), .Y(n_722) );
OAI21xp5_ASAP7_75t_L g903 ( .A1(n_723), .A2(n_904), .B(n_906), .Y(n_903) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2x1_ASAP7_75t_SL g724 ( .A(n_725), .B(n_727), .Y(n_724) );
BUFx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_726), .B(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_726), .B(n_830), .Y(n_859) );
INVx2_ASAP7_75t_L g868 ( .A(n_726), .Y(n_868) );
AND2x4_ASAP7_75t_SL g873 ( .A(n_726), .B(n_815), .Y(n_873) );
NOR2x1_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_730), .B(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g793 ( .A(n_730), .B(n_794), .Y(n_793) );
INVx2_ASAP7_75t_L g800 ( .A(n_730), .Y(n_800) );
OR2x2_ASAP7_75t_L g739 ( .A(n_731), .B(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g794 ( .A(n_731), .Y(n_794) );
INVx1_ASAP7_75t_L g871 ( .A(n_731), .Y(n_871) );
AOI21xp33_ASAP7_75t_SL g732 ( .A1(n_733), .A2(n_737), .B(n_739), .Y(n_732) );
AOI32xp33_ASAP7_75t_L g862 ( .A1(n_733), .A2(n_830), .A3(n_863), .B1(n_864), .B2(n_869), .Y(n_862) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVx3_ASAP7_75t_L g792 ( .A(n_735), .Y(n_792) );
OR2x2_ASAP7_75t_L g745 ( .A(n_736), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g833 ( .A(n_736), .Y(n_833) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_737), .A2(n_798), .B1(n_801), .B2(n_803), .Y(n_797) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND2xp33_ASAP7_75t_L g860 ( .A(n_739), .B(n_861), .Y(n_860) );
INVx2_ASAP7_75t_L g776 ( .A(n_740), .Y(n_776) );
BUFx2_ASAP7_75t_L g849 ( .A(n_740), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_747), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g806 ( .A1(n_744), .A2(n_778), .B1(n_807), .B2(n_810), .C(n_813), .Y(n_806) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g782 ( .A(n_746), .Y(n_782) );
INVx1_ASAP7_75t_L g815 ( .A(n_746), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_748), .B(n_812), .Y(n_811) );
AND2x2_ASAP7_75t_L g854 ( .A(n_748), .B(n_776), .Y(n_854) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OR2x6_ASAP7_75t_L g900 ( .A(n_751), .B(n_901), .Y(n_900) );
NAND3xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_763), .C(n_787), .Y(n_752) );
OAI21xp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .B(n_758), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OAI22xp33_ASAP7_75t_L g888 ( .A1(n_756), .A2(n_789), .B1(n_889), .B2(n_890), .Y(n_888) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVx2_ASAP7_75t_L g902 ( .A(n_761), .Y(n_902) );
OR2x2_ASAP7_75t_L g772 ( .A(n_762), .B(n_773), .Y(n_772) );
NOR2x1_ASAP7_75t_SL g812 ( .A(n_762), .B(n_773), .Y(n_812) );
AOI221xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_767), .B1(n_771), .B2(n_777), .C(n_779), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g777 ( .A(n_766), .B(n_778), .Y(n_777) );
INVxp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
OR2x2_ASAP7_75t_L g916 ( .A(n_769), .B(n_775), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_774), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx1_ASAP7_75t_L g877 ( .A(n_775), .Y(n_877) );
AND2x2_ASAP7_75t_L g828 ( .A(n_776), .B(n_829), .Y(n_828) );
AND2x2_ASAP7_75t_L g863 ( .A(n_776), .B(n_852), .Y(n_863) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_783), .B(n_784), .Y(n_779) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_780), .A2(n_898), .B1(n_900), .B2(n_902), .Y(n_897) );
BUFx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_781), .B(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g857 ( .A(n_783), .Y(n_857) );
OR2x2_ASAP7_75t_L g889 ( .A(n_783), .B(n_856), .Y(n_889) );
INVx4_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AOI321xp33_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_790), .A3(n_791), .B1(n_793), .B2(n_795), .C(n_797), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx2_ASAP7_75t_SL g809 ( .A(n_799), .Y(n_809) );
AND2x4_ASAP7_75t_L g851 ( .A(n_799), .B(n_852), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_799), .B(n_871), .Y(n_870) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx4_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
AND5x1_ASAP7_75t_L g805 ( .A(n_806), .B(n_825), .C(n_850), .D(n_862), .E(n_872), .Y(n_805) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
OAI22xp33_ASAP7_75t_L g838 ( .A1(n_808), .A2(n_839), .B1(n_842), .B2(n_847), .Y(n_838) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OAI32xp33_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_816), .A3(n_818), .B1(n_819), .B2(n_822), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g893 ( .A(n_823), .Y(n_893) );
NOR2xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_838), .Y(n_825) );
OAI32xp33_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_830), .A3(n_831), .B1(n_834), .B2(n_836), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g901 ( .A(n_829), .Y(n_901) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
A2O1A1Ixp33_ASAP7_75t_L g892 ( .A1(n_834), .A2(n_846), .B(n_893), .C(n_894), .Y(n_892) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVxp33_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_837), .B(n_868), .Y(n_879) );
AND2x2_ASAP7_75t_L g885 ( .A(n_837), .B(n_856), .Y(n_885) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx4_ASAP7_75t_L g844 ( .A(n_841), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_845), .Y(n_842) );
AOI322xp5_ASAP7_75t_L g850 ( .A1(n_843), .A2(n_851), .A3(n_853), .B1(n_854), .B2(n_855), .C1(n_858), .C2(n_860), .Y(n_850) );
INVx6_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVxp67_ASAP7_75t_L g890 ( .A(n_851), .Y(n_890) );
AND2x2_ASAP7_75t_L g855 ( .A(n_856), .B(n_857), .Y(n_855) );
INVx1_ASAP7_75t_L g876 ( .A(n_856), .Y(n_876) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_863), .A2(n_873), .B1(n_874), .B2(n_878), .Y(n_872) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g912 ( .A(n_865), .Y(n_912) );
OR2x2_ASAP7_75t_L g865 ( .A(n_866), .B(n_868), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
OAI31xp33_ASAP7_75t_L g911 ( .A1(n_873), .A2(n_912), .A3(n_913), .B(n_915), .Y(n_911) );
INVx2_ASAP7_75t_SL g878 ( .A(n_879), .Y(n_878) );
AND4x1_ASAP7_75t_L g880 ( .A(n_881), .B(n_891), .C(n_903), .D(n_911), .Y(n_880) );
O2A1O1Ixp33_ASAP7_75t_SL g881 ( .A1(n_882), .A2(n_885), .B(n_886), .C(n_888), .Y(n_881) );
HB1xp67_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
NOR2xp33_ASAP7_75t_SL g891 ( .A(n_892), .B(n_897), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_895), .B(n_896), .Y(n_894) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_909), .B(n_910), .Y(n_908) );
INVx2_ASAP7_75t_SL g915 ( .A(n_916), .Y(n_915) );
BUFx4f_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
OR2x6_ASAP7_75t_L g919 ( .A(n_920), .B(n_923), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_921), .B(n_922), .Y(n_920) );
INVx3_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx2_ASAP7_75t_L g933 ( .A(n_924), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_924), .B(n_939), .Y(n_938) );
OAI21xp5_ASAP7_75t_L g926 ( .A1(n_927), .A2(n_930), .B(n_932), .Y(n_926) );
CKINVDCx5p33_ASAP7_75t_R g927 ( .A(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
BUFx3_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
BUFx3_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
BUFx3_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
endmodule