module fake_jpeg_1346_n_149 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_149);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_53),
.Y(n_69)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_37),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_67),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_42),
.B1(n_50),
.B2(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_68),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_52),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_48),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_79),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_43),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_46),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_72),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_51),
.B(n_40),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_81),
.A2(n_41),
.B(n_55),
.Y(n_90)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_55),
.Y(n_96)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_70),
.B1(n_59),
.B2(n_36),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_0),
.B(n_2),
.C(n_4),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_95),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_60),
.B1(n_54),
.B2(n_50),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_97),
.B(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_101),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_42),
.B1(n_44),
.B2(n_3),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_74),
.C(n_78),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_112),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_33),
.Y(n_103)
);

NOR3xp33_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_107),
.C(n_22),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_105),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_109),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_15),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_99),
.B(n_0),
.Y(n_109)
);

NAND2x1_ASAP7_75t_SL g111 ( 
.A(n_89),
.B(n_2),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_6),
.B(n_7),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_16),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_117),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_4),
.B(n_5),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_6),
.B(n_8),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_20),
.C(n_32),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_87),
.B(n_14),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_5),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_120),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_122),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_23),
.B(n_31),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_127),
.B1(n_129),
.B2(n_10),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_24),
.B(n_29),
.Y(n_129)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_105),
.A3(n_117),
.B1(n_112),
.B2(n_8),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_124),
.B1(n_126),
.B2(n_130),
.Y(n_140)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_133),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_134),
.B(n_136),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_142),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_138),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_132),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_128),
.C(n_131),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_105),
.B(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_13),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_28),
.Y(n_149)
);


endmodule