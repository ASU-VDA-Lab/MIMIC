module fake_aes_7096_n_668 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_668);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_668;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_384;
wire n_434;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_575;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_69), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_31), .Y(n_78) );
INVxp67_ASAP7_75t_SL g79 ( .A(n_50), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_42), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_43), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_53), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_18), .Y(n_83) );
CKINVDCx14_ASAP7_75t_R g84 ( .A(n_25), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_8), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_59), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_41), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_30), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_35), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_44), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_12), .Y(n_91) );
INVxp33_ASAP7_75t_L g92 ( .A(n_16), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_9), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_23), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_12), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_55), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_40), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_67), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_51), .Y(n_99) );
BUFx3_ASAP7_75t_L g100 ( .A(n_60), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_1), .Y(n_101) );
BUFx2_ASAP7_75t_L g102 ( .A(n_15), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_73), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_70), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_7), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_68), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_15), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_56), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_72), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_8), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_61), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_62), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_48), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_58), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_5), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_20), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_9), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_46), .Y(n_118) );
INVx3_ASAP7_75t_L g119 ( .A(n_24), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_49), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_39), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_65), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_22), .Y(n_123) );
AND2x6_ASAP7_75t_L g124 ( .A(n_119), .B(n_29), .Y(n_124) );
BUFx3_ASAP7_75t_L g125 ( .A(n_119), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_95), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_95), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_119), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_77), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_114), .B(n_0), .Y(n_130) );
AND2x6_ASAP7_75t_L g131 ( .A(n_100), .B(n_32), .Y(n_131) );
BUFx8_ASAP7_75t_L g132 ( .A(n_114), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_77), .Y(n_133) );
INVx4_ASAP7_75t_L g134 ( .A(n_100), .Y(n_134) );
BUFx2_ASAP7_75t_L g135 ( .A(n_102), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_81), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_85), .B(n_0), .Y(n_137) );
AND2x6_ASAP7_75t_L g138 ( .A(n_81), .B(n_33), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_86), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_102), .B(n_1), .Y(n_140) );
OR2x2_ASAP7_75t_L g141 ( .A(n_85), .B(n_2), .Y(n_141) );
OR2x6_ASAP7_75t_L g142 ( .A(n_93), .B(n_2), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_88), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_88), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_91), .B(n_3), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_90), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_93), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_115), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_101), .B(n_3), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_117), .B(n_4), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_92), .B(n_4), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_90), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_117), .Y(n_155) );
OAI21x1_ASAP7_75t_L g156 ( .A1(n_118), .A2(n_36), .B(n_75), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_118), .Y(n_157) );
INVx5_ASAP7_75t_L g158 ( .A(n_80), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_121), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_105), .B(n_5), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_121), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_122), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_107), .B(n_6), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_122), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_110), .B(n_6), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_123), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_124), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_158), .B(n_82), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_158), .B(n_89), .Y(n_169) );
NOR2xp33_ASAP7_75t_SL g170 ( .A(n_132), .B(n_83), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_158), .B(n_83), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_125), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_135), .B(n_84), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_132), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_128), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_128), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_128), .Y(n_177) );
AND2x6_ASAP7_75t_L g178 ( .A(n_130), .B(n_123), .Y(n_178) );
BUFx4f_ASAP7_75t_L g179 ( .A(n_142), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_125), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_142), .A2(n_94), .B1(n_99), .B2(n_79), .Y(n_181) );
INVx8_ASAP7_75t_L g182 ( .A(n_158), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_128), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_128), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_125), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_136), .Y(n_186) );
NAND2x1p5_ASAP7_75t_L g187 ( .A(n_137), .B(n_104), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_124), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_136), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_137), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_124), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_124), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_135), .B(n_94), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_136), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_137), .Y(n_195) );
BUFx2_ASAP7_75t_L g196 ( .A(n_132), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_148), .B(n_99), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_136), .Y(n_198) );
BUFx2_ASAP7_75t_L g199 ( .A(n_132), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_158), .B(n_106), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_136), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_144), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_144), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_158), .B(n_130), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_144), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_144), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_130), .B(n_108), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_130), .B(n_116), .Y(n_208) );
INVx4_ASAP7_75t_L g209 ( .A(n_124), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_144), .Y(n_210) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_153), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_145), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_145), .Y(n_213) );
INVx1_ASAP7_75t_SL g214 ( .A(n_146), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_145), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_146), .Y(n_216) );
INVx1_ASAP7_75t_SL g217 ( .A(n_153), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_129), .B(n_103), .Y(n_218) );
NAND2x1p5_ASAP7_75t_L g219 ( .A(n_137), .B(n_98), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_145), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_149), .B(n_120), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_152), .B(n_97), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_145), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_174), .B(n_142), .Y(n_224) );
BUFx2_ASAP7_75t_L g225 ( .A(n_174), .Y(n_225) );
INVx2_ASAP7_75t_SL g226 ( .A(n_179), .Y(n_226) );
BUFx3_ASAP7_75t_L g227 ( .A(n_188), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_190), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_221), .B(n_147), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_196), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_197), .Y(n_231) );
NOR2x2_ASAP7_75t_L g232 ( .A(n_170), .B(n_142), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_197), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_196), .Y(n_234) );
OR2x2_ASAP7_75t_L g235 ( .A(n_214), .B(n_140), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_188), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_217), .A2(n_142), .B1(n_152), .B2(n_164), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_190), .Y(n_238) );
INVx2_ASAP7_75t_SL g239 ( .A(n_179), .Y(n_239) );
INVx2_ASAP7_75t_SL g240 ( .A(n_179), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_175), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_221), .B(n_157), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_211), .B(n_147), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_190), .Y(n_244) );
BUFx2_ASAP7_75t_L g245 ( .A(n_199), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_195), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_175), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_182), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_182), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_175), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_208), .B(n_143), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_195), .Y(n_252) );
INVx5_ASAP7_75t_L g253 ( .A(n_182), .Y(n_253) );
BUFx12f_ASAP7_75t_L g254 ( .A(n_199), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_208), .B(n_143), .Y(n_255) );
BUFx2_ASAP7_75t_L g256 ( .A(n_178), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_175), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_182), .Y(n_258) );
NOR2x1_ASAP7_75t_L g259 ( .A(n_193), .B(n_152), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_216), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_193), .B(n_157), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_195), .A2(n_152), .B(n_129), .C(n_164), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_172), .Y(n_263) );
BUFx2_ASAP7_75t_L g264 ( .A(n_178), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_178), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_178), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_178), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_182), .Y(n_268) );
INVx3_ASAP7_75t_L g269 ( .A(n_178), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_181), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_175), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_176), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_173), .B(n_154), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_187), .A2(n_141), .B1(n_133), .B2(n_154), .Y(n_274) );
INVx5_ASAP7_75t_L g275 ( .A(n_178), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_176), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_172), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_180), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_181), .Y(n_279) );
INVxp67_ASAP7_75t_L g280 ( .A(n_173), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_180), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_187), .Y(n_282) );
AND2x4_ASAP7_75t_L g283 ( .A(n_207), .B(n_141), .Y(n_283) );
INVx4_ASAP7_75t_L g284 ( .A(n_167), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_185), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_244), .Y(n_286) );
BUFx4f_ASAP7_75t_L g287 ( .A(n_254), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_254), .Y(n_288) );
A2O1A1Ixp33_ASAP7_75t_L g289 ( .A1(n_273), .A2(n_218), .B(n_222), .C(n_159), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_244), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g291 ( .A1(n_243), .A2(n_133), .B1(n_159), .B2(n_151), .C(n_160), .Y(n_291) );
AOI21x1_ASAP7_75t_L g292 ( .A1(n_228), .A2(n_185), .B(n_204), .Y(n_292) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_260), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_225), .B(n_204), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_283), .A2(n_187), .B1(n_219), .B2(n_207), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_244), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_283), .B(n_207), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_283), .B(n_207), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_228), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_238), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_275), .B(n_167), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_238), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_246), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_274), .A2(n_219), .B1(n_222), .B2(n_168), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_246), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_252), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_252), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_224), .A2(n_222), .B1(n_219), .B2(n_138), .Y(n_308) );
INVx3_ASAP7_75t_L g309 ( .A(n_253), .Y(n_309) );
AO32x2_ASAP7_75t_L g310 ( .A1(n_226), .A2(n_134), .A3(n_167), .B1(n_209), .B2(n_191), .Y(n_310) );
CKINVDCx11_ASAP7_75t_R g311 ( .A(n_225), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_263), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_245), .B(n_222), .Y(n_313) );
AND2x6_ASAP7_75t_L g314 ( .A(n_224), .B(n_192), .Y(n_314) );
AOI222xp33_ASAP7_75t_L g315 ( .A1(n_270), .A2(n_163), .B1(n_165), .B2(n_150), .C1(n_155), .C2(n_149), .Y(n_315) );
INVx4_ASAP7_75t_L g316 ( .A(n_253), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_229), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_242), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_245), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g320 ( .A(n_230), .Y(n_320) );
INVx6_ASAP7_75t_L g321 ( .A(n_224), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_253), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_251), .Y(n_323) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_262), .A2(n_162), .B(n_161), .C(n_139), .Y(n_324) );
INVx4_ASAP7_75t_L g325 ( .A(n_253), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_253), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_L g327 ( .A1(n_261), .A2(n_162), .B(n_161), .C(n_139), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_263), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_275), .B(n_167), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_253), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_255), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_259), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_277), .Y(n_333) );
AND3x1_ASAP7_75t_SL g334 ( .A(n_270), .B(n_78), .C(n_96), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_277), .Y(n_335) );
BUFx12f_ASAP7_75t_L g336 ( .A(n_230), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_312), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_333), .Y(n_338) );
BUFx2_ASAP7_75t_L g339 ( .A(n_314), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_294), .A2(n_279), .B1(n_233), .B2(n_231), .Y(n_340) );
AND2x4_ASAP7_75t_SL g341 ( .A(n_313), .B(n_282), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_322), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_295), .A2(n_237), .B1(n_282), .B2(n_235), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_317), .B(n_235), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_292), .A2(n_156), .B(n_285), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_294), .A2(n_279), .B1(n_280), .B2(n_282), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_322), .B(n_275), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_319), .B(n_234), .Y(n_348) );
INVx2_ASAP7_75t_SL g349 ( .A(n_316), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_335), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_318), .B(n_234), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_323), .B(n_226), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_308), .A2(n_239), .B1(n_240), .B2(n_256), .Y(n_353) );
BUFx10_ASAP7_75t_L g354 ( .A(n_314), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_313), .A2(n_239), .B1(n_240), .B2(n_264), .Y(n_355) );
INVx3_ASAP7_75t_L g356 ( .A(n_316), .Y(n_356) );
INVx1_ASAP7_75t_SL g357 ( .A(n_311), .Y(n_357) );
INVxp67_ASAP7_75t_SL g358 ( .A(n_320), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_331), .B(n_256), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_308), .A2(n_266), .B1(n_264), .B2(n_275), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_325), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_325), .B(n_275), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_304), .A2(n_266), .B1(n_232), .B2(n_265), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_288), .B(n_169), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_314), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_315), .A2(n_269), .B1(n_265), .B2(n_267), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_314), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_328), .Y(n_368) );
HB1xp67_ASAP7_75t_SL g369 ( .A(n_348), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_344), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_343), .A2(n_311), .B1(n_332), .B2(n_291), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_340), .A2(n_300), .B1(n_303), .B2(n_306), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_338), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_363), .A2(n_289), .B1(n_321), .B2(n_297), .Y(n_374) );
AOI22xp33_ASAP7_75t_SL g375 ( .A1(n_357), .A2(n_320), .B1(n_336), .B2(n_287), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_351), .B(n_348), .Y(n_376) );
OAI211xp5_ASAP7_75t_SL g377 ( .A1(n_346), .A2(n_126), .B(n_127), .C(n_334), .Y(n_377) );
AOI222xp33_ASAP7_75t_L g378 ( .A1(n_357), .A2(n_287), .B1(n_293), .B2(n_289), .C1(n_298), .C2(n_334), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_337), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_341), .B(n_309), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_351), .Y(n_381) );
OAI33xp33_ASAP7_75t_L g382 ( .A1(n_338), .A2(n_327), .A3(n_111), .B1(n_113), .B2(n_112), .B3(n_109), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_368), .A2(n_321), .B1(n_327), .B2(n_324), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_368), .A2(n_321), .B1(n_324), .B2(n_305), .Y(n_384) );
OAI22xp33_ASAP7_75t_L g385 ( .A1(n_358), .A2(n_293), .B1(n_326), .B2(n_330), .Y(n_385) );
OAI211xp5_ASAP7_75t_L g386 ( .A1(n_364), .A2(n_155), .B(n_150), .C(n_149), .Y(n_386) );
OAI22xp5_ASAP7_75t_SL g387 ( .A1(n_364), .A2(n_330), .B1(n_326), .B2(n_309), .Y(n_387) );
AOI21xp33_ASAP7_75t_L g388 ( .A1(n_349), .A2(n_299), .B(n_302), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_341), .B(n_150), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_350), .A2(n_307), .B1(n_155), .B2(n_166), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_352), .B(n_126), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g392 ( .A1(n_339), .A2(n_314), .B1(n_124), .B2(n_138), .Y(n_392) );
AOI222xp33_ASAP7_75t_L g393 ( .A1(n_350), .A2(n_127), .B1(n_126), .B2(n_200), .C1(n_124), .C2(n_138), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_359), .A2(n_127), .B1(n_278), .B2(n_285), .C(n_281), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_337), .A2(n_166), .B1(n_278), .B2(n_281), .Y(n_395) );
NOR2xp33_ASAP7_75t_R g396 ( .A(n_354), .B(n_265), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_371), .A2(n_366), .B1(n_355), .B2(n_359), .C(n_353), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_379), .B(n_356), .Y(n_398) );
OAI221xp5_ASAP7_75t_L g399 ( .A1(n_371), .A2(n_349), .B1(n_361), .B2(n_290), .C(n_356), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_379), .B(n_356), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_370), .B(n_342), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_373), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_380), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_384), .Y(n_404) );
INVx1_ASAP7_75t_SL g405 ( .A(n_369), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_380), .B(n_339), .Y(n_406) );
INVxp67_ASAP7_75t_L g407 ( .A(n_381), .Y(n_407) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_378), .A2(n_361), .B1(n_365), .B2(n_342), .C(n_87), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_374), .B(n_365), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_387), .A2(n_367), .B1(n_354), .B2(n_347), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_383), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_377), .A2(n_138), .B1(n_131), .B2(n_367), .Y(n_412) );
OAI31xp33_ASAP7_75t_L g413 ( .A1(n_385), .A2(n_360), .A3(n_200), .B(n_362), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_376), .B(n_367), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_382), .A2(n_138), .B1(n_131), .B2(n_367), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_372), .B(n_367), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_372), .B(n_345), .Y(n_417) );
OAI221xp5_ASAP7_75t_L g418 ( .A1(n_375), .A2(n_296), .B1(n_286), .B2(n_166), .C(n_171), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_389), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_391), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_388), .B(n_286), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_390), .B(n_345), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_395), .A2(n_166), .B1(n_347), .B2(n_362), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_386), .A2(n_166), .B1(n_134), .B2(n_203), .C(n_201), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_394), .B(n_347), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_396), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_395), .Y(n_427) );
OAI31xp33_ASAP7_75t_SL g428 ( .A1(n_392), .A2(n_156), .A3(n_362), .B(n_347), .Y(n_428) );
OAI211xp5_ASAP7_75t_L g429 ( .A1(n_390), .A2(n_134), .B(n_220), .C(n_215), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_393), .Y(n_430) );
OAI221xp5_ASAP7_75t_SL g431 ( .A1(n_413), .A2(n_194), .B1(n_223), .B2(n_220), .C(n_215), .Y(n_431) );
OAI21xp33_ASAP7_75t_L g432 ( .A1(n_428), .A2(n_405), .B(n_407), .Y(n_432) );
INVx2_ASAP7_75t_SL g433 ( .A(n_398), .Y(n_433) );
NOR3xp33_ASAP7_75t_L g434 ( .A(n_408), .B(n_134), .C(n_210), .Y(n_434) );
AOI33xp33_ASAP7_75t_L g435 ( .A1(n_405), .A2(n_194), .A3(n_223), .B1(n_198), .B2(n_201), .B3(n_210), .Y(n_435) );
OAI211xp5_ASAP7_75t_SL g436 ( .A1(n_428), .A2(n_198), .B(n_203), .C(n_205), .Y(n_436) );
AOI211xp5_ASAP7_75t_SL g437 ( .A1(n_423), .A2(n_362), .B(n_354), .C(n_269), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_413), .B(n_176), .C(n_205), .Y(n_438) );
BUFx3_ASAP7_75t_L g439 ( .A(n_403), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_402), .B(n_7), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g441 ( .A1(n_420), .A2(n_206), .B1(n_213), .B2(n_212), .C(n_186), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_402), .B(n_10), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_420), .A2(n_206), .B1(n_213), .B2(n_212), .C(n_186), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_402), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_420), .B(n_10), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_417), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_417), .B(n_11), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_423), .A2(n_329), .B(n_301), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_414), .B(n_11), .Y(n_449) );
INVx3_ASAP7_75t_L g450 ( .A(n_426), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_414), .B(n_13), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_416), .B(n_13), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_430), .A2(n_267), .B1(n_269), .B2(n_354), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_401), .Y(n_454) );
NAND4xp75_ASAP7_75t_L g455 ( .A(n_430), .B(n_396), .C(n_14), .D(n_301), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_416), .B(n_14), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_401), .B(n_138), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_426), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_411), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_398), .B(n_17), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_411), .A2(n_329), .B(n_191), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_411), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_400), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_400), .B(n_19), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_421), .Y(n_465) );
BUFx2_ASAP7_75t_L g466 ( .A(n_426), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_422), .B(n_21), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_422), .B(n_26), .Y(n_468) );
AND2x2_ASAP7_75t_SL g469 ( .A(n_409), .B(n_192), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_430), .B(n_138), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_409), .B(n_27), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_404), .B(n_28), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_421), .B(n_183), .Y(n_473) );
AOI22xp33_ASAP7_75t_SL g474 ( .A1(n_406), .A2(n_131), .B1(n_267), .B2(n_192), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_404), .B(n_34), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_404), .B(n_183), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_427), .B(n_37), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_419), .B(n_131), .Y(n_478) );
AOI211xp5_ASAP7_75t_SL g479 ( .A1(n_432), .A2(n_397), .B(n_418), .C(n_399), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_454), .B(n_403), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_442), .Y(n_481) );
NAND3xp33_ASAP7_75t_L g482 ( .A(n_447), .B(n_424), .C(n_410), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_446), .B(n_427), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_455), .A2(n_412), .B(n_425), .Y(n_484) );
INVx5_ASAP7_75t_L g485 ( .A(n_450), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_442), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_433), .B(n_403), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_463), .B(n_427), .Y(n_488) );
BUFx2_ASAP7_75t_L g489 ( .A(n_466), .Y(n_489) );
OAI21xp33_ASAP7_75t_L g490 ( .A1(n_447), .A2(n_415), .B(n_425), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_433), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_446), .B(n_403), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_437), .A2(n_406), .B(n_429), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_449), .B(n_403), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_465), .B(n_403), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_444), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_449), .B(n_406), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_444), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_452), .B(n_406), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_451), .B(n_131), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_466), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_452), .B(n_184), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_462), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_451), .B(n_131), .Y(n_504) );
INVxp67_ASAP7_75t_L g505 ( .A(n_440), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_456), .B(n_131), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_440), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_456), .B(n_445), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_439), .B(n_38), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_459), .B(n_184), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_467), .B(n_177), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_467), .B(n_177), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_445), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_462), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_473), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_459), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_450), .B(n_248), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_473), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_468), .B(n_45), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_450), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_468), .B(n_202), .Y(n_521) );
AO21x1_ASAP7_75t_L g522 ( .A1(n_471), .A2(n_189), .B(n_202), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_460), .B(n_189), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g524 ( .A(n_435), .B(n_176), .C(n_272), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_460), .B(n_47), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_469), .B(n_192), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_458), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_439), .B(n_52), .Y(n_528) );
INVx2_ASAP7_75t_SL g529 ( .A(n_458), .Y(n_529) );
BUFx2_ASAP7_75t_L g530 ( .A(n_458), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_471), .B(n_54), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_464), .B(n_57), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_471), .B(n_63), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_476), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_438), .A2(n_209), .B1(n_191), .B2(n_192), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_491), .B(n_464), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_489), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_513), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g539 ( .A(n_479), .B(n_436), .C(n_434), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_483), .B(n_469), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_508), .B(n_515), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_518), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_483), .B(n_477), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_496), .Y(n_544) );
BUFx2_ASAP7_75t_L g545 ( .A(n_501), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_507), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_499), .B(n_477), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_488), .B(n_472), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_498), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_480), .Y(n_550) );
AOI32xp33_ASAP7_75t_L g551 ( .A1(n_531), .A2(n_478), .A3(n_453), .B1(n_475), .B2(n_472), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_499), .B(n_475), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_495), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_495), .B(n_497), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_527), .Y(n_555) );
OAI21xp33_ASAP7_75t_L g556 ( .A1(n_520), .A2(n_431), .B(n_470), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_530), .Y(n_557) );
AOI211xp5_ASAP7_75t_L g558 ( .A1(n_482), .A2(n_448), .B(n_457), .C(n_476), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_494), .B(n_534), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_516), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_505), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_529), .B(n_461), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_534), .B(n_455), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_481), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_486), .B(n_64), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_526), .A2(n_474), .B(n_443), .Y(n_566) );
INVxp67_ASAP7_75t_L g567 ( .A(n_529), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_503), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_485), .B(n_441), .Y(n_569) );
NOR2x1_ASAP7_75t_R g570 ( .A(n_485), .B(n_249), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_514), .B(n_66), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_487), .Y(n_572) );
NAND4xp25_ASAP7_75t_SL g573 ( .A(n_531), .B(n_71), .C(n_74), .D(n_76), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_485), .Y(n_574) );
AND3x1_ASAP7_75t_L g575 ( .A(n_533), .B(n_257), .C(n_276), .Y(n_575) );
BUFx3_ASAP7_75t_L g576 ( .A(n_485), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_492), .B(n_257), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_490), .B(n_250), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_492), .B(n_310), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_510), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_502), .Y(n_581) );
NAND2x1_ASAP7_75t_L g582 ( .A(n_545), .B(n_533), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_538), .B(n_502), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_561), .B(n_485), .Y(n_584) );
XOR2x2_ASAP7_75t_L g585 ( .A(n_575), .B(n_526), .Y(n_585) );
AOI211xp5_ASAP7_75t_L g586 ( .A1(n_570), .A2(n_484), .B(n_522), .C(n_493), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_564), .B(n_512), .Y(n_587) );
NOR3xp33_ASAP7_75t_L g588 ( .A(n_539), .B(n_532), .C(n_525), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_546), .B(n_512), .Y(n_589) );
OAI21xp33_ASAP7_75t_L g590 ( .A1(n_557), .A2(n_519), .B(n_511), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_541), .B(n_522), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_572), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_555), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_567), .Y(n_594) );
AND2x4_ASAP7_75t_SL g595 ( .A(n_537), .B(n_509), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_550), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_559), .B(n_511), .Y(n_597) );
OAI211xp5_ASAP7_75t_L g598 ( .A1(n_569), .A2(n_506), .B(n_504), .C(n_500), .Y(n_598) );
XOR2xp5_ASAP7_75t_L g599 ( .A(n_536), .B(n_517), .Y(n_599) );
OAI21xp5_ASAP7_75t_L g600 ( .A1(n_569), .A2(n_524), .B(n_517), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_554), .B(n_528), .Y(n_601) );
NOR2xp67_ASAP7_75t_L g602 ( .A(n_573), .B(n_509), .Y(n_602) );
AOI321xp33_ASAP7_75t_L g603 ( .A1(n_558), .A2(n_521), .A3(n_528), .B1(n_523), .B2(n_509), .C(n_535), .Y(n_603) );
AND2x4_ASAP7_75t_SL g604 ( .A(n_581), .B(n_250), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_542), .B(n_241), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_553), .B(n_241), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_580), .B(n_276), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_549), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_543), .B(n_272), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_552), .B(n_547), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_567), .B(n_540), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_560), .Y(n_612) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_544), .Y(n_613) );
AOI21xp5_ASAP7_75t_SL g614 ( .A1(n_576), .A2(n_249), .B(n_268), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_568), .Y(n_615) );
OAI21xp33_ASAP7_75t_L g616 ( .A1(n_556), .A2(n_271), .B(n_247), .Y(n_616) );
AOI22xp5_ASAP7_75t_SL g617 ( .A1(n_576), .A2(n_248), .B1(n_268), .B2(n_258), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_563), .B(n_247), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_540), .A2(n_191), .B1(n_209), .B2(n_284), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_573), .A2(n_209), .B1(n_284), .B2(n_258), .Y(n_620) );
OAI21xp33_ASAP7_75t_L g621 ( .A1(n_548), .A2(n_227), .B(n_236), .Y(n_621) );
XNOR2x1_ASAP7_75t_L g622 ( .A(n_565), .B(n_227), .Y(n_622) );
INVx1_ASAP7_75t_SL g623 ( .A(n_574), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_579), .B(n_236), .Y(n_624) );
NOR2x1_ASAP7_75t_L g625 ( .A(n_566), .B(n_571), .Y(n_625) );
AO21x1_ASAP7_75t_L g626 ( .A1(n_566), .A2(n_571), .B(n_562), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_562), .B(n_551), .Y(n_627) );
OAI21xp33_ASAP7_75t_L g628 ( .A1(n_578), .A2(n_432), .B(n_538), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_577), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_577), .B(n_578), .Y(n_630) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_576), .Y(n_631) );
AOI222xp33_ASAP7_75t_L g632 ( .A1(n_539), .A2(n_371), .B1(n_405), .B2(n_432), .C1(n_407), .C2(n_376), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_538), .B(n_561), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_627), .A2(n_632), .B1(n_625), .B2(n_626), .Y(n_634) );
NAND3xp33_ASAP7_75t_SL g635 ( .A(n_586), .B(n_632), .C(n_600), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_633), .A2(n_591), .B1(n_596), .B2(n_628), .C(n_588), .Y(n_636) );
BUFx2_ASAP7_75t_L g637 ( .A(n_594), .Y(n_637) );
AOI322xp5_ASAP7_75t_L g638 ( .A1(n_592), .A2(n_611), .A3(n_591), .B1(n_610), .B2(n_594), .C1(n_582), .C2(n_601), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_623), .B(n_631), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_602), .A2(n_599), .B1(n_623), .B2(n_631), .Y(n_640) );
AOI22x1_ASAP7_75t_L g641 ( .A1(n_603), .A2(n_631), .B1(n_617), .B2(n_613), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_588), .A2(n_630), .B1(n_590), .B2(n_616), .Y(n_642) );
OAI21xp5_ASAP7_75t_L g643 ( .A1(n_585), .A2(n_614), .B(n_620), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_608), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_585), .A2(n_584), .B(n_595), .Y(n_645) );
XOR2xp5_ASAP7_75t_L g646 ( .A(n_622), .B(n_583), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_595), .A2(n_613), .B(n_587), .Y(n_647) );
OAI211xp5_ASAP7_75t_SL g648 ( .A1(n_634), .A2(n_598), .B(n_621), .C(n_589), .Y(n_648) );
XNOR2xp5_ASAP7_75t_L g649 ( .A(n_640), .B(n_593), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_644), .Y(n_650) );
OR3x2_ASAP7_75t_L g651 ( .A(n_635), .B(n_597), .C(n_609), .Y(n_651) );
XNOR2xp5_ASAP7_75t_L g652 ( .A(n_641), .B(n_629), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_637), .Y(n_653) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_643), .B(n_618), .C(n_624), .D(n_619), .Y(n_654) );
NOR5xp2_ASAP7_75t_L g655 ( .A(n_643), .B(n_615), .C(n_612), .D(n_604), .E(n_606), .Y(n_655) );
AND3x1_ASAP7_75t_L g656 ( .A(n_653), .B(n_636), .C(n_645), .Y(n_656) );
INVxp67_ASAP7_75t_SL g657 ( .A(n_655), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_650), .Y(n_658) );
OAI22xp5_ASAP7_75t_SL g659 ( .A1(n_652), .A2(n_646), .B1(n_642), .B2(n_638), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_659), .A2(n_651), .B1(n_648), .B2(n_649), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_658), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_657), .A2(n_654), .B1(n_647), .B2(n_639), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_661), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_660), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_664), .A2(n_662), .B1(n_656), .B2(n_654), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_665), .Y(n_666) );
OAI31xp33_ASAP7_75t_L g667 ( .A1(n_666), .A2(n_664), .A3(n_663), .B(n_619), .Y(n_667) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_667), .A2(n_605), .B(n_607), .Y(n_668) );
endmodule