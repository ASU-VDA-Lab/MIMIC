module fake_jpeg_8717_n_30 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_30);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_30;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_29;
wire n_15;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

OA22x2_ASAP7_75t_L g17 ( 
.A1(n_7),
.A2(n_2),
.B1(n_1),
.B2(n_5),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_21),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_6),
.B1(n_11),
.B2(n_10),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_20),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_0),
.Y(n_21)
);

AOI32xp33_ASAP7_75t_L g22 ( 
.A1(n_17),
.A2(n_14),
.A3(n_16),
.B1(n_9),
.B2(n_12),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_SL g25 ( 
.A1(n_22),
.A2(n_14),
.B(n_16),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_24),
.C(n_26),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_20),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_28),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_23),
.B(n_3),
.Y(n_30)
);


endmodule