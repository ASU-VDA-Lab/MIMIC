module fake_jpeg_30221_n_488 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_488);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_488;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_55),
.Y(n_109)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_61),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_64),
.Y(n_149)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_74),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_45),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_24),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_75),
.B(n_79),
.Y(n_136)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

BUFx4f_ASAP7_75t_SL g79 ( 
.A(n_22),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_24),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_80),
.B(n_81),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_35),
.B(n_16),
.C(n_15),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_25),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_82),
.B(n_85),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

BUFx16f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

BUFx16f_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_38),
.B1(n_41),
.B2(n_33),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_100),
.A2(n_41),
.B1(n_33),
.B2(n_26),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_56),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_102),
.B(n_113),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_103),
.B(n_55),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_53),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_82),
.A2(n_20),
.B(n_44),
.C(n_42),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_127),
.B(n_29),
.Y(n_194)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

BUFx12_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

HAxp5_ASAP7_75t_SL g137 ( 
.A(n_51),
.B(n_20),
.CON(n_137),
.SN(n_137)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_74),
.Y(n_162)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_60),
.Y(n_153)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_157),
.Y(n_238)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_159),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_160),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_161),
.A2(n_168),
.B1(n_169),
.B2(n_172),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_162),
.B(n_141),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_109),
.B(n_79),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_164),
.B(n_198),
.Y(n_225)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_165),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_109),
.B(n_29),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_166),
.B(n_171),
.Y(n_212)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

INVx4_ASAP7_75t_SL g220 ( 
.A(n_167),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_137),
.A2(n_52),
.B1(n_63),
.B2(n_89),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_124),
.A2(n_87),
.B1(n_83),
.B2(n_77),
.Y(n_169)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_145),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_106),
.A2(n_61),
.B1(n_69),
.B2(n_91),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_108),
.Y(n_177)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_104),
.Y(n_180)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_101),
.Y(n_183)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_184),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_139),
.B(n_40),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_185),
.B(n_194),
.Y(n_247)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_126),
.Y(n_186)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_186),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_42),
.B(n_26),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_103),
.C(n_122),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_188),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_107),
.A2(n_65),
.B1(n_72),
.B2(n_62),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_189),
.A2(n_195),
.B1(n_146),
.B2(n_154),
.Y(n_228)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_112),
.Y(n_190)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_192),
.Y(n_248)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_121),
.Y(n_193)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_193),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_132),
.A2(n_72),
.B1(n_62),
.B2(n_91),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_L g196 ( 
.A1(n_123),
.A2(n_64),
.B1(n_49),
.B2(n_44),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_196),
.A2(n_200),
.B1(n_123),
.B2(n_147),
.Y(n_240)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_128),
.Y(n_197)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_197),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_145),
.B(n_49),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_117),
.Y(n_199)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_136),
.A2(n_40),
.B1(n_25),
.B2(n_24),
.Y(n_200)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_136),
.B(n_16),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_205),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_128),
.B(n_15),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_142),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_114),
.B(n_15),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_209),
.Y(n_221)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_119),
.Y(n_208)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_156),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_211),
.B(n_219),
.Y(n_284)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_162),
.B(n_120),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_251),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_181),
.B(n_125),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_227),
.B(n_167),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

INVx13_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_240),
.A2(n_199),
.B1(n_183),
.B2(n_191),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_196),
.A2(n_150),
.B1(n_152),
.B2(n_135),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_242),
.A2(n_208),
.B1(n_175),
.B2(n_174),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_187),
.B(n_151),
.C(n_116),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_243),
.B(n_21),
.Y(n_290)
);

O2A1O1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_161),
.A2(n_133),
.B(n_37),
.C(n_110),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_193),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_189),
.A2(n_131),
.B(n_111),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_246),
.A2(n_157),
.B1(n_192),
.B2(n_158),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_253),
.A2(n_285),
.B1(n_218),
.B2(n_215),
.Y(n_303)
);

AND2x6_ASAP7_75t_L g255 ( 
.A(n_213),
.B(n_211),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_258),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_230),
.A2(n_195),
.B(n_177),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_256),
.A2(n_269),
.B(n_287),
.Y(n_295)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_257),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_233),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_259),
.B(n_267),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_206),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_260),
.B(n_265),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_262),
.A2(n_289),
.B1(n_220),
.B2(n_222),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_221),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_263),
.B(n_282),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_173),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_238),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_266),
.Y(n_317)
);

AND2x6_ASAP7_75t_L g267 ( 
.A(n_212),
.B(n_178),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_216),
.A2(n_201),
.B1(n_170),
.B2(n_203),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_268),
.A2(n_224),
.B1(n_231),
.B2(n_248),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_251),
.A2(n_165),
.B1(n_159),
.B2(n_209),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_270),
.Y(n_300)
);

AND2x6_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_219),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_271),
.B(n_272),
.Y(n_319)
);

NAND3xp33_ASAP7_75t_L g272 ( 
.A(n_217),
.B(n_235),
.C(n_219),
.Y(n_272)
);

INVx13_ASAP7_75t_L g273 ( 
.A(n_223),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_273),
.Y(n_316)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_244),
.Y(n_274)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_274),
.Y(n_302)
);

AND2x6_ASAP7_75t_L g275 ( 
.A(n_216),
.B(n_163),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_275),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_237),
.B(n_184),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_276),
.B(n_281),
.Y(n_323)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_277),
.Y(n_305)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_238),
.Y(n_278)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_234),
.Y(n_279)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_279),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_280),
.A2(n_220),
.B1(n_222),
.B2(n_214),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_226),
.B(n_188),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_242),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_239),
.Y(n_283)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_283),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_234),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_288),
.Y(n_309)
);

NOR3xp33_ASAP7_75t_SL g287 ( 
.A(n_245),
.B(n_163),
.C(n_188),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_226),
.B(n_184),
.Y(n_288)
);

OA22x2_ASAP7_75t_L g289 ( 
.A1(n_240),
.A2(n_176),
.B1(n_37),
.B2(n_149),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_224),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_231),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_291),
.B(n_313),
.C(n_315),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_292),
.A2(n_304),
.B1(n_308),
.B2(n_279),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_293),
.B(n_105),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_296),
.B(n_306),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_214),
.B1(n_248),
.B2(n_218),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_297),
.A2(n_303),
.B1(n_310),
.B2(n_322),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_256),
.A2(n_254),
.B(n_284),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_299),
.A2(n_312),
.B(n_268),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_301),
.A2(n_317),
.B(n_320),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_263),
.A2(n_215),
.B1(n_232),
.B2(n_229),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_229),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_254),
.A2(n_232),
.B1(n_239),
.B2(n_202),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_289),
.A2(n_252),
.B1(n_241),
.B2(n_176),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_264),
.A2(n_236),
.B(n_223),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_210),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_264),
.B(n_255),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_262),
.A2(n_252),
.B1(n_241),
.B2(n_236),
.Y(n_322)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_274),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_325),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_275),
.C(n_271),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_329),
.B(n_355),
.C(n_296),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_298),
.B(n_267),
.Y(n_330)
);

NAND3xp33_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_335),
.C(n_300),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_331),
.A2(n_334),
.B1(n_342),
.B2(n_349),
.Y(n_372)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_302),
.Y(n_332)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_332),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_333),
.B(n_297),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_318),
.A2(n_304),
.B1(n_292),
.B2(n_307),
.Y(n_334)
);

NOR3xp33_ASAP7_75t_SL g335 ( 
.A(n_319),
.B(n_287),
.C(n_261),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_294),
.B(n_257),
.Y(n_336)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_336),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_307),
.B(n_277),
.Y(n_337)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_337),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_323),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_338),
.B(n_341),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_295),
.A2(n_289),
.B1(n_280),
.B2(n_278),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_339),
.A2(n_351),
.B1(n_317),
.B2(n_21),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_309),
.B(n_289),
.Y(n_340)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_340),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_270),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_295),
.A2(n_261),
.B1(n_266),
.B2(n_283),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_316),
.B(n_273),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_343),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_302),
.B(n_266),
.Y(n_344)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_344),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_345),
.B(n_346),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_299),
.A2(n_210),
.B(n_105),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_312),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_322),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_306),
.A2(n_14),
.B1(n_13),
.B2(n_3),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_305),
.Y(n_350)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_350),
.Y(n_377)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_305),
.Y(n_352)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_352),
.Y(n_380)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_325),
.Y(n_353)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_353),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_324),
.A2(n_21),
.B1(n_1),
.B2(n_3),
.Y(n_354)
);

INVxp33_ASAP7_75t_L g376 ( 
.A(n_354),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_291),
.B(n_21),
.C(n_14),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_316),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_356),
.B(n_338),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_355),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_313),
.C(n_321),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_359),
.B(n_368),
.C(n_371),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_361),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_293),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_363),
.B(n_378),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_367),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_329),
.B(n_314),
.C(n_320),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_370),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_347),
.B(n_314),
.C(n_300),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_374),
.B(n_326),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_337),
.B(n_317),
.Y(n_375)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_375),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_347),
.B(n_311),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_348),
.B(n_311),
.C(n_324),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_379),
.B(n_345),
.C(n_333),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_381),
.A2(n_331),
.B1(n_340),
.B2(n_334),
.Y(n_389)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_344),
.Y(n_383)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_383),
.Y(n_403)
);

AOI21x1_ASAP7_75t_SL g384 ( 
.A1(n_351),
.A2(n_0),
.B(n_1),
.Y(n_384)
);

AO21x1_ASAP7_75t_L g400 ( 
.A1(n_384),
.A2(n_351),
.B(n_353),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_358),
.B(n_330),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_385),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_384),
.A2(n_356),
.B1(n_346),
.B2(n_332),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_388),
.A2(n_381),
.B1(n_362),
.B2(n_369),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_389),
.A2(n_362),
.B1(n_369),
.B2(n_383),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_391),
.B(n_405),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_397),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_379),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_400),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_352),
.Y(n_396)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_396),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_377),
.Y(n_397)
);

INVxp33_ASAP7_75t_L g398 ( 
.A(n_366),
.Y(n_398)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_398),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_401),
.C(n_407),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_368),
.B(n_350),
.C(n_327),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_402),
.B(n_374),
.Y(n_417)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_377),
.Y(n_404)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_404),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_349),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_327),
.Y(n_406)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_406),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_326),
.C(n_335),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_371),
.B(n_13),
.C(n_1),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_408),
.B(n_359),
.C(n_365),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_387),
.A2(n_370),
.B(n_372),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_411),
.A2(n_400),
.B(n_389),
.Y(n_434)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_396),
.Y(n_415)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_415),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_421),
.Y(n_433)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_406),
.Y(n_418)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_418),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_419),
.A2(n_387),
.B1(n_394),
.B2(n_399),
.Y(n_429)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_403),
.Y(n_420)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_420),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_357),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_422),
.A2(n_427),
.B1(n_418),
.B2(n_409),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_423),
.B(n_391),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_386),
.B(n_364),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_426),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_438),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_401),
.C(n_393),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_441),
.C(n_390),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_431),
.B(n_439),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_434),
.A2(n_438),
.B(n_437),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_410),
.A2(n_407),
.B1(n_382),
.B2(n_380),
.Y(n_435)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_435),
.Y(n_451)
);

INVx13_ASAP7_75t_L g436 ( 
.A(n_416),
.Y(n_436)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_436),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_419),
.A2(n_402),
.B1(n_398),
.B2(n_408),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_395),
.C(n_390),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_416),
.B(n_382),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_442),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_436),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_443),
.B(n_450),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_428),
.B(n_424),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_446),
.B(n_447),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_439),
.B(n_417),
.Y(n_448)
);

AO21x1_ASAP7_75t_L g464 ( 
.A1(n_448),
.A2(n_449),
.B(n_456),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_441),
.A2(n_414),
.B(n_423),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_434),
.A2(n_414),
.B(n_411),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_395),
.C(n_413),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_453),
.B(n_454),
.C(n_376),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_433),
.B(n_413),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_421),
.C(n_429),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_458),
.C(n_461),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_453),
.B(n_433),
.C(n_437),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_454),
.B(n_442),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_460),
.B(n_466),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_455),
.B(n_432),
.C(n_420),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_451),
.A2(n_415),
.B1(n_432),
.B2(n_440),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_462),
.B(n_444),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_440),
.C(n_425),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_465),
.B(n_443),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_445),
.B(n_380),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_467),
.B(n_450),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_468),
.B(n_470),
.Y(n_477)
);

AOI322xp5_ASAP7_75t_L g476 ( 
.A1(n_471),
.A2(n_473),
.A3(n_474),
.B1(n_464),
.B2(n_376),
.C1(n_4),
.C2(n_5),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_459),
.A2(n_444),
.B(n_452),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_463),
.A2(n_448),
.B(n_456),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_470),
.A2(n_464),
.B1(n_463),
.B2(n_467),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_475),
.B(n_476),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_472),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_478),
.B(n_12),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_477),
.B(n_469),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_480),
.B(n_481),
.Y(n_483)
);

NAND2x1_ASAP7_75t_L g482 ( 
.A(n_479),
.B(n_475),
.Y(n_482)
);

AOI31xp33_ASAP7_75t_L g484 ( 
.A1(n_482),
.A2(n_6),
.A3(n_7),
.B(n_10),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_484),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_485),
.Y(n_486)
);

OAI321xp33_ASAP7_75t_L g487 ( 
.A1(n_486),
.A2(n_482),
.A3(n_483),
.B1(n_11),
.B2(n_6),
.C(n_7),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_487),
.A2(n_7),
.B1(n_11),
.B2(n_356),
.Y(n_488)
);


endmodule