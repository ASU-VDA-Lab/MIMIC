module real_jpeg_18678_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_535),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_0),
.B(n_536),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_1),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_1),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_1),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_1),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_1),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_1),
.B(n_189),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_1),
.B(n_94),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_2),
.Y(n_94)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_2),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_2),
.Y(n_381)
);

BUFx5_ASAP7_75t_L g390 ( 
.A(n_2),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_3),
.Y(n_96)
);

NAND2x1_ASAP7_75t_L g97 ( 
.A(n_3),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_3),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_3),
.B(n_253),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_3),
.B(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_3),
.B(n_339),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_3),
.B(n_385),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_3),
.B(n_94),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_4),
.Y(n_112)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_4),
.Y(n_157)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_4),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g396 ( 
.A(n_4),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_5),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_5),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_5),
.B(n_34),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_5),
.B(n_300),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_5),
.B(n_341),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_5),
.B(n_446),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_5),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_5),
.B(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_6),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_6),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_6),
.B(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_6),
.B(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_6),
.B(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_6),
.B(n_489),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_6),
.B(n_497),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_7),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_7),
.Y(n_298)
);

BUFx5_ASAP7_75t_L g438 ( 
.A(n_7),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_8),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_8),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_8),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_8),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_8),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_8),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_8),
.B(n_48),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_8),
.A2(n_12),
.B1(n_274),
.B2(n_277),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_8),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_9),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_9),
.B(n_70),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_9),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_9),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_9),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_9),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_9),
.B(n_298),
.Y(n_297)
);

AND2x2_ASAP7_75t_SL g334 ( 
.A(n_9),
.B(n_94),
.Y(n_334)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_10),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g249 ( 
.A(n_10),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_10),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_11),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_11),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_11),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_11),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_11),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_12),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_12),
.B(n_230),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_12),
.B(n_337),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_12),
.B(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_12),
.B(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_12),
.B(n_438),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_12),
.B(n_442),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_12),
.B(n_474),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_13),
.Y(n_240)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_14),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_14),
.Y(n_206)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_14),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_14),
.Y(n_290)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_14),
.Y(n_417)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_15),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_16),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_16),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_16),
.B(n_36),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_16),
.B(n_232),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_16),
.B(n_294),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g333 ( 
.A(n_16),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_16),
.B(n_388),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_17),
.Y(n_102)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_18),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_18),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_168),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_166),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_140),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_23),
.B(n_140),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_103),
.C(n_115),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_24),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_74),
.C(n_90),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_26),
.B(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_42),
.C(n_58),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_27),
.B(n_42),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_28),
.B(n_33),
.C(n_38),
.Y(n_114)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_30),
.B(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_37),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g337 ( 
.A(n_37),
.Y(n_337)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.C(n_51),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_43),
.B(n_51),
.Y(n_184)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_47),
.B(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_50),
.Y(n_339)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_58),
.B(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_69),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_60),
.A2(n_61),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_61),
.B(n_65),
.C(n_69),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_SL g130 ( 
.A(n_61),
.B(n_106),
.C(n_109),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_64),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_65),
.A2(n_66),
.B1(n_93),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_93),
.C(n_95),
.Y(n_92)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_68),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_68),
.Y(n_499)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_73),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_74),
.B(n_90),
.Y(n_177)
);

XNOR2x1_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_81),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_85),
.C(n_89),
.Y(n_128)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_80),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_89),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g436 ( 
.A(n_88),
.Y(n_436)
);

MAJx2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.C(n_99),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_91),
.A2(n_92),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_93),
.B(n_186),
.C(n_188),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_93),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_93),
.A2(n_188),
.B1(n_196),
.B2(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_95),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_95),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_95),
.A2(n_193),
.B1(n_282),
.B2(n_330),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_97),
.B(n_99),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_97),
.B(n_245),
.C(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_97),
.Y(n_270)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_99),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_99),
.A2(n_208),
.B1(n_211),
.B2(n_257),
.Y(n_256)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_102),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_103),
.A2(n_115),
.B1(n_116),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_113),
.C(n_114),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_104),
.B(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_106),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_108),
.B(n_132),
.C(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_113),
.B(n_114),
.Y(n_179)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_129),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_130),
.C(n_131),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_128),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_122),
.C(n_128),
.Y(n_142)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_127),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

XOR2x1_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_147),
.B1(n_148),
.B2(n_152),
.Y(n_146)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_165),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_158),
.B2(n_159),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_153),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_156),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_160),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_162),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_215),
.B(n_532),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_170),
.A2(n_533),
.B(n_534),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

NOR2xp67_ASAP7_75t_SL g534 ( 
.A(n_171),
.B(n_174),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.C(n_180),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_178),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_180),
.B(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_197),
.C(n_212),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.C(n_192),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_183),
.B(n_185),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_190),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_191),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_192),
.B(n_313),
.Y(n_312)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_193),
.B(n_281),
.C(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_212),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_208),
.C(n_211),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_198),
.B(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.C(n_207),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_207),
.Y(n_242)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_203),
.B(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_208),
.Y(n_257)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_210),
.Y(n_292)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_213),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_261),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_258),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_218),
.B(n_258),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.C(n_223),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_219),
.B(n_221),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_223),
.B(n_351),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_243),
.C(n_255),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_224),
.B(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.C(n_241),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_225),
.B(n_228),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.C(n_236),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_229),
.A2(n_236),
.B1(n_237),
.B2(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_229),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_231),
.B(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_235),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_236),
.B(n_411),
.C(n_413),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_236),
.A2(n_237),
.B1(n_411),
.B2(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2x2_ASAP7_75t_SL g322 ( 
.A(n_241),
.B(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_243),
.B(n_255),
.Y(n_311)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_250),
.C(n_251),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_244),
.B(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_246),
.Y(n_271)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_250),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_251),
.A2(n_252),
.B1(n_392),
.B2(n_393),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_252),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_254),
.Y(n_375)
);

AO21x2_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_355),
.B(n_529),
.Y(n_261)
);

NOR2xp67_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_349),
.Y(n_262)
);

AND2x2_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_316),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_264),
.B(n_316),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_309),
.Y(n_264)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_265),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_285),
.C(n_304),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_267),
.B(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_272),
.C(n_280),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_268),
.B(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_272),
.A2(n_273),
.B1(n_280),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_273),
.A2(n_371),
.B(n_376),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx6_ASAP7_75t_L g447 ( 
.A(n_275),
.Y(n_447)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_276),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_280),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_281),
.B(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_282),
.Y(n_330)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_284),
.B(n_333),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_285),
.A2(n_305),
.B1(n_306),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_285),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_296),
.C(n_299),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_286),
.B(n_344),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_291),
.C(n_293),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_287),
.A2(n_293),
.B1(n_368),
.B2(n_369),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_287),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_287),
.B(n_433),
.Y(n_432)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_291),
.B(n_367),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_293),
.Y(n_369)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_296),
.A2(n_297),
.B1(n_299),
.B2(n_345),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_299),
.Y(n_345)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_310),
.A2(n_312),
.B1(n_314),
.B2(n_315),
.Y(n_309)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_310),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_312),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_312),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_314),
.B(n_353),
.C(n_354),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_322),
.C(n_324),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_318),
.A2(n_319),
.B1(n_322),
.B2(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_322),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_359),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_343),
.C(n_346),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_326),
.B(n_364),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_331),
.C(n_335),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_328),
.B(n_422),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_331),
.B(n_335),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_334),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_332),
.B(n_334),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_338),
.C(n_340),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_336),
.A2(n_338),
.B1(n_407),
.B2(n_408),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_336),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_338),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_338),
.A2(n_408),
.B1(n_483),
.B2(n_484),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_338),
.B(n_479),
.C(n_483),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_340),
.B(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_346),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_349),
.A2(n_530),
.B(n_531),
.Y(n_529)
);

AND2x2_ASAP7_75t_SL g349 ( 
.A(n_350),
.B(n_352),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_350),
.B(n_352),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_425),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_361),
.C(n_400),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_358),
.B(n_362),
.Y(n_528)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_365),
.C(n_397),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_363),
.B(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_365),
.B(n_397),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_370),
.C(n_382),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_366),
.B(n_370),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_368),
.B(n_434),
.C(n_437),
.Y(n_458)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_403),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_391),
.C(n_392),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_383),
.B(n_515),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_387),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_384),
.B(n_387),
.Y(n_465)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_384),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_384),
.A2(n_472),
.B1(n_473),
.B2(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

NOR2x1_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_423),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_423),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.C(n_420),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_402),
.B(n_526),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_404),
.B(n_421),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_409),
.C(n_418),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_405),
.B(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_410),
.B(n_419),
.Y(n_520)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_411),
.Y(n_461)
);

XOR2x2_ASAP7_75t_L g459 ( 
.A(n_413),
.B(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_417),
.Y(n_485)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NAND3xp33_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_427),
.C(n_528),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_428),
.A2(n_523),
.B(n_527),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_509),
.B(n_522),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_468),
.B(n_508),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_456),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_431),
.B(n_456),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_439),
.C(n_448),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_432),
.B(n_504),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_437),
.Y(n_433)
);

INVx5_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_438),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_439),
.A2(n_440),
.B1(n_448),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_445),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_441),
.B(n_445),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx6_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_448),
.Y(n_505)
);

AO22x1_ASAP7_75t_SL g448 ( 
.A1(n_449),
.A2(n_453),
.B1(n_454),
.B2(n_455),
.Y(n_448)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_449),
.Y(n_454)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_453),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_453),
.B(n_454),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_455),
.B(n_496),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_462),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_458),
.B(n_459),
.C(n_462),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

MAJx2_ASAP7_75t_L g517 ( 
.A(n_463),
.B(n_465),
.C(n_466),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_469),
.A2(n_502),
.B(n_507),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_470),
.A2(n_486),
.B(n_501),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_478),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_471),
.B(n_478),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_473),
.Y(n_494)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx4_ASAP7_75t_SL g475 ( 
.A(n_476),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_479),
.A2(n_480),
.B1(n_481),
.B2(n_482),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_487),
.A2(n_495),
.B(n_500),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_493),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_493),
.Y(n_500)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_503),
.B(n_506),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_503),
.B(n_506),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_510),
.B(n_521),
.Y(n_509)
);

NOR2xp67_ASAP7_75t_SL g522 ( 
.A(n_510),
.B(n_521),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_511),
.A2(n_512),
.B1(n_518),
.B2(n_519),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_513),
.A2(n_514),
.B1(n_516),
.B2(n_517),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_517),
.C(n_518),
.Y(n_524)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

NOR2x1_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_525),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_524),
.B(n_525),
.Y(n_527)
);


endmodule