module fake_jpeg_30398_n_178 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_22),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_3),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_25),
.Y(n_70)
);

INVx11_ASAP7_75t_SL g71 ( 
.A(n_4),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_76),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_0),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_80),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_1),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_1),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_54),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_76),
.B(n_70),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_59),
.B1(n_50),
.B2(n_48),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_93),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_50),
.B1(n_48),
.B2(n_62),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_60),
.Y(n_102)
);

CKINVDCx9p33_ASAP7_75t_R g96 ( 
.A(n_74),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_96),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_65),
.B1(n_61),
.B2(n_68),
.Y(n_97)
);

OR2x4_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_65),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_107),
.Y(n_131)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

NAND2x1_ASAP7_75t_SL g105 ( 
.A(n_96),
.B(n_73),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_5),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g107 ( 
.A(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_49),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_111),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_87),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_83),
.B(n_72),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_8),
.B1(n_10),
.B2(n_47),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_114),
.Y(n_135)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_101),
.A3(n_111),
.B1(n_99),
.B2(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_130),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_109),
.B(n_64),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_121),
.B(n_124),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_51),
.B1(n_66),
.B2(n_58),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_126),
.B1(n_133),
.B2(n_137),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_2),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_117),
.A2(n_51),
.B1(n_73),
.B2(n_6),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_4),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_128),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_28),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_114),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_8),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_15),
.Y(n_150)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_10),
.B(n_11),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_146),
.B(n_153),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_12),
.B(n_14),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_147),
.B(n_149),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_135),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_151),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_16),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_154),
.B(n_20),
.Y(n_162)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_156),
.B(n_148),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_136),
.A3(n_128),
.B1(n_135),
.B2(n_21),
.Y(n_157)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_162),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_155),
.A2(n_17),
.B(n_18),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_143),
.C(n_144),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_164),
.C(n_156),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_141),
.Y(n_167)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_167),
.A2(n_163),
.B(n_158),
.C(n_145),
.D(n_149),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_170),
.C(n_168),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_166),
.B1(n_167),
.B2(n_32),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_29),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_30),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_33),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_154),
.C(n_36),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_35),
.C(n_38),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_42),
.Y(n_178)
);


endmodule