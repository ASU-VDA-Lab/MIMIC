module real_jpeg_11642_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_300;
wire n_292;
wire n_215;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_285;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

INVx4_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_5),
.A2(n_56),
.B1(n_58),
.B2(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_5),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_5),
.A2(n_61),
.B1(n_62),
.B2(n_105),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_5),
.A2(n_38),
.B1(n_42),
.B2(n_105),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_105),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_6),
.A2(n_38),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_6),
.A2(n_45),
.B1(n_61),
.B2(n_62),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_45),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_7),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_8),
.A2(n_56),
.B1(n_58),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_8),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_8),
.A2(n_61),
.B1(n_62),
.B2(n_146),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_8),
.A2(n_38),
.B1(n_42),
.B2(n_146),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_146),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_9),
.A2(n_34),
.B1(n_56),
.B2(n_58),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_9),
.A2(n_34),
.B1(n_38),
.B2(n_42),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_9),
.A2(n_34),
.B1(n_61),
.B2(n_62),
.Y(n_149)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_11),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_11),
.B(n_107),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_11),
.B(n_27),
.C(n_41),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_11),
.A2(n_38),
.B1(n_42),
.B2(n_161),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_11),
.A2(n_24),
.B1(n_31),
.B2(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_11),
.B(n_83),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_12),
.A2(n_56),
.B1(n_58),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_12),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_12),
.A2(n_61),
.B1(n_62),
.B2(n_169),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_12),
.A2(n_38),
.B1(n_42),
.B2(n_169),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_169),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_13),
.A2(n_61),
.B1(n_62),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_13),
.A2(n_38),
.B1(n_42),
.B2(n_77),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_13),
.A2(n_56),
.B1(n_58),
.B2(n_77),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_77),
.Y(n_158)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_15),
.A2(n_38),
.B1(n_42),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_15),
.A2(n_48),
.B1(n_56),
.B2(n_58),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_48),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_15),
.A2(n_48),
.B1(n_61),
.B2(n_62),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_130),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_108),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_19),
.B(n_108),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_67),
.C(n_86),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_20),
.A2(n_21),
.B1(n_67),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_49),
.Y(n_21)
);

AOI21xp33_ASAP7_75t_L g109 ( 
.A1(n_22),
.A2(n_23),
.B(n_51),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_23),
.A2(n_50),
.B1(n_51),
.B2(n_66),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_23),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_23),
.A2(n_35),
.B1(n_66),
.B2(n_178),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B(n_32),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_24),
.A2(n_137),
.B(n_139),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_24),
.A2(n_31),
.B1(n_251),
.B2(n_259),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_24),
.A2(n_95),
.B(n_253),
.Y(n_273)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_25),
.B(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_25),
.A2(n_30),
.B1(n_138),
.B2(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_25),
.A2(n_33),
.B(n_140),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_25),
.A2(n_30),
.B1(n_250),
.B2(n_252),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_27),
.B1(n_39),
.B2(n_41),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_26),
.B(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_30),
.B(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_31),
.B(n_94),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_31),
.A2(n_92),
.B(n_158),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_31),
.B(n_161),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_35),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_44),
.B(n_46),
.Y(n_35)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_36),
.A2(n_44),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_36),
.A2(n_71),
.B(n_98),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_36),
.A2(n_46),
.B(n_71),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_36),
.A2(n_69),
.B(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_36),
.A2(n_98),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_36),
.A2(n_98),
.B1(n_225),
.B2(n_248),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_37)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

OA22x2_ASAP7_75t_SL g82 ( 
.A1(n_38),
.A2(n_42),
.B1(n_80),
.B2(n_81),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_38),
.A2(n_80),
.B(n_220),
.C(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_38),
.B(n_244),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_SL g41 ( 
.A(n_39),
.Y(n_41)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_L g221 ( 
.A(n_42),
.B(n_62),
.C(n_81),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_43),
.A2(n_73),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_73),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_63),
.B(n_64),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_52),
.A2(n_107),
.B1(n_160),
.B2(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_53),
.A2(n_104),
.B(n_106),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_53),
.B(n_65),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_53),
.A2(n_60),
.B1(n_104),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_53),
.A2(n_60),
.B1(n_145),
.B2(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_55),
.A2(n_62),
.B(n_160),
.C(n_162),
.Y(n_159)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_56),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

HAxp5_ASAP7_75t_SL g160 ( 
.A(n_58),
.B(n_161),
.CON(n_160),
.SN(n_160)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_58),
.B(n_59),
.C(n_61),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_62),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g220 ( 
.A(n_62),
.B(n_161),
.CON(n_220),
.SN(n_220)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_67),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_74),
.B(n_85),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_74),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_72),
.A2(n_97),
.B(n_98),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B1(n_83),
.B2(n_84),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_82),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_101),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_78),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_78),
.A2(n_122),
.B(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_78),
.A2(n_83),
.B1(n_197),
.B2(n_220),
.Y(n_222)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_102),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_82),
.A2(n_119),
.B1(n_164),
.B2(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_82),
.A2(n_119),
.B1(n_188),
.B2(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_83),
.B(n_149),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_111),
.B1(n_112),
.B2(n_127),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_86),
.A2(n_87),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_99),
.C(n_103),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_88),
.A2(n_89),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_96),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_90),
.A2(n_91),
.B1(n_96),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_96),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_98),
.B(n_161),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_99),
.B(n_103),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_116),
.B1(n_125),
.B2(n_126),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_123),
.B2(n_124),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B(n_121),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_119),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_123),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_294),
.B(n_300),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_180),
.B(n_293),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_170),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_133),
.B(n_170),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_150),
.C(n_152),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_134),
.B(n_150),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_142),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_143),
.C(n_148),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_141),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_136),
.B(n_141),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_147),
.B2(n_148),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_152),
.B(n_291),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_163),
.C(n_166),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_153),
.A2(n_154),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_155),
.A2(n_156),
.B1(n_159),
.B2(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_166),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_179),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_172),
.B(n_177),
.C(n_179),
.Y(n_299)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_208),
.B(n_288),
.C(n_292),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_201),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_201),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_191),
.C(n_194),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_183),
.B(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_186),
.C(n_190),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_189),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_194),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.C(n_200),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_195),
.B(n_229),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_202),
.B(n_206),
.C(n_207),
.Y(n_289)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_203),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_282),
.B(n_287),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_237),
.B(n_281),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_227),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_213),
.B(n_227),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_222),
.C(n_223),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_214),
.A2(n_215),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_216),
.B(n_219),
.Y(n_232)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_222),
.B(n_223),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_226),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_228),
.B(n_233),
.C(n_235),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_275),
.B(n_280),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_265),
.B(n_274),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_254),
.B(n_264),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_249),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_249),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_260),
.B(n_263),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_262),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_267),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_273),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_272),
.C(n_273),
.Y(n_279)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_279),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_279),
.Y(n_280)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_286),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_290),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_299),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_299),
.Y(n_300)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);


endmodule