module fake_jpeg_1787_n_203 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_203);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

INVx11_ASAP7_75t_SL g54 ( 
.A(n_11),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_22),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_33),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_76),
.Y(n_83)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_79),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_0),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_94),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_50),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_51),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_62),
.B1(n_71),
.B2(n_79),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_97),
.B(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_49),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_49),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_52),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_106),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_69),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_77),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_107),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_108),
.B(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_69),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_74),
.B1(n_71),
.B2(n_55),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_67),
.B1(n_55),
.B2(n_64),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_112),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_67),
.B1(n_70),
.B2(n_66),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_53),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_113),
.B(n_24),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_95),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_131),
.C(n_119),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_63),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_115),
.B(n_128),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_61),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_120),
.Y(n_141)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_121),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_80),
.B(n_82),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_63),
.B(n_59),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_57),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_129),
.Y(n_145)
);

XNOR2x1_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_94),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_56),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_82),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_130),
.B(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_21),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_31),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_110),
.B(n_63),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_137),
.C(n_148),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_123),
.A2(n_63),
.B1(n_59),
.B2(n_4),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_140),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_134),
.A2(n_122),
.B1(n_126),
.B2(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_138),
.B(n_10),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_59),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_147),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_126),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_149),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_26),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_5),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_SL g149 ( 
.A(n_132),
.B(n_20),
.C(n_46),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_154),
.C(n_157),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_153)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_32),
.C(n_45),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_43),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_47),
.C(n_44),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_8),
.B(n_9),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_145),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_168),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_171),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_34),
.C(n_41),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_175),
.C(n_147),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_150),
.B(n_12),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_174),
.B1(n_13),
.B2(n_14),
.Y(n_184)
);

XNOR2x2_ASAP7_75t_SL g172 ( 
.A(n_142),
.B(n_12),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_38),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_177),
.B(n_178),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_184),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_144),
.C(n_175),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_158),
.C(n_161),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_173),
.A2(n_143),
.B(n_141),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_173),
.B(n_179),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_166),
.A2(n_149),
.B1(n_14),
.B2(n_15),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_182),
.A2(n_169),
.B1(n_167),
.B2(n_159),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_160),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_186),
.Y(n_192)
);

INVxp67_ASAP7_75t_SL g187 ( 
.A(n_176),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_187),
.A2(n_190),
.B(n_191),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_189),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_185),
.A2(n_172),
.B(n_180),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_195),
.B(n_162),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_187),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_194),
.Y(n_199)
);

AO22x1_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_162),
.B1(n_188),
.B2(n_177),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_198),
.B(n_35),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_199),
.A2(n_200),
.B(n_36),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_201),
.B(n_37),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_16),
.Y(n_203)
);


endmodule