module real_jpeg_13432_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_345, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_345;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_2),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_168),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_2),
.A2(n_65),
.B1(n_66),
.B2(n_168),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_2),
.A2(n_58),
.B1(n_59),
.B2(n_168),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_4),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_62),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_62),
.Y(n_250)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_6),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_7),
.A2(n_45),
.B1(n_46),
.B2(n_54),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_7),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_54),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_7),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_8),
.A2(n_44),
.B1(n_65),
.B2(n_66),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_8),
.A2(n_44),
.B1(n_58),
.B2(n_59),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_44),
.Y(n_261)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_75),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_75),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_10),
.A2(n_65),
.B1(n_66),
.B2(n_75),
.Y(n_206)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_12),
.A2(n_65),
.B1(n_66),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_12),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_86),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_86),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_86),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_13),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_13),
.B(n_34),
.C(n_49),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_13),
.B(n_84),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_13),
.A2(n_119),
.B(n_172),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_13),
.A2(n_65),
.B(n_83),
.C(n_199),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_156),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_13),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_13),
.B(n_58),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_14),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_128),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_128),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_14),
.A2(n_65),
.B1(n_66),
.B2(n_128),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_20),
.B(n_342),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_17),
.B(n_343),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_18),
.A2(n_33),
.B1(n_34),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_18),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_18),
.A2(n_40),
.B1(n_65),
.B2(n_66),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_18),
.A2(n_40),
.B1(n_58),
.B2(n_59),
.Y(n_331)
);

AOI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_337),
.B(n_340),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_329),
.B(n_333),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_316),
.B(n_328),
.Y(n_22)
);

AO21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_144),
.B(n_313),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_131),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_106),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_26),
.B(n_106),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_76),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_27),
.B(n_77),
.C(n_92),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B(n_56),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_28),
.A2(n_29),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_41),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_30),
.A2(n_31),
.B1(n_56),
.B2(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_30),
.A2(n_31),
.B1(n_41),
.B2(n_42),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_37),
.B(n_38),
.Y(n_31)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_32),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_32),
.A2(n_37),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_32),
.B(n_173),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_32),
.A2(n_37),
.B1(n_118),
.B2(n_261),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_37),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_34),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_33),
.B(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_37),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_37),
.B(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_39),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_47),
.B1(n_52),
.B2(n_55),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_43),
.A2(n_47),
.B1(n_55),
.B2(n_123),
.Y(n_122)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

AO22x1_ASAP7_75t_SL g84 ( 
.A1(n_45),
.A2(n_46),
.B1(n_82),
.B2(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_45),
.B(n_160),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_46),
.A2(n_82),
.B(n_156),
.Y(n_199)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_47),
.A2(n_55),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_47),
.B(n_158),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_47),
.A2(n_55),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_47),
.A2(n_55),
.B1(n_123),
.B2(n_250),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_51),
.A2(n_53),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_51),
.A2(n_167),
.B(n_169),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_51),
.B(n_156),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_51),
.A2(n_169),
.B(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_55),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_63),
.B(n_69),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_63),
.B1(n_71),
.B2(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_59),
.B1(n_64),
.B2(n_68),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_59),
.A2(n_71),
.B(n_156),
.C(n_243),
.Y(n_242)
);

AOI32xp33_ASAP7_75t_L g256 ( 
.A1(n_59),
.A2(n_65),
.A3(n_68),
.B1(n_244),
.B2(n_257),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_63),
.B(n_74),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_63),
.A2(n_71),
.B1(n_95),
.B2(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_63),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_63),
.A2(n_69),
.B(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_63),
.A2(n_71),
.B1(n_127),
.B2(n_271),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_63)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g257 ( 
.A(n_64),
.B(n_66),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_66),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_70),
.A2(n_224),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_70),
.A2(n_224),
.B1(n_323),
.B2(n_331),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_70),
.A2(n_224),
.B(n_331),
.Y(n_339)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_71),
.A2(n_127),
.B(n_129),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_92),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_77),
.A2(n_78),
.B(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_89),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_79),
.A2(n_85),
.B1(n_87),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_79),
.A2(n_87),
.B1(n_100),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_79),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_79),
.A2(n_87),
.B1(n_219),
.B2(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_79),
.A2(n_205),
.B(n_247),
.Y(n_269)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_84),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_80),
.B(n_206),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_80),
.A2(n_84),
.B(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_84),
.B(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_87),
.A2(n_219),
.B(n_220),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_87),
.A2(n_125),
.B(n_220),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_SL g154 ( 
.A1(n_90),
.A2(n_155),
.B(n_157),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_90),
.A2(n_157),
.B(n_232),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_105),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_94),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_SL g142 ( 
.A(n_94),
.B(n_97),
.C(n_102),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_94),
.B(n_135),
.C(n_142),
.Y(n_327)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_101),
.B1(n_102),
.B2(n_104),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_102),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_102),
.B(n_136),
.C(n_140),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_112),
.C(n_113),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_107),
.A2(n_108),
.B1(n_112),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_112),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_113),
.B(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_124),
.C(n_126),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_114),
.A2(n_115),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_116),
.A2(n_121),
.B1(n_122),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_116),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_119),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_119),
.A2(n_120),
.B1(n_201),
.B2(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_119),
.A2(n_120),
.B1(n_227),
.B2(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_120),
.A2(n_178),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_120),
.B(n_156),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_120),
.A2(n_186),
.B(n_201),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_124),
.B(n_126),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_130),
.B(n_242),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_L g313 ( 
.A1(n_131),
.A2(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_143),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_132),
.B(n_143),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_142),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_137),
.Y(n_322)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_141),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_307),
.B(n_312),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_295),
.B(n_306),
.Y(n_145)
);

OAI321xp33_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_263),
.A3(n_288),
.B1(n_293),
.B2(n_294),
.C(n_345),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_236),
.B(n_262),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_213),
.B(n_235),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_194),
.B(n_212),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_174),
.B(n_193),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_161),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_152),
.B(n_161),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_159),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_153),
.A2(n_154),
.B1(n_159),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_159),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_170),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_166),
.C(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_171),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_182),
.B(n_192),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_180),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_176),
.B(n_180),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_187),
.B(n_191),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_184),
.B(n_185),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_195),
.B(n_196),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_202),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_207),
.C(n_211),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_200),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_202)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_207),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_209),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_214),
.B(n_215),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_228),
.B2(n_229),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_231),
.C(n_233),
.Y(n_237)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_222),
.C(n_226),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_233),
.B2(n_234),
.Y(n_229)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_230),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_231),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_237),
.B(n_238),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_252),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_239),
.B(n_253),
.C(n_254),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_245),
.B2(n_251),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_240),
.B(n_246),
.C(n_248),
.Y(n_277)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_245),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_259),
.Y(n_273)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_278),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_278),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_274),
.C(n_277),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_265),
.A2(n_266),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_273),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_272),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_272),
.C(n_273),
.Y(n_287)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_270),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_274),
.B(n_277),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_276),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_287),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_282),
.C(n_287),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_285),
.C(n_286),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_289),
.B(n_290),
.Y(n_293)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_305),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_305),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_300),
.C(n_301),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_309),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_327),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_327),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_326),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_321),
.B1(n_324),
.B2(n_325),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_319),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_321),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_324),
.C(n_326),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_332),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_330),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_338),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_332),
.Y(n_336)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_339),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_339),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_341),
.Y(n_340)
);


endmodule