module fake_netlist_6_1232_n_381 (n_52, n_16, n_1, n_91, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_55, n_94, n_97, n_108, n_58, n_64, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_381);

input n_52;
input n_16;
input n_1;
input n_91;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_94;
input n_97;
input n_108;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_381;

wire n_326;
wire n_256;
wire n_209;
wire n_367;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_208;
wire n_161;
wire n_316;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_297;
wire n_342;
wire n_358;
wire n_160;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_350;
wire n_142;
wire n_143;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_140;
wire n_337;
wire n_214;
wire n_246;
wire n_289;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_230;
wire n_141;
wire n_200;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_314;
wire n_378;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_360;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_344;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_371;
wire n_189;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_155;
wire n_122;
wire n_218;
wire n_234;
wire n_236;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_196;
wire n_352;
wire n_374;
wire n_366;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_293;
wire n_334;
wire n_370;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_260;
wire n_265;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_363;
wire n_323;
wire n_152;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_204;
wire n_261;
wire n_312;
wire n_130;
wire n_164;
wire n_292;
wire n_121;
wire n_307;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_237;
wire n_244;
wire n_243;
wire n_124;
wire n_282;
wire n_116;
wire n_211;
wire n_117;
wire n_175;
wire n_322;
wire n_345;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_311;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_159;
wire n_157;
wire n_162;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_221;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_277;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_317;
wire n_149;
wire n_347;
wire n_328;
wire n_373;
wire n_195;
wire n_285;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_324;
wire n_335;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_267;
wire n_339;
wire n_315;
wire n_288;
wire n_135;
wire n_165;
wire n_351;
wire n_259;
wire n_177;
wire n_364;
wire n_295;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVxp67_ASAP7_75t_SL g117 ( 
.A(n_93),
.Y(n_117)
);

INVxp33_ASAP7_75t_SL g118 ( 
.A(n_73),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_25),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_13),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_12),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_14),
.Y(n_125)
);

INVxp67_ASAP7_75t_SL g126 ( 
.A(n_79),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_18),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_23),
.Y(n_131)
);

BUFx10_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_3),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_16),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_54),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_7),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_62),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_5),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_51),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_3),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_107),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_44),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_47),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_1),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_10),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_115),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_50),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_41),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_66),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_0),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_74),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_6),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_55),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_32),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_43),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_33),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_11),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_21),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_42),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_35),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_29),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_70),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_8),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_49),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_90),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_0),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_129),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_2),
.Y(n_186)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g192 ( 
.A(n_123),
.B(n_4),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_116),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_137),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_195)
);

AND2x4_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_8),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_194),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_9),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_187),
.B(n_118),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_118),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_186),
.B(n_157),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_159),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_192),
.B(n_157),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_192),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_183),
.B(n_174),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_172),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_135),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_176),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_165),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_185),
.A2(n_195),
.B1(n_177),
.B2(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_165),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_121),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_178),
.B(n_174),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_121),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_160),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_189),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_197),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_204),
.B(n_119),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_120),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_189),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_203),
.A2(n_117),
.B(n_126),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_139),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_175),
.B1(n_171),
.B2(n_124),
.Y(n_234)
);

BUFx6f_ASAP7_75t_SL g235 ( 
.A(n_215),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_122),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_L g238 ( 
.A1(n_207),
.A2(n_170),
.B1(n_160),
.B2(n_167),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_144),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_170),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_148),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_152),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_125),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_198),
.B(n_127),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_205),
.B(n_128),
.Y(n_248)
);

AND2x4_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_130),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_SL g250 ( 
.A1(n_219),
.A2(n_168),
.B(n_166),
.C(n_164),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_198),
.B(n_131),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_224),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_134),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_138),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_140),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_202),
.B(n_142),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_218),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_154),
.B(n_146),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_145),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_228),
.A2(n_161),
.B(n_149),
.Y(n_265)
);

OAI21x1_ASAP7_75t_L g266 ( 
.A1(n_231),
.A2(n_163),
.B(n_162),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_245),
.A2(n_155),
.B(n_153),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_147),
.B(n_210),
.C(n_201),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_241),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_228),
.A2(n_9),
.B1(n_10),
.B2(n_15),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_230),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_241),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_239),
.A2(n_17),
.B(n_19),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_20),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_226),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_249),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_226),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_256),
.A2(n_22),
.B(n_24),
.C(n_26),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_249),
.Y(n_280)
);

O2A1O1Ixp5_ASAP7_75t_L g281 ( 
.A1(n_248),
.A2(n_27),
.B(n_28),
.C(n_30),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_243),
.Y(n_282)
);

AOI21x1_ASAP7_75t_L g283 ( 
.A1(n_253),
.A2(n_31),
.B(n_34),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_254),
.A2(n_36),
.B(n_37),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_236),
.A2(n_38),
.B(n_39),
.Y(n_285)
);

O2A1O1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_248),
.A2(n_40),
.B(n_45),
.C(n_46),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_261),
.B(n_242),
.C(n_263),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_L g288 ( 
.A1(n_261),
.A2(n_242),
.B(n_236),
.C(n_232),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_269),
.B(n_272),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_263),
.A2(n_236),
.B(n_229),
.C(n_234),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_260),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_238),
.Y(n_292)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_258),
.A2(n_257),
.B(n_234),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_262),
.A2(n_246),
.B(n_233),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_237),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_237),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_270),
.A2(n_275),
.B1(n_264),
.B2(n_259),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_272),
.A2(n_251),
.B1(n_247),
.B2(n_235),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_276),
.A2(n_250),
.B(n_235),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

BUFx8_ASAP7_75t_L g301 ( 
.A(n_277),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_278),
.Y(n_302)
);

AO31x2_ASAP7_75t_L g303 ( 
.A1(n_262),
.A2(n_250),
.A3(n_53),
.B(n_56),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_48),
.Y(n_304)
);

AOI31xp67_ASAP7_75t_L g305 ( 
.A1(n_266),
.A2(n_60),
.A3(n_61),
.B(n_63),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_277),
.A2(n_64),
.B(n_68),
.Y(n_306)
);

AOI21xp33_ASAP7_75t_L g307 ( 
.A1(n_273),
.A2(n_69),
.B(n_71),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_288),
.A2(n_285),
.B(n_274),
.Y(n_308)
);

NAND2x1p5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_285),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g310 ( 
.A1(n_289),
.A2(n_283),
.B(n_281),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_L g311 ( 
.A1(n_287),
.A2(n_290),
.B(n_292),
.C(n_293),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_286),
.B(n_279),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_265),
.Y(n_314)
);

AO21x2_ASAP7_75t_L g315 ( 
.A1(n_294),
.A2(n_284),
.B(n_265),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_296),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_267),
.Y(n_317)
);

AOI221xp5_ASAP7_75t_L g318 ( 
.A1(n_291),
.A2(n_284),
.B1(n_75),
.B2(n_76),
.C(n_77),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_298),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_114),
.Y(n_320)
);

OA21x2_ASAP7_75t_L g321 ( 
.A1(n_311),
.A2(n_308),
.B(n_317),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_316),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_299),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_301),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_303),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_314),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_320),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_315),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_312),
.A2(n_307),
.B(n_305),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_303),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_309),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_326),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_303),
.Y(n_334)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_306),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_327),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_309),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_325),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_325),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_323),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_322),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_328),
.B(n_310),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_340),
.B(n_321),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_338),
.B(n_321),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_336),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_321),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_328),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_321),
.Y(n_348)
);

NAND3xp33_ASAP7_75t_L g349 ( 
.A(n_331),
.B(n_318),
.C(n_330),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_329),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_329),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_327),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_336),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_330),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_347),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_335),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_345),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_352),
.B(n_348),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_332),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_354),
.B(n_332),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_357),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_360),
.B(n_345),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_358),
.B(n_346),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_362),
.B(n_355),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_363),
.B(n_361),
.Y(n_365)
);

O2A1O1Ixp5_ASAP7_75t_SL g366 ( 
.A1(n_364),
.A2(n_359),
.B(n_349),
.C(n_356),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g367 ( 
.A(n_365),
.Y(n_367)
);

AOI211xp5_ASAP7_75t_L g368 ( 
.A1(n_366),
.A2(n_349),
.B(n_363),
.C(n_344),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_R g369 ( 
.A(n_367),
.B(n_72),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_368),
.B(n_343),
.Y(n_370)
);

NAND5xp2_ASAP7_75t_L g371 ( 
.A(n_369),
.B(n_334),
.C(n_81),
.D(n_82),
.E(n_86),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_370),
.B(n_353),
.Y(n_372)
);

AND3x2_ASAP7_75t_L g373 ( 
.A(n_372),
.B(n_371),
.C(n_334),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_373),
.Y(n_374)
);

AO22x2_ASAP7_75t_L g375 ( 
.A1(n_374),
.A2(n_78),
.B1(n_88),
.B2(n_89),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_375),
.A2(n_91),
.B1(n_92),
.B2(n_95),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_375),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_376),
.A2(n_113),
.B(n_102),
.Y(n_378)
);

NAND3xp33_ASAP7_75t_L g379 ( 
.A(n_377),
.B(n_101),
.C(n_103),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_378),
.A2(n_379),
.B(n_104),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_380),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_381)
);


endmodule