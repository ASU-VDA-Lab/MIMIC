module real_jpeg_13752_n_16 (n_5, n_4, n_8, n_0, n_12, n_326, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_326;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_2),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_3),
.A2(n_49),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_3),
.A2(n_32),
.B1(n_36),
.B2(n_49),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_3),
.A2(n_49),
.B1(n_76),
.B2(n_77),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_4),
.A2(n_76),
.B1(n_77),
.B2(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_4),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_137),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_137),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_4),
.A2(n_32),
.B1(n_36),
.B2(n_137),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_6),
.A2(n_76),
.B1(n_77),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_6),
.A2(n_64),
.B1(n_65),
.B2(n_84),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_84),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_6),
.A2(n_32),
.B1(n_36),
.B2(n_84),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_7),
.A2(n_76),
.B1(n_77),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_7),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_7),
.A2(n_64),
.B1(n_65),
.B2(n_160),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_160),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_7),
.A2(n_32),
.B1(n_36),
.B2(n_160),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_10),
.A2(n_58),
.B1(n_64),
.B2(n_65),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_10),
.A2(n_32),
.B1(n_36),
.B2(n_58),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_10),
.A2(n_58),
.B1(n_76),
.B2(n_77),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_11),
.A2(n_32),
.B1(n_36),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_11),
.A2(n_40),
.B1(n_64),
.B2(n_65),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_11),
.A2(n_40),
.B1(n_46),
.B2(n_47),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_11),
.A2(n_40),
.B1(n_76),
.B2(n_77),
.Y(n_116)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_13),
.A2(n_75),
.B(n_76),
.C(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_13),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_13),
.A2(n_76),
.B1(n_77),
.B2(n_151),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_13),
.B(n_86),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_151),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_13),
.A2(n_104),
.B1(n_105),
.B2(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_13),
.B(n_92),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_14),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_14),
.A2(n_35),
.B1(n_76),
.B2(n_77),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_14),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_14),
.A2(n_35),
.B1(n_64),
.B2(n_65),
.Y(n_133)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_319),
.C(n_323),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_317),
.B(n_321),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_309),
.B(n_316),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_275),
.B(n_306),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_138),
.B(n_274),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_118),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_22),
.B(n_118),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_88),
.B2(n_117),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_23),
.B(n_89),
.C(n_101),
.Y(n_304)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_59),
.C(n_71),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_25),
.A2(n_26),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_42),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_27),
.A2(n_28),
.B1(n_42),
.B2(n_43),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_37),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_29),
.A2(n_104),
.B(n_233),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_30),
.A2(n_41),
.B1(n_128),
.B2(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_30),
.A2(n_41),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_31),
.A2(n_41),
.B(n_130),
.Y(n_204)
);

CKINVDCx6p67_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_32),
.A2(n_36),
.B1(n_52),
.B2(n_53),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_36),
.B(n_53),
.C(n_151),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_36),
.B(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_37),
.A2(n_105),
.B(n_148),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_39),
.B(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_50),
.B1(n_56),
.B2(n_57),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_45),
.A2(n_55),
.B(n_97),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

OA22x2_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_47),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_SL g200 ( 
.A1(n_46),
.A2(n_61),
.B(n_201),
.C(n_203),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_46),
.B(n_223),
.Y(n_222)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

NOR3xp33_ASAP7_75t_L g203 ( 
.A(n_47),
.B(n_62),
.C(n_64),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_50),
.A2(n_57),
.B(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_50),
.A2(n_96),
.B(n_109),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_50),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_50),
.A2(n_56),
.B1(n_208),
.B2(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_50),
.A2(n_56),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_50),
.A2(n_56),
.B1(n_216),
.B2(n_226),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_50),
.A2(n_56),
.B(n_96),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_55),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_55),
.B(n_99),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_55),
.B(n_151),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_59),
.B(n_71),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B(n_66),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_60),
.B(n_70),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_60),
.A2(n_155),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_63),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_65),
.B1(n_75),
.B2(n_80),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_64),
.A2(n_80),
.B(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

HAxp5_ASAP7_75t_SL g202 ( 
.A(n_65),
.B(n_151),
.CON(n_202),
.SN(n_202)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_66),
.B(n_156),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_67),
.A2(n_133),
.B(n_134),
.Y(n_132)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_67),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_67),
.A2(n_92),
.B1(n_154),
.B2(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_67),
.A2(n_92),
.B1(n_189),
.B2(n_202),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_67),
.A2(n_92),
.B(n_133),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_82),
.B(n_85),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_72),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_72),
.A2(n_81),
.B1(n_158),
.B2(n_161),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_72),
.A2(n_115),
.B(n_313),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_73),
.A2(n_83),
.B1(n_86),
.B2(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_73),
.A2(n_86),
.B1(n_159),
.B2(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_73),
.B(n_116),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_73),
.A2(n_86),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_73),
.A2(n_86),
.B(n_87),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_81),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_80),
.Y(n_74)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_81),
.A2(n_288),
.B(n_289),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_85),
.B(n_289),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_116),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_101),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_94),
.B(n_100),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_94),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_92),
.B(n_133),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_93),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_95),
.A2(n_206),
.B(n_207),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_100),
.B(n_278),
.C(n_291),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_100),
.B(n_278),
.CI(n_291),
.CON(n_305),
.SN(n_305)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_110),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g291 ( 
.A1(n_102),
.A2(n_103),
.B(n_112),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_103),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_107),
.B1(n_108),
.B2(n_111),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B(n_106),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_127),
.B(n_129),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_104),
.A2(n_105),
.B1(n_231),
.B2(n_239),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_105),
.B(n_151),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.C(n_124),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_119),
.A2(n_120),
.B1(n_123),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_123),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_124),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_132),
.C(n_135),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_131),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_131),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_135),
.Y(n_165)
);

INVxp33_ASAP7_75t_L g284 ( 
.A(n_134),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_268),
.B(n_273),
.Y(n_138)
);

AOI221xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_177),
.B1(n_193),
.B2(n_267),
.C(n_326),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_166),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_141),
.B(n_166),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_162),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_142),
.B(n_163),
.C(n_164),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_152),
.C(n_157),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_144),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_152),
.B(n_157),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_155),
.B(n_156),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g282 ( 
.A1(n_155),
.A2(n_283),
.B(n_284),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.C(n_176),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_176),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.C(n_174),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_172),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_191),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_178),
.B(n_191),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.C(n_183),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_179),
.B(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_181),
.B(n_183),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.C(n_187),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_187),
.B(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_266),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_261),
.B(n_265),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_217),
.B(n_260),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_212),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_197),
.B(n_212),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_209),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_205),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_199),
.B(n_205),
.C(n_209),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_200),
.B(n_204),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.C(n_215),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_215),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_255),
.B(n_259),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_245),
.B(n_254),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_234),
.B(n_244),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_229),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_224),
.B1(n_227),
.B2(n_228),
.Y(n_221)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_222),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_224),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_227),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_240),
.B(n_243),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_242),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_247),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_250),
.C(n_253),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_252),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_258),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_264),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_303),
.Y(n_275)
);

AOI21xp33_ASAP7_75t_L g306 ( 
.A1(n_276),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_292),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_292),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_287),
.B2(n_290),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_285),
.B2(n_286),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_286),
.C(n_287),
.Y(n_293)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_286),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_296),
.C(n_301),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_287),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_290),
.B1(n_295),
.B2(n_302),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_293),
.C(n_302),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_288),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_299),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_298),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_300),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_305),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_305),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_315),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_315),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_310),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_319),
.Y(n_322)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_312),
.CI(n_314),
.CON(n_310),
.SN(n_310)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_320),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);


endmodule