module fake_jpeg_16956_n_107 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_0),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_0),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_51),
.A2(n_43),
.B1(n_41),
.B2(n_40),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_58),
.B(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_47),
.B(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_57),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_50),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_32),
.B1(n_31),
.B2(n_33),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_62)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_71),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_53),
.B(n_63),
.C(n_4),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_13),
.C(n_14),
.Y(n_82)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_36),
.B1(n_3),
.B2(n_4),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_76),
.B1(n_9),
.B2(n_11),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_75),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_81),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_74),
.B(n_12),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_15),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_84),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_76),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_85),
.C(n_83),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_91),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_94),
.B1(n_77),
.B2(n_90),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_92),
.A2(n_88),
.B1(n_70),
.B2(n_79),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_98),
.C(n_93),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_99),
.C(n_20),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_18),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_103),
.A2(n_22),
.B(n_23),
.Y(n_104)
);

BUFx24_ASAP7_75t_SL g105 ( 
.A(n_104),
.Y(n_105)
);

AO21x1_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_24),
.B(n_25),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_26),
.Y(n_107)
);


endmodule