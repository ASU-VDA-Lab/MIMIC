module fake_jpeg_12521_n_174 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_9),
.B(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_7),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_31),
.B(n_32),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_13),
.B(n_0),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_41),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_19),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_24),
.B1(n_17),
.B2(n_18),
.Y(n_56)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_4),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_22),
.Y(n_43)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_15),
.B(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_16),
.B(n_6),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_4),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_24),
.Y(n_79)
);

XNOR2x1_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_74),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_26),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_69),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_26),
.Y(n_69)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_16),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_81),
.Y(n_92)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_42),
.A2(n_27),
.B1(n_20),
.B2(n_28),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_5),
.B1(n_20),
.B2(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_52),
.B(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_18),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_21),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_68),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_46),
.C(n_49),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_85),
.B(n_97),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_87),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_58),
.B1(n_65),
.B2(n_66),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_95),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_78),
.C(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_63),
.B(n_84),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_60),
.B(n_97),
.Y(n_109)
);

AO22x1_ASAP7_75t_SL g102 ( 
.A1(n_59),
.A2(n_54),
.B1(n_71),
.B2(n_64),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_103),
.Y(n_113)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_54),
.C(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_85),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_57),
.A2(n_67),
.B(n_68),
.C(n_78),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_105),
.B(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_109),
.B(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_114),
.B(n_115),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_96),
.Y(n_116)
);

NOR2x1_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_102),
.Y(n_138)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_91),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_122),
.B(n_90),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_94),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_123),
.B(n_89),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_88),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_134),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_124),
.C(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_136),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_95),
.B(n_89),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_113),
.B(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_100),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_106),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_102),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_138),
.Y(n_143)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_144),
.A2(n_132),
.B(n_129),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_129),
.C(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_109),
.C(n_112),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_130),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_125),
.B1(n_115),
.B2(n_119),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_151),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_152),
.B(n_157),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_125),
.B1(n_111),
.B2(n_137),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_155),
.B(n_156),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_144),
.A2(n_114),
.B(n_138),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_146),
.C(n_149),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_110),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_145),
.B(n_143),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_143),
.C(n_140),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_165),
.C(n_166),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_154),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_164),
.B(n_126),
.Y(n_168)
);

NAND2xp33_ASAP7_75t_SL g165 ( 
.A(n_160),
.B(n_135),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_148),
.B1(n_161),
.B2(n_118),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_168),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_108),
.C(n_118),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_108),
.C(n_120),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_170),
.C(n_120),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_120),
.Y(n_174)
);


endmodule