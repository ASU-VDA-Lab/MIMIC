module fake_jpeg_852_n_676 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_676);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_676;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_59),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_61),
.Y(n_149)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_62),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_63),
.Y(n_199)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_65),
.B(n_69),
.Y(n_160)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_68),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_70),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_10),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_72),
.B(n_76),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_74),
.Y(n_177)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_75),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_33),
.B(n_9),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_78),
.Y(n_188)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_79),
.Y(n_190)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_80),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_81),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_82),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_83),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_84),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_85),
.Y(n_187)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_87),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_35),
.B(n_9),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_107),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_89),
.Y(n_223)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_32),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_91),
.B(n_100),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_93),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_94),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_96),
.Y(n_186)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_98),
.Y(n_191)
);

BUFx4f_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g205 ( 
.A1(n_101),
.A2(n_39),
.B(n_11),
.Y(n_205)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_103),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_104),
.Y(n_194)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_106),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_40),
.B(n_18),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_108),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_26),
.Y(n_109)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_109),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_23),
.Y(n_110)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_110),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_111),
.Y(n_196)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_26),
.Y(n_112)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_35),
.B(n_9),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_115),
.Y(n_155)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_22),
.Y(n_114)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_114),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_46),
.B(n_18),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_34),
.Y(n_116)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_116),
.Y(n_220)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_38),
.Y(n_117)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_34),
.Y(n_118)
);

BUFx4f_ASAP7_75t_L g209 ( 
.A(n_118),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_34),
.Y(n_119)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_47),
.Y(n_120)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_122),
.B(n_128),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_46),
.B(n_18),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_13),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_43),
.Y(n_124)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_43),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_125),
.B(n_127),
.Y(n_182)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_126),
.Y(n_202)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_36),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_51),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_51),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_129),
.B(n_130),
.Y(n_184)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_51),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_131),
.Y(n_137)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_36),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_132),
.B(n_130),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_61),
.A2(n_50),
.B1(n_47),
.B2(n_54),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_134),
.A2(n_140),
.B1(n_152),
.B2(n_161),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_50),
.B1(n_54),
.B2(n_37),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_136),
.A2(n_143),
.B1(n_210),
.B2(n_0),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_78),
.A2(n_82),
.B1(n_70),
.B2(n_63),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_87),
.A2(n_53),
.B1(n_37),
.B2(n_41),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_99),
.B(n_56),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_145),
.B(n_159),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_83),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_147),
.B(n_180),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_63),
.A2(n_55),
.B1(n_56),
.B2(n_45),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_62),
.B(n_45),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_158),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_108),
.B(n_48),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_70),
.A2(n_55),
.B1(n_48),
.B2(n_27),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_112),
.A2(n_55),
.B1(n_53),
.B2(n_41),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_162),
.A2(n_221),
.B1(n_121),
.B2(n_119),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_89),
.A2(n_27),
.B1(n_55),
.B2(n_20),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_164),
.A2(n_74),
.B1(n_73),
.B2(n_2),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_166),
.B(n_171),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_103),
.B(n_55),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_122),
.A2(n_20),
.B1(n_29),
.B2(n_57),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_175),
.A2(n_203),
.B1(n_204),
.B2(n_228),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_75),
.B(n_12),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_178),
.B(n_192),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_116),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_92),
.A2(n_20),
.B1(n_57),
.B2(n_39),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_185),
.A2(n_6),
.B1(n_7),
.B2(n_221),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_79),
.A2(n_57),
.B(n_39),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_189),
.A2(n_84),
.B(n_81),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_80),
.B(n_9),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_95),
.B(n_131),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_197),
.B(n_198),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_96),
.B(n_14),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_59),
.A2(n_57),
.B1(n_39),
.B2(n_12),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_85),
.A2(n_57),
.B1(n_39),
.B2(n_11),
.Y(n_204)
);

HAxp5_ASAP7_75t_SL g255 ( 
.A(n_205),
.B(n_0),
.CON(n_255),
.SN(n_255)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_60),
.A2(n_8),
.B1(n_17),
.B2(n_16),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_212),
.B(n_214),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_93),
.B(n_8),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_128),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_217),
.B(n_222),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_98),
.B(n_8),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_218),
.B(n_231),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_71),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_109),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_104),
.B(n_17),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_224),
.B(n_227),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_110),
.B(n_16),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_111),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_118),
.B(n_0),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_232),
.Y(n_335)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_233),
.Y(n_318)
);

OA22x2_ASAP7_75t_L g234 ( 
.A1(n_164),
.A2(n_189),
.B1(n_169),
.B2(n_216),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_234),
.B(n_267),
.Y(n_339)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_133),
.A2(n_15),
.B(n_14),
.C(n_124),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_235),
.A2(n_304),
.B(n_247),
.C(n_244),
.Y(n_321)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_236),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_237),
.A2(n_249),
.B1(n_258),
.B2(n_296),
.Y(n_347)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_238),
.Y(n_370)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_240),
.Y(n_329)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_242),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_165),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_243),
.B(n_248),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_244),
.A2(n_249),
.B(n_253),
.Y(n_357)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_245),
.Y(n_348)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_246),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_158),
.B(n_0),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_247),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_182),
.Y(n_248)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_250),
.Y(n_354)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_135),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_252),
.B(n_254),
.Y(n_333)
);

AOI32xp33_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_15),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_255),
.A2(n_211),
.B(n_167),
.Y(n_320)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_170),
.Y(n_256)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_256),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_162),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_259),
.A2(n_301),
.B1(n_307),
.B2(n_309),
.Y(n_322)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_170),
.Y(n_260)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_260),
.Y(n_331)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_138),
.Y(n_261)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_261),
.Y(n_336)
);

INVx6_ASAP7_75t_SL g262 ( 
.A(n_150),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g372 ( 
.A(n_262),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_160),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_263),
.B(n_287),
.Y(n_353)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_181),
.Y(n_264)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_264),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_213),
.B(n_146),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_265),
.Y(n_332)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_200),
.Y(n_266)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_266),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_168),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_184),
.Y(n_269)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_144),
.B(n_1),
.CI(n_3),
.CON(n_270),
.SN(n_270)
);

FAx1_ASAP7_75t_SL g342 ( 
.A(n_270),
.B(n_177),
.CI(n_193),
.CON(n_342),
.SN(n_342)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_200),
.Y(n_272)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_272),
.Y(n_334)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_220),
.Y(n_273)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_273),
.Y(n_337)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_169),
.Y(n_274)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_274),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_197),
.B(n_3),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_277),
.B(n_279),
.Y(n_330)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_220),
.Y(n_278)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_278),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_155),
.B(n_3),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_139),
.B(n_4),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_281),
.B(n_285),
.Y(n_344)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_195),
.Y(n_282)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_282),
.Y(n_364)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_174),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_283),
.Y(n_361)
);

OR2x2_ASAP7_75t_SL g284 ( 
.A(n_168),
.B(n_6),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_284),
.B(n_308),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_139),
.B(n_148),
.Y(n_285)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_195),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_213),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_288),
.B(n_292),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_289),
.B(n_290),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_213),
.B(n_156),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_146),
.B(n_156),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_291),
.B(n_298),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_176),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_154),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_293),
.B(n_294),
.Y(n_359)
);

AOI32xp33_ASAP7_75t_L g294 ( 
.A1(n_229),
.A2(n_196),
.A3(n_225),
.B1(n_148),
.B2(n_157),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_137),
.A2(n_163),
.B1(n_201),
.B2(n_209),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_295),
.A2(n_305),
.B1(n_315),
.B2(n_138),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_179),
.A2(n_208),
.B1(n_206),
.B2(n_223),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_181),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_297),
.B(n_299),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_174),
.B(n_216),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_179),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_202),
.B(n_153),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_300),
.B(n_193),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_229),
.A2(n_188),
.B1(n_149),
.B2(n_208),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_206),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_302),
.B(n_310),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_215),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_303),
.B(n_306),
.Y(n_378)
);

A2O1A1Ixp33_ASAP7_75t_L g304 ( 
.A1(n_196),
.A2(n_215),
.B(n_230),
.C(n_194),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_209),
.A2(n_219),
.B1(n_223),
.B2(n_142),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_209),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_141),
.A2(n_191),
.B1(n_186),
.B2(n_151),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_149),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_188),
.A2(n_230),
.B1(n_194),
.B2(n_225),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_190),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_172),
.B(n_187),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_311),
.B(n_312),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_172),
.B(n_187),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_190),
.B(n_207),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_313),
.B(n_316),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_141),
.A2(n_186),
.B1(n_191),
.B2(n_151),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_207),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_317),
.A2(n_303),
.B1(n_233),
.B2(n_240),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_320),
.A2(n_352),
.B(n_298),
.Y(n_387)
);

O2A1O1Ixp33_ASAP7_75t_L g397 ( 
.A1(n_321),
.A2(n_246),
.B(n_242),
.C(n_236),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_237),
.A2(n_289),
.B1(n_268),
.B2(n_275),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_338),
.A2(n_351),
.B1(n_368),
.B2(n_374),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_269),
.A2(n_142),
.B1(n_167),
.B2(n_177),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_340),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_275),
.B(n_268),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_341),
.B(n_349),
.C(n_358),
.Y(n_382)
);

OR2x2_ASAP7_75t_SL g404 ( 
.A(n_342),
.B(n_358),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_346),
.B(n_291),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_211),
.C(n_276),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_277),
.B(n_281),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_350),
.B(n_270),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_286),
.A2(n_251),
.B1(n_239),
.B2(n_234),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_247),
.A2(n_235),
.B(n_271),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_357),
.A2(n_373),
.B(n_320),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_314),
.B(n_285),
.C(n_265),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_241),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_328),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_307),
.A2(n_262),
.B1(n_310),
.B2(n_316),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_365),
.Y(n_412)
);

MAJx2_ASAP7_75t_L g366 ( 
.A(n_279),
.B(n_255),
.C(n_265),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_366),
.B(n_367),
.C(n_371),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_234),
.A2(n_257),
.B1(n_290),
.B2(n_295),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_304),
.A2(n_234),
.B(n_284),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_290),
.A2(n_270),
.B1(n_280),
.B2(n_261),
.Y(n_374)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_369),
.Y(n_379)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_379),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_380),
.B(n_383),
.Y(n_443)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_369),
.Y(n_381)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_381),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_357),
.A2(n_291),
.B1(n_298),
.B2(n_283),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_384),
.A2(n_389),
.B1(n_394),
.B2(n_396),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_385),
.B(n_406),
.Y(n_463)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_355),
.Y(n_386)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_386),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_387),
.A2(n_401),
.B(n_334),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_341),
.B(n_274),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_388),
.B(n_390),
.C(n_407),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_373),
.A2(n_260),
.B1(n_256),
.B2(n_266),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_SL g390 ( 
.A(n_351),
.B(n_308),
.C(n_299),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_360),
.B(n_302),
.Y(n_391)
);

NOR3xp33_ASAP7_75t_L g452 ( 
.A(n_391),
.B(n_420),
.C(n_378),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_350),
.B(n_278),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_392),
.B(n_395),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_347),
.A2(n_272),
.B1(n_273),
.B2(n_287),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_344),
.B(n_330),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_347),
.A2(n_238),
.B1(n_282),
.B2(n_293),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_397),
.A2(n_375),
.B(n_353),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_359),
.A2(n_306),
.B1(n_264),
.B2(n_267),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_398),
.A2(n_424),
.B1(n_425),
.B2(n_372),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_399),
.A2(n_402),
.B1(n_409),
.B2(n_426),
.Y(n_459)
);

INVx5_ASAP7_75t_L g400 ( 
.A(n_329),
.Y(n_400)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_400),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_338),
.A2(n_297),
.B1(n_250),
.B2(n_245),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_344),
.B(n_232),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_403),
.B(n_404),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_330),
.B(n_374),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_405),
.B(n_411),
.Y(n_456)
);

FAx1_ASAP7_75t_SL g406 ( 
.A(n_366),
.B(n_352),
.CI(n_349),
.CON(n_406),
.SN(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_366),
.B(n_376),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_328),
.B(n_326),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_408),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_368),
.A2(n_339),
.B1(n_359),
.B2(n_371),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_355),
.Y(n_410)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_410),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_343),
.B(n_376),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_318),
.Y(n_413)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_413),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_372),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_414),
.B(n_416),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_343),
.B(n_346),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_318),
.Y(n_417)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_417),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_326),
.B(n_353),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_418),
.Y(n_453)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_319),
.Y(n_419)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_419),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_321),
.B(n_367),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_378),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_428),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_422),
.B(n_327),
.Y(n_433)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_329),
.Y(n_423)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_423),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_339),
.A2(n_371),
.B1(n_367),
.B2(n_342),
.Y(n_424)
);

OAI22xp33_ASAP7_75t_L g425 ( 
.A1(n_322),
.A2(n_339),
.B1(n_332),
.B2(n_342),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_317),
.A2(n_333),
.B1(n_327),
.B2(n_356),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_336),
.Y(n_427)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_427),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_335),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_382),
.B(n_356),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_432),
.B(n_433),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_435),
.A2(n_441),
.B(n_464),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_436),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_401),
.A2(n_363),
.B(n_333),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_437),
.A2(n_422),
.B(n_384),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_SL g441 ( 
.A1(n_415),
.A2(n_354),
.B1(n_348),
.B2(n_370),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_382),
.B(n_375),
.C(n_361),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_444),
.B(n_448),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_398),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_450),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_407),
.B(n_375),
.C(n_319),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_400),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_420),
.A2(n_378),
.B(n_363),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_451),
.A2(n_462),
.B(n_397),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_452),
.B(n_457),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_423),
.Y(n_457)
);

OA21x2_ASAP7_75t_L g462 ( 
.A1(n_393),
.A2(n_324),
.B(n_325),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_SL g464 ( 
.A1(n_412),
.A2(n_354),
.B1(n_348),
.B2(n_370),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_393),
.A2(n_336),
.B1(n_324),
.B2(n_325),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_465),
.A2(n_394),
.B1(n_396),
.B2(n_417),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_466),
.A2(n_411),
.B(n_416),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_388),
.B(n_334),
.C(n_362),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_467),
.B(n_323),
.Y(n_509)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_386),
.Y(n_469)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_469),
.Y(n_478)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_410),
.Y(n_470)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_470),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g541 ( 
.A1(n_471),
.A2(n_475),
.B(n_480),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_462),
.Y(n_474)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_474),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_466),
.A2(n_387),
.B(n_412),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_435),
.A2(n_409),
.B1(n_405),
.B2(n_426),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_476),
.A2(n_493),
.B1(n_496),
.B2(n_498),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_446),
.B(n_395),
.Y(n_477)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_477),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_451),
.A2(n_424),
.B(n_421),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_446),
.B(n_392),
.Y(n_482)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_482),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_429),
.B(n_381),
.Y(n_484)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_484),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_485),
.A2(n_492),
.B(n_439),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_456),
.B(n_383),
.Y(n_486)
);

INVxp33_ASAP7_75t_L g521 ( 
.A(n_486),
.Y(n_521)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_434),
.Y(n_488)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_488),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_489),
.A2(n_495),
.B1(n_500),
.B2(n_507),
.Y(n_519)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_434),
.Y(n_491)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_491),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_447),
.A2(n_402),
.B1(n_390),
.B2(n_403),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_445),
.Y(n_494)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_494),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_459),
.A2(n_389),
.B1(n_379),
.B2(n_391),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_456),
.A2(n_404),
.B1(n_406),
.B2(n_380),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_429),
.B(n_413),
.Y(n_497)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_497),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_437),
.A2(n_406),
.B1(n_414),
.B2(n_419),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_445),
.Y(n_499)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_499),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_459),
.A2(n_428),
.B1(n_427),
.B2(n_370),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_440),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_501),
.B(n_502),
.Y(n_516)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_455),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_453),
.B(n_427),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_503),
.B(n_508),
.Y(n_535)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_455),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_504),
.B(n_505),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_430),
.B(n_362),
.Y(n_505)
);

FAx1_ASAP7_75t_SL g506 ( 
.A(n_436),
.B(n_335),
.CI(n_337),
.CON(n_506),
.SN(n_506)
);

FAx1_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_451),
.CI(n_483),
.CON(n_512),
.SN(n_512)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_462),
.A2(n_364),
.B1(n_337),
.B2(n_345),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_430),
.B(n_364),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_509),
.B(n_467),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_474),
.A2(n_449),
.B1(n_454),
.B2(n_443),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_510),
.A2(n_511),
.B1(n_513),
.B2(n_518),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_495),
.A2(n_449),
.B1(n_454),
.B2(n_443),
.Y(n_511)
);

NOR2x1p5_ASAP7_75t_L g567 ( 
.A(n_512),
.B(n_483),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_471),
.A2(n_462),
.B1(n_431),
.B2(n_463),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_514),
.B(n_539),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_490),
.B(n_444),
.C(n_487),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_517),
.B(n_529),
.C(n_538),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_471),
.A2(n_431),
.B1(n_463),
.B2(n_465),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_476),
.A2(n_438),
.B1(n_432),
.B2(n_433),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_520),
.A2(n_528),
.B1(n_542),
.B2(n_475),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_490),
.B(n_438),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_SL g549 ( 
.A(n_522),
.B(n_496),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_503),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_525),
.B(n_473),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_501),
.B(n_486),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_526),
.B(n_530),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_472),
.A2(n_470),
.B1(n_469),
.B2(n_460),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_490),
.B(n_448),
.C(n_458),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_473),
.B(n_345),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_497),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_534),
.B(n_484),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_487),
.B(n_460),
.C(n_458),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_472),
.A2(n_439),
.B1(n_457),
.B2(n_450),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_498),
.B(n_442),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_543),
.B(n_508),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_480),
.A2(n_468),
.B1(n_442),
.B2(n_461),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_544),
.A2(n_493),
.B1(n_507),
.B2(n_500),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_492),
.B(n_461),
.C(n_331),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_546),
.B(n_529),
.C(n_517),
.Y(n_557)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_548),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_549),
.B(n_557),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_537),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_550),
.B(n_554),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_516),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_551),
.B(n_576),
.Y(n_587)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_537),
.Y(n_552)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_552),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_516),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_515),
.A2(n_480),
.B1(n_475),
.B2(n_477),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_556),
.A2(n_513),
.B1(n_518),
.B2(n_510),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_558),
.A2(n_575),
.B1(n_540),
.B2(n_512),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_534),
.B(n_505),
.Y(n_559)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_559),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_522),
.B(n_509),
.C(n_485),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_560),
.B(n_563),
.C(n_572),
.Y(n_584)
);

XOR2x2_ASAP7_75t_L g600 ( 
.A(n_561),
.B(n_569),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_562),
.B(n_536),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_538),
.B(n_482),
.C(n_504),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g564 ( 
.A(n_535),
.Y(n_564)
);

INVx13_ASAP7_75t_L g589 ( 
.A(n_564),
.Y(n_589)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_531),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_566),
.B(n_567),
.Y(n_582)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_531),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_568),
.B(n_570),
.Y(n_588)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_532),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_SL g571 ( 
.A(n_520),
.B(n_483),
.Y(n_571)
);

OAI322xp33_ASAP7_75t_L g594 ( 
.A1(n_571),
.A2(n_512),
.A3(n_524),
.B1(n_527),
.B2(n_541),
.C1(n_515),
.C2(n_506),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_514),
.B(n_491),
.C(n_502),
.Y(n_572)
);

CKINVDCx16_ASAP7_75t_R g573 ( 
.A(n_528),
.Y(n_573)
);

BUFx12_ASAP7_75t_L g580 ( 
.A(n_573),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_546),
.B(n_479),
.C(n_499),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_574),
.B(n_577),
.C(n_488),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_519),
.A2(n_489),
.B1(n_506),
.B2(n_479),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_521),
.B(n_335),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_543),
.B(n_478),
.C(n_494),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_578),
.A2(n_585),
.B1(n_597),
.B2(n_598),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_574),
.B(n_542),
.Y(n_583)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_583),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_554),
.A2(n_511),
.B1(n_523),
.B2(n_540),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_586),
.B(n_591),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_557),
.B(n_539),
.C(n_541),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_593),
.A2(n_575),
.B1(n_558),
.B2(n_570),
.Y(n_616)
);

XOR2x2_ASAP7_75t_L g611 ( 
.A(n_594),
.B(n_569),
.Y(n_611)
);

AOI322xp5_ASAP7_75t_SL g595 ( 
.A1(n_565),
.A2(n_524),
.A3(n_527),
.B1(n_506),
.B2(n_481),
.C1(n_533),
.C2(n_536),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_SL g618 ( 
.A(n_595),
.B(n_377),
.Y(n_618)
);

A2O1A1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_567),
.A2(n_523),
.B(n_544),
.C(n_545),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_596),
.B(n_548),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_556),
.A2(n_481),
.B1(n_545),
.B2(n_532),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_547),
.B(n_533),
.C(n_478),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_601),
.B(n_547),
.C(n_586),
.Y(n_603)
);

FAx1_ASAP7_75t_L g602 ( 
.A(n_567),
.B(n_468),
.CI(n_331),
.CON(n_602),
.SN(n_602)
);

A2O1A1Ixp33_ASAP7_75t_SL g614 ( 
.A1(n_602),
.A2(n_568),
.B(n_566),
.C(n_552),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_603),
.B(n_611),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_601),
.B(n_572),
.C(n_553),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_604),
.B(n_608),
.C(n_612),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_605),
.B(n_607),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_582),
.B(n_559),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_584),
.B(n_553),
.C(n_560),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_582),
.A2(n_550),
.B(n_555),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_609),
.A2(n_602),
.B(n_596),
.Y(n_625)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_598),
.Y(n_610)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_610),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_584),
.B(n_577),
.C(n_563),
.Y(n_612)
);

NOR2xp67_ASAP7_75t_L g613 ( 
.A(n_591),
.B(n_571),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_613),
.B(n_614),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_600),
.B(n_555),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_615),
.B(n_583),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_616),
.A2(n_593),
.B1(n_602),
.B2(n_581),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_600),
.B(n_549),
.C(n_323),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_617),
.B(n_622),
.C(n_599),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_618),
.B(n_621),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_587),
.B(n_377),
.Y(n_619)
);

CKINVDCx16_ASAP7_75t_R g629 ( 
.A(n_619),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_578),
.A2(n_585),
.B1(n_592),
.B2(n_581),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_583),
.B(n_590),
.C(n_597),
.Y(n_622)
);

INVx6_ASAP7_75t_L g624 ( 
.A(n_620),
.Y(n_624)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_624),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_625),
.A2(n_633),
.B(n_614),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_628),
.B(n_623),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_SL g633 ( 
.A(n_605),
.B(n_579),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_607),
.B(n_588),
.Y(n_635)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_635),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_636),
.A2(n_616),
.B1(n_617),
.B2(n_580),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_614),
.B(n_588),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_637),
.B(n_638),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_603),
.B(n_590),
.C(n_579),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_639),
.B(n_640),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_614),
.B(n_592),
.Y(n_640)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_641),
.Y(n_655)
);

XOR2xp5_ASAP7_75t_L g657 ( 
.A(n_644),
.B(n_649),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_630),
.B(n_612),
.C(n_604),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_645),
.B(n_648),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_633),
.A2(n_606),
.B(n_623),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_L g660 ( 
.A1(n_646),
.A2(n_625),
.B(n_626),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_SL g648 ( 
.A(n_630),
.B(n_608),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_639),
.B(n_622),
.C(n_615),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_629),
.B(n_609),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_651),
.A2(n_653),
.B(n_634),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_SL g654 ( 
.A(n_652),
.B(n_631),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_638),
.B(n_611),
.C(n_580),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_654),
.B(n_661),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_656),
.A2(n_658),
.B(n_660),
.Y(n_667)
);

O2A1O1Ixp33_ASAP7_75t_SL g658 ( 
.A1(n_643),
.A2(n_627),
.B(n_626),
.C(n_631),
.Y(n_658)
);

OAI21xp33_ASAP7_75t_L g661 ( 
.A1(n_653),
.A2(n_632),
.B(n_627),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g662 ( 
.A1(n_650),
.A2(n_632),
.B(n_637),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_662),
.B(n_635),
.Y(n_668)
);

AO221x1_ASAP7_75t_L g664 ( 
.A1(n_659),
.A2(n_624),
.B1(n_636),
.B2(n_642),
.C(n_645),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_SL g670 ( 
.A1(n_664),
.A2(n_644),
.B(n_580),
.Y(n_670)
);

XOR2xp5_ASAP7_75t_L g665 ( 
.A(n_657),
.B(n_649),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_665),
.B(n_666),
.Y(n_671)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_659),
.B(n_647),
.C(n_646),
.Y(n_666)
);

OAI21xp33_ASAP7_75t_SL g669 ( 
.A1(n_668),
.A2(n_640),
.B(n_655),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_L g673 ( 
.A(n_669),
.B(n_670),
.C(n_628),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_671),
.A2(n_667),
.B1(n_666),
.B2(n_663),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g674 ( 
.A(n_672),
.B(n_673),
.C(n_665),
.Y(n_674)
);

XOR2xp5_ASAP7_75t_L g675 ( 
.A(n_674),
.B(n_589),
.Y(n_675)
);

XNOR2xp5_ASAP7_75t_L g676 ( 
.A(n_675),
.B(n_589),
.Y(n_676)
);


endmodule