module fake_jpeg_31483_n_196 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_196);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_196;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx2_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx12f_ASAP7_75t_SL g35 ( 
.A(n_22),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_49),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_13),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_38),
.B(n_41),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_1),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_44),
.B(n_54),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_20),
.B(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_61),
.Y(n_67)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_57),
.Y(n_96)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_15),
.B(n_2),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

CKINVDCx6p67_ASAP7_75t_R g94 ( 
.A(n_62),
.Y(n_94)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_40),
.A2(n_30),
.B1(n_25),
.B2(n_23),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_70),
.A2(n_97),
.B1(n_45),
.B2(n_50),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_99),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_36),
.B(n_18),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_25),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_2),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_54),
.B(n_7),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_64),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_9),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_33),
.A2(n_6),
.B1(n_3),
.B2(n_5),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_6),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_54),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_102),
.B(n_103),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_55),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_62),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_108),
.Y(n_130)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_62),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_74),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_84),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_114),
.Y(n_138)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_52),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_99),
.C(n_97),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_115),
.A2(n_98),
.B1(n_82),
.B2(n_65),
.Y(n_129)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_32),
.B1(n_68),
.B2(n_88),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_117),
.B(n_78),
.Y(n_124)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_85),
.Y(n_123)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_64),
.B(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_121),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_124),
.B1(n_129),
.B2(n_135),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_76),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_104),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_87),
.B(n_74),
.C(n_75),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_119),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_71),
.B1(n_69),
.B2(n_93),
.Y(n_135)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_100),
.B1(n_120),
.B2(n_110),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_152),
.B1(n_133),
.B2(n_126),
.Y(n_164)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_147),
.Y(n_160)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_100),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_101),
.B(n_138),
.C(n_124),
.D(n_136),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_128),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_150),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_101),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_151),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_100),
.B1(n_107),
.B2(n_116),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_125),
.C(n_130),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_157),
.C(n_163),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_104),
.C(n_137),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_152),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_136),
.C(n_135),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_164),
.B(n_141),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_141),
.B1(n_142),
.B2(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_166),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_162),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_169),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_170),
.A2(n_171),
.B(n_172),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_158),
.A2(n_129),
.B1(n_150),
.B2(n_134),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_156),
.C(n_161),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_178),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_168),
.A2(n_150),
.B(n_153),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_173),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_180),
.A2(n_181),
.B(n_183),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_158),
.B(n_172),
.Y(n_181)
);

OA21x2_ASAP7_75t_SL g182 ( 
.A1(n_174),
.A2(n_170),
.B(n_159),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_176),
.Y(n_186)
);

XOR2x2_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_132),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_186),
.B(n_187),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_143),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_140),
.Y(n_188)
);

AOI31xp67_ASAP7_75t_SL g191 ( 
.A1(n_188),
.A2(n_109),
.A3(n_73),
.B(n_72),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_185),
.A2(n_105),
.B(n_112),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_81),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_192),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_189),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_193),
.Y(n_196)
);


endmodule