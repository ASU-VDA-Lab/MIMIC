module fake_jpeg_8304_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_35),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_28),
.B1(n_36),
.B2(n_47),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_30),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_28),
.B1(n_36),
.B2(n_47),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_55),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_17),
.B1(n_22),
.B2(n_32),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_71),
.B1(n_72),
.B2(n_31),
.Y(n_101)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_60),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_10),
.Y(n_110)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_65),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_27),
.B1(n_32),
.B2(n_22),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_74),
.Y(n_91)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

OR2x2_ASAP7_75t_SL g100 ( 
.A(n_70),
.B(n_44),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_17),
.B1(n_29),
.B2(n_18),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_29),
.B1(n_18),
.B2(n_20),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_34),
.B1(n_43),
.B2(n_39),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_80),
.A2(n_114),
.B1(n_120),
.B2(n_33),
.Y(n_129)
);

OAI32xp33_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_43),
.A3(n_34),
.B1(n_48),
.B2(n_21),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_81),
.A2(n_51),
.B1(n_73),
.B2(n_19),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_86),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_64),
.A2(n_30),
.B1(n_24),
.B2(n_21),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_84),
.A2(n_101),
.B1(n_110),
.B2(n_33),
.Y(n_133)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g132 ( 
.A(n_87),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_89),
.B(n_99),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_48),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_90),
.B(n_112),
.C(n_119),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_92),
.A2(n_97),
.B1(n_118),
.B2(n_0),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_93),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_55),
.A2(n_21),
.B1(n_24),
.B2(n_19),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_61),
.A2(n_26),
.B1(n_24),
.B2(n_42),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_100),
.A2(n_0),
.B(n_1),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_42),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_42),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_44),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_69),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_116),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_44),
.C(n_45),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_75),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_113),
.A2(n_76),
.B1(n_33),
.B2(n_9),
.Y(n_125)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_65),
.B(n_19),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_66),
.A2(n_26),
.B1(n_19),
.B2(n_33),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_66),
.B(n_45),
.C(n_51),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_121),
.A2(n_137),
.B1(n_147),
.B2(n_95),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_81),
.A2(n_73),
.B1(n_45),
.B2(n_76),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_124),
.A2(n_130),
.B1(n_102),
.B2(n_103),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_33),
.B1(n_16),
.B2(n_14),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_133),
.A2(n_117),
.B1(n_93),
.B2(n_99),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_104),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_148),
.B1(n_102),
.B2(n_120),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_79),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_116),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_145),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_92),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_90),
.A2(n_11),
.B1(n_10),
.B2(n_2),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_98),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_100),
.B(n_88),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_107),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_159),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_156),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_112),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_155),
.A2(n_152),
.B(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_164),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_119),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_147),
.C(n_130),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_131),
.B(n_108),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_108),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_170),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_180),
.B1(n_183),
.B2(n_184),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_126),
.B(n_110),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_163),
.B(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_126),
.B(n_110),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_141),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_122),
.B(n_138),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_167),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_169),
.A2(n_178),
.B(n_182),
.Y(n_185)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_140),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_172),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_132),
.B1(n_139),
.B2(n_150),
.Y(n_199)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_175),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_122),
.A2(n_111),
.B(n_85),
.C(n_118),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_114),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_177),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_148),
.B(n_97),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_124),
.A2(n_85),
.B1(n_96),
.B2(n_109),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_87),
.Y(n_181)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_143),
.B(n_1),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_137),
.A2(n_121),
.B1(n_133),
.B2(n_127),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_186),
.B(n_201),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_188),
.A2(n_161),
.B1(n_177),
.B2(n_178),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_169),
.A2(n_129),
.B(n_136),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_SL g239 ( 
.A(n_190),
.B(n_212),
.C(n_4),
.Y(n_239)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_193),
.B(n_200),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_198),
.C(n_201),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_168),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_205),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_199),
.A2(n_157),
.B1(n_156),
.B2(n_173),
.Y(n_222)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_132),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_210),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_160),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_162),
.A2(n_135),
.B1(n_123),
.B2(n_134),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_207),
.A2(n_182),
.B1(n_153),
.B2(n_179),
.Y(n_225)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_154),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_211),
.Y(n_228)
);

A2O1A1O1Ixp25_ASAP7_75t_L g212 ( 
.A1(n_155),
.A2(n_82),
.B(n_135),
.C(n_123),
.D(n_134),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_155),
.B(n_149),
.C(n_139),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_149),
.C(n_3),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_175),
.A2(n_149),
.B1(n_139),
.B2(n_86),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_235)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_175),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_217),
.A2(n_170),
.B(n_164),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_222),
.B1(n_235),
.B2(n_244),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_220),
.A2(n_242),
.B(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_223),
.Y(n_256)
);

FAx1_ASAP7_75t_SL g223 ( 
.A(n_213),
.B(n_166),
.CI(n_167),
.CON(n_223),
.SN(n_223)
);

OAI32xp33_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_183),
.A3(n_165),
.B1(n_163),
.B2(n_174),
.Y(n_224)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_227),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_232),
.C(n_236),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

OA21x2_ASAP7_75t_SL g231 ( 
.A1(n_186),
.A2(n_179),
.B(n_180),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_185),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_2),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_233),
.A2(n_239),
.B(n_189),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_4),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_213),
.A2(n_188),
.B1(n_187),
.B2(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_4),
.C(n_5),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_241),
.C(n_189),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_5),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_192),
.B(n_5),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_187),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_185),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_254),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_248),
.A2(n_257),
.B(n_263),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_245),
.A2(n_208),
.B1(n_215),
.B2(n_194),
.Y(n_251)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_238),
.A2(n_191),
.B1(n_202),
.B2(n_192),
.Y(n_252)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_200),
.B1(n_209),
.B2(n_210),
.Y(n_253)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_220),
.A2(n_224),
.B1(n_219),
.B2(n_237),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_255),
.A2(n_223),
.B1(n_226),
.B2(n_235),
.Y(n_272)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_228),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_219),
.B(n_212),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_264),
.C(n_232),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_191),
.C(n_193),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_241),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_274),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_258),
.A2(n_221),
.B1(n_227),
.B2(n_199),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_271),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_272),
.B(n_247),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_234),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_252),
.B(n_203),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_286),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_240),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_280),
.Y(n_298)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_279),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_256),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_223),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_282),
.C(n_283),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_225),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_228),
.C(n_211),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_262),
.B(n_251),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_195),
.Y(n_288)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_273),
.A2(n_267),
.B1(n_261),
.B2(n_259),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_290),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_313)
);

OAI21x1_ASAP7_75t_L g291 ( 
.A1(n_269),
.A2(n_257),
.B(n_263),
.Y(n_291)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_297),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_250),
.B(n_265),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_294),
.A2(n_199),
.B(n_203),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_SL g297 ( 
.A1(n_281),
.A2(n_266),
.A3(n_248),
.B1(n_233),
.B2(n_264),
.C1(n_199),
.C2(n_242),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_242),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_301),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_195),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_283),
.C(n_271),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_304),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_285),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_294),
.B(n_289),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_307),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_282),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_310),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_290),
.A2(n_280),
.B(n_268),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_295),
.A2(n_268),
.B(n_277),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_300),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_313),
.B(n_7),
.Y(n_316)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_315),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_319),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_300),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_310),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_298),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_306),
.B(n_298),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_322),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_287),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_SL g325 ( 
.A(n_318),
.B(n_314),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_328),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_320),
.A2(n_305),
.B1(n_311),
.B2(n_303),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_326),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_324),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_332),
.C(n_309),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_302),
.C(n_318),
.Y(n_332)
);

INVx11_ASAP7_75t_L g333 ( 
.A(n_331),
.Y(n_333)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_333),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_329),
.B(n_333),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_334),
.B(n_333),
.Y(n_337)
);

AOI322xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_334),
.A3(n_333),
.B1(n_314),
.B2(n_307),
.C1(n_287),
.C2(n_8),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_334),
.Y(n_339)
);


endmodule