module fake_jpeg_20532_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx6_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_9),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_3),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_20),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_24),
.Y(n_29)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_1),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_27),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_35),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_21),
.A2(n_19),
.B(n_14),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_11),
.B(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_13),
.Y(n_45)
);

FAx1_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_16),
.CI(n_14),
.CON(n_42),
.SN(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_12),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_25),
.B1(n_23),
.B2(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_17),
.B1(n_26),
.B2(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_26),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_43),
.C(n_7),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_45),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_8),
.B1(n_5),
.B2(n_6),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_38),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_42),
.Y(n_54)
);

NAND3xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_7),
.C(n_8),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_54),
.B1(n_55),
.B2(n_47),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_59),
.A2(n_60),
.B1(n_39),
.B2(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_52),
.C(n_53),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_64),
.C(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_66),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_56),
.C(n_40),
.Y(n_66)
);

BUFx24_ASAP7_75t_SL g67 ( 
.A(n_63),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_67),
.B(n_62),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

MAJx2_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_64),
.C(n_43),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_43),
.B(n_49),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_70),
.Y(n_73)
);


endmodule