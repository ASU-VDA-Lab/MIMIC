module real_jpeg_1712_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_286;
wire n_176;
wire n_166;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_1),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_83),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_83),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_1),
.A2(n_59),
.B1(n_63),
.B2(n_83),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_2),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_176),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_176),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_2),
.A2(n_59),
.B1(n_63),
.B2(n_176),
.Y(n_286)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_3),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_4),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_122),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_122),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_4),
.A2(n_59),
.B1(n_63),
.B2(n_122),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_5),
.A2(n_25),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_5),
.B(n_25),
.Y(n_29)
);

AO22x2_ASAP7_75t_L g30 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_5),
.A2(n_11),
.B(n_25),
.C(n_225),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_7),
.A2(n_37),
.B1(n_59),
.B2(n_63),
.Y(n_114)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_10),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_144),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_144),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_10),
.A2(n_59),
.B1(n_63),
.B2(n_144),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_11),
.B(n_41),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_11),
.B(n_52),
.Y(n_213)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_11),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_11),
.B(n_30),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_226),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_11),
.B(n_59),
.C(n_62),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_226),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_11),
.B(n_112),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_11),
.B(n_57),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_51),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_12),
.A2(n_51),
.B1(n_59),
.B2(n_63),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_43),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_13),
.A2(n_43),
.B1(n_59),
.B2(n_63),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_15),
.A2(n_41),
.B1(n_42),
.B2(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_15),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_75),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_75),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_15),
.A2(n_59),
.B1(n_63),
.B2(n_75),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_89),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_88),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_21),
.B(n_76),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_55),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_38),
.B1(n_53),
.B2(n_54),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_35),
.Y(n_23)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_24),
.B(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_24),
.A2(n_30),
.B1(n_193),
.B2(n_210),
.Y(n_238)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_25),
.A2(n_26),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

AOI32xp33_ASAP7_75t_L g196 ( 
.A1(n_25),
.A2(n_42),
.A3(n_46),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g198 ( 
.A(n_26),
.B(n_47),
.Y(n_198)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_30),
.B(n_173),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_31),
.A2(n_32),
.B1(n_61),
.B2(n_62),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_31),
.A2(n_34),
.B(n_226),
.Y(n_225)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_32),
.B(n_271),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_36),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_50),
.B2(n_52),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_45),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_42),
.A2(n_73),
.B(n_226),
.C(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_44),
.B(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_44),
.A2(n_52),
.B1(n_143),
.B2(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_73),
.B1(n_74),
.B2(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_45),
.A2(n_82),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_45),
.B(n_121),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_45),
.A2(n_119),
.B(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_68),
.C(n_72),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_68),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g84 ( 
.A(n_56),
.B(n_81),
.C(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_64),
.B(n_66),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_57),
.A2(n_64),
.B1(n_117),
.B2(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_57),
.A2(n_64),
.B1(n_138),
.B2(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_57),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_67),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_58),
.A2(n_98),
.B1(n_99),
.B2(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_58),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_58),
.A2(n_242),
.B(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_58),
.A2(n_98),
.B1(n_219),
.B2(n_253),
.Y(n_264)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_59),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_59),
.B(n_282),
.Y(n_281)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_64),
.A2(n_218),
.B(n_220),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_64),
.B(n_222),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_71),
.B1(n_87),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_69),
.A2(n_71),
.B1(n_96),
.B2(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_69),
.A2(n_192),
.B(n_194),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_69),
.A2(n_194),
.B(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_71),
.A2(n_140),
.B(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_71),
.A2(n_172),
.B(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_73),
.A2(n_142),
.B(n_145),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.C(n_84),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_77),
.A2(n_81),
.B1(n_101),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_81),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_84),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_152),
.B(n_323),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_147),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_123),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_92),
.B(n_123),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_104),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_95),
.B(n_97),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_94),
.B(n_100),
.C(n_104),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_98),
.A2(n_221),
.B(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B(n_118),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_106),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_115),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_108),
.B1(n_118),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_107),
.A2(n_108),
.B1(n_115),
.B2(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_112),
.B(n_113),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_109),
.A2(n_112),
.B1(n_135),
.B2(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_109),
.A2(n_226),
.B(n_259),
.Y(n_283)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_110),
.A2(n_111),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_110),
.A2(n_111),
.B1(n_201),
.B2(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_110),
.B(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_110),
.A2(n_257),
.B(n_258),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_110),
.A2(n_111),
.B1(n_257),
.B2(n_291),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_111),
.A2(n_216),
.B(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_111),
.B(n_230),
.Y(n_259)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_112),
.A2(n_229),
.B(n_286),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_115),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.C(n_130),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_125),
.B1(n_129),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_139),
.C(n_141),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_132),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_133),
.A2(n_136),
.B1(n_137),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_141),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_146),
.B(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_147),
.A2(n_324),
.B(n_325),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_148),
.B(n_151),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_177),
.B(n_322),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_154),
.B(n_157),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.C(n_163),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_170),
.C(n_174),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_165),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_166),
.B(n_168),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_167),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_169),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_171),
.B1(n_174),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

OAI21x1_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_203),
.B(n_321),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_179),
.B(n_181),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.C(n_188),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_182),
.B(n_186),
.Y(n_306)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_188),
.B(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.C(n_195),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_189),
.B(n_191),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_195),
.B(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_196),
.A2(n_199),
.B1(n_200),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_196),
.Y(n_245)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI31xp33_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_303),
.A3(n_313),
.B(n_318),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_247),
.B(n_302),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_231),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_206),
.B(n_231),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_217),
.C(n_223),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_207),
.B(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_212),
.C(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_217),
.B(n_223),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_224),
.B(n_227),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_243),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_232),
.B(n_244),
.C(n_246),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_233),
.B(n_238),
.C(n_239),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_297),
.B(n_301),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_266),
.B(n_296),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_260),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_250),
.B(n_260),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.C(n_255),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_256),
.B1(n_275),
.B2(n_277),
.Y(n_274)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_265),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_264),
.C(n_265),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_278),
.B(n_295),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_274),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_274),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_269),
.A2(n_270),
.B1(n_272),
.B2(n_293),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_275),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_289),
.B(n_294),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_284),
.B(n_288),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_287),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_286),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_292),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_300),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_307),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_310),
.C(n_311),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_315),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_317),
.Y(n_319)
);


endmodule