module fake_jpeg_29999_n_436 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_436);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_436;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

INVx8_ASAP7_75t_SL g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_47),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_44),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_65),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_55),
.B(n_87),
.Y(n_126)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_0),
.B(n_1),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_62),
.B(n_1),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_68),
.Y(n_118)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_21),
.B(n_15),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_69),
.B(n_83),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVxp67_ASAP7_75t_SL g91 ( 
.A(n_74),
.Y(n_91)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_82),
.Y(n_92)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_39),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_85),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_86),
.Y(n_123)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_37),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_51),
.A2(n_33),
.B1(n_32),
.B2(n_37),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_108),
.A2(n_83),
.B1(n_87),
.B2(n_75),
.Y(n_159)
);

AND2x4_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_33),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_131),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_132),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_81),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_45),
.A2(n_39),
.B1(n_42),
.B2(n_21),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_122),
.B1(n_31),
.B2(n_24),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_49),
.A2(n_39),
.B1(n_42),
.B2(n_26),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_41),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_58),
.B(n_26),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_80),
.B(n_39),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_134),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_72),
.B(n_36),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_144),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_143),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_113),
.A2(n_25),
.B1(n_112),
.B2(n_31),
.Y(n_144)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_31),
.C(n_36),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_157),
.Y(n_178)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_147),
.Y(n_195)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_148),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_108),
.A2(n_88),
.B1(n_64),
.B2(n_66),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_150),
.B1(n_159),
.B2(n_104),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_73),
.B1(n_63),
.B2(n_79),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_125),
.B(n_38),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_167),
.Y(n_179)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_118),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_160),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_94),
.B(n_24),
.Y(n_160)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_163),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_101),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_175),
.B1(n_128),
.B2(n_136),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_100),
.A2(n_77),
.B1(n_70),
.B2(n_38),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_135),
.B1(n_130),
.B2(n_109),
.Y(n_199)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_95),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_171),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_41),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_174),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_173),
.A2(n_99),
.B1(n_128),
.B2(n_97),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_93),
.B(n_81),
.Y(n_174)
);

AND2x6_ASAP7_75t_L g175 ( 
.A(n_112),
.B(n_59),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_189),
.A2(n_191),
.B1(n_176),
.B2(n_196),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_123),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_190),
.B(n_198),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_164),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_147),
.A2(n_115),
.B1(n_96),
.B2(n_93),
.Y(n_197)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_140),
.B(n_169),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_130),
.B1(n_109),
.B2(n_102),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_140),
.B(n_135),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_202),
.B(n_141),
.Y(n_223)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_205),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_178),
.B(n_155),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_222),
.Y(n_231)
);

AND2x6_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_175),
.Y(n_207)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_155),
.C(n_169),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g240 ( 
.A1(n_209),
.A2(n_206),
.B(n_212),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_189),
.A2(n_149),
.B1(n_150),
.B2(n_144),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_217),
.B(n_220),
.Y(n_233)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_211),
.Y(n_236)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_202),
.C(n_179),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_181),
.C(n_184),
.Y(n_241)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_215),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_191),
.A2(n_164),
.B(n_151),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_218),
.A2(n_226),
.B1(n_142),
.B2(n_120),
.Y(n_250)
);

OA21x2_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_170),
.B(n_168),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_228),
.B1(n_196),
.B2(n_186),
.Y(n_235)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_225),
.Y(n_232)
);

INVx13_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_227),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_157),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_191),
.A2(n_106),
.B1(n_103),
.B2(n_97),
.Y(n_226)
);

INVx13_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_178),
.B(n_166),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_229),
.B(n_182),
.Y(n_254)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_235),
.A2(n_242),
.B1(n_252),
.B2(n_226),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_179),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_246),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_217),
.C(n_209),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_223),
.A2(n_186),
.B1(n_183),
.B2(n_148),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_216),
.A2(n_195),
.B1(n_187),
.B2(n_177),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_243),
.A2(n_187),
.B1(n_230),
.B2(n_177),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_181),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_184),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_249),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_200),
.B(n_195),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_248),
.A2(n_255),
.B(n_220),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_185),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_250),
.A2(n_216),
.B1(n_230),
.B2(n_204),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_210),
.A2(n_143),
.B1(n_153),
.B2(n_187),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_163),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_254),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_185),
.B(n_182),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_205),
.B(n_213),
.Y(n_256)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_256),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_256),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_258),
.B(n_264),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_257),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_259),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_260),
.B(n_241),
.C(n_246),
.Y(n_296)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_257),
.Y(n_261)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_229),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_265),
.A2(n_274),
.B1(n_283),
.B2(n_251),
.Y(n_311)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_266),
.Y(n_297)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_267),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_269),
.A2(n_277),
.B(n_278),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_254),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_270),
.Y(n_313)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_220),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_272),
.B(n_282),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_253),
.A2(n_219),
.B1(n_220),
.B2(n_210),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_275),
.B(n_239),
.Y(n_303)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_276),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_233),
.A2(n_216),
.B(n_207),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_207),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_154),
.Y(n_309)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_280),
.B(n_286),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_284),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_180),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_252),
.A2(n_208),
.B1(n_222),
.B2(n_218),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_245),
.Y(n_284)
);

AND2x6_ASAP7_75t_L g285 ( 
.A(n_234),
.B(n_233),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_285),
.A2(n_288),
.B(n_236),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_239),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_255),
.A2(n_204),
.B(n_180),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_275),
.B(n_288),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_291),
.A2(n_292),
.B(n_306),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_234),
.B(n_235),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_232),
.B(n_249),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_293),
.A2(n_303),
.B(n_312),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_300),
.C(n_308),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_232),
.C(n_242),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_270),
.B(n_245),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_203),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_285),
.A2(n_243),
.B(n_236),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_263),
.A2(n_262),
.B1(n_286),
.B2(n_273),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_265),
.B1(n_263),
.B2(n_283),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_260),
.B(n_250),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_310),
.C(n_315),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_268),
.B(n_215),
.C(n_211),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_311),
.A2(n_273),
.B1(n_271),
.B2(n_267),
.Y(n_323)
);

AOI221xp5_ASAP7_75t_L g314 ( 
.A1(n_262),
.A2(n_236),
.B1(n_251),
.B2(n_167),
.C(n_158),
.Y(n_314)
);

OAI21xp33_ASAP7_75t_L g325 ( 
.A1(n_314),
.A2(n_259),
.B(n_280),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_204),
.C(n_171),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_317),
.A2(n_321),
.B1(n_322),
.B2(n_334),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_304),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_324),
.Y(n_354)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_320),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_292),
.A2(n_284),
.B1(n_266),
.B2(n_276),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_306),
.A2(n_307),
.B1(n_291),
.B2(n_303),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_323),
.A2(n_327),
.B1(n_332),
.B2(n_289),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_259),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_295),
.Y(n_345)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_326),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_311),
.A2(n_261),
.B1(n_203),
.B2(n_173),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_301),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_333),
.Y(n_359)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_331),
.Y(n_356)
);

NOR2x1_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_227),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_297),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_297),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_295),
.A2(n_138),
.B1(n_145),
.B2(n_161),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_335),
.A2(n_336),
.B1(n_340),
.B2(n_290),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_313),
.B(n_14),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_296),
.B(n_139),
.C(n_162),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_338),
.B(n_310),
.C(n_315),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_142),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_339),
.B(n_301),
.Y(n_347)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_302),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_341),
.B(n_345),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_319),
.B(n_329),
.C(n_338),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_342),
.B(n_346),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_319),
.B(n_309),
.Y(n_346)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_347),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_329),
.B(n_300),
.C(n_308),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_348),
.B(n_349),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_312),
.C(n_298),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_350),
.A2(n_326),
.B1(n_334),
.B2(n_333),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_298),
.C(n_293),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_352),
.B(n_353),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_322),
.B(n_289),
.C(n_302),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_321),
.B(n_305),
.C(n_294),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_355),
.B(n_362),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_357),
.A2(n_224),
.B1(n_136),
.B2(n_107),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_317),
.B(n_305),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_358),
.Y(n_364)
);

NOR3xp33_ASAP7_75t_SL g360 ( 
.A(n_336),
.B(n_339),
.C(n_337),
.Y(n_360)
);

NOR3xp33_ASAP7_75t_SL g363 ( 
.A(n_360),
.B(n_331),
.C(n_337),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_327),
.A2(n_290),
.B1(n_294),
.B2(n_173),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_361),
.B(n_152),
.Y(n_376)
);

FAx1_ASAP7_75t_SL g362 ( 
.A(n_323),
.B(n_91),
.CI(n_227),
.CON(n_362),
.SN(n_362)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_363),
.A2(n_371),
.B1(n_376),
.B2(n_362),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_349),
.A2(n_332),
.B(n_320),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_367),
.A2(n_352),
.B(n_351),
.Y(n_385)
);

INVx13_ASAP7_75t_L g368 ( 
.A(n_360),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_368),
.B(n_375),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_354),
.Y(n_370)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_370),
.Y(n_384)
);

NOR3xp33_ASAP7_75t_SL g371 ( 
.A(n_359),
.B(n_318),
.C(n_330),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_355),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_353),
.A2(n_340),
.B1(n_152),
.B2(n_96),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_373),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_347),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_379),
.A2(n_103),
.B1(n_97),
.B2(n_106),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_343),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_91),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_341),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_387),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_342),
.C(n_348),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_393),
.C(n_373),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_363),
.A2(n_344),
.B1(n_356),
.B2(n_345),
.Y(n_383)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_383),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_386),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_372),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_379),
.A2(n_107),
.B1(n_106),
.B2(n_103),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_391),
.B(n_394),
.Y(n_404)
);

BUFx24_ASAP7_75t_SL g392 ( 
.A(n_368),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_392),
.B(n_378),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_224),
.C(n_137),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_389),
.A2(n_371),
.B1(n_367),
.B2(n_376),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_395),
.B(n_396),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_378),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_400),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_402),
.B(n_403),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_386),
.B(n_364),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_393),
.A2(n_369),
.B(n_374),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_405),
.B(n_406),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_381),
.B(n_15),
.Y(n_406)
);

A2O1A1Ixp33_ASAP7_75t_SL g407 ( 
.A1(n_402),
.A2(n_388),
.B(n_398),
.C(n_401),
.Y(n_407)
);

AOI322xp5_ASAP7_75t_L g420 ( 
.A1(n_407),
.A2(n_14),
.A3(n_2),
.B1(n_3),
.B2(n_5),
.C1(n_6),
.C2(n_1),
.Y(n_420)
);

INVx11_ASAP7_75t_L g409 ( 
.A(n_404),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_409),
.A2(n_11),
.B(n_2),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_397),
.A2(n_388),
.B1(n_384),
.B2(n_390),
.Y(n_411)
);

AOI322xp5_ASAP7_75t_L g419 ( 
.A1(n_411),
.A2(n_27),
.A3(n_14),
.B1(n_117),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_419)
);

INVx6_ASAP7_75t_L g412 ( 
.A(n_401),
.Y(n_412)
);

AOI322xp5_ASAP7_75t_L g423 ( 
.A1(n_412),
.A2(n_410),
.A3(n_411),
.B1(n_407),
.B2(n_413),
.C1(n_6),
.C2(n_7),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_400),
.A2(n_90),
.B1(n_27),
.B2(n_99),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_414),
.B(n_416),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_86),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_85),
.C(n_82),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_417),
.B(n_418),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_415),
.B(n_27),
.C(n_117),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_419),
.B(n_420),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_422),
.B(n_423),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_420),
.A2(n_410),
.B(n_407),
.Y(n_426)
);

AOI322xp5_ASAP7_75t_L g431 ( 
.A1(n_426),
.A2(n_5),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.C1(n_11),
.C2(n_428),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_421),
.B(n_1),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_427),
.B(n_2),
.C(n_3),
.Y(n_430)
);

A2O1A1Ixp33_ASAP7_75t_L g429 ( 
.A1(n_424),
.A2(n_2),
.B(n_3),
.C(n_5),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_429),
.A2(n_430),
.B(n_431),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_432),
.A2(n_425),
.B(n_8),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_433),
.B(n_7),
.C(n_8),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_434),
.B(n_10),
.C(n_11),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_435),
.B(n_11),
.Y(n_436)
);


endmodule