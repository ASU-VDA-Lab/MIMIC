module real_aes_14853_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_92;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_87;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
OA21x2_ASAP7_75t_L g93 ( .A1(n_0), .A2(n_43), .B(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g176 ( .A(n_0), .Y(n_176) );
INVx1_ASAP7_75t_L g596 ( .A(n_1), .Y(n_596) );
AND2x2_ASAP7_75t_L g129 ( .A(n_2), .B(n_130), .Y(n_129) );
AOI221xp5_ASAP7_75t_L g168 ( .A1(n_3), .A2(n_75), .B1(n_153), .B2(n_169), .C(n_170), .Y(n_168) );
BUFx3_ASAP7_75t_L g522 ( .A(n_4), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_5), .B(n_136), .Y(n_258) );
INVx3_ASAP7_75t_L g605 ( .A(n_6), .Y(n_605) );
INVx1_ASAP7_75t_L g573 ( .A(n_7), .Y(n_573) );
INVx2_ASAP7_75t_L g528 ( .A(n_8), .Y(n_528) );
INVx1_ASAP7_75t_L g539 ( .A(n_8), .Y(n_539) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_9), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_10), .B(n_98), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_11), .B(n_248), .Y(n_247) );
BUFx3_ASAP7_75t_L g100 ( .A(n_12), .Y(n_100) );
INVx1_ASAP7_75t_L g111 ( .A(n_12), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_13), .B(n_113), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g718 ( .A(n_14), .Y(n_718) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_15), .Y(n_205) );
BUFx10_ASAP7_75t_L g731 ( .A(n_16), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_17), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g749 ( .A(n_17), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_18), .B(n_121), .Y(n_202) );
OAI21xp33_ASAP7_75t_L g286 ( .A1(n_18), .A2(n_59), .B(n_287), .Y(n_286) );
O2A1O1Ixp5_ASAP7_75t_L g171 ( .A1(n_19), .A2(n_158), .B(n_160), .C(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g618 ( .A(n_20), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g641 ( .A(n_20), .B(n_29), .Y(n_641) );
INVxp33_ASAP7_75t_L g659 ( .A(n_20), .Y(n_659) );
INVx1_ASAP7_75t_L g690 ( .A(n_20), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_21), .A2(n_55), .B1(n_560), .B2(n_561), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_21), .A2(n_44), .B1(n_669), .B2(n_671), .Y(n_668) );
INVx1_ASAP7_75t_L g119 ( .A(n_22), .Y(n_119) );
INVx2_ASAP7_75t_L g615 ( .A(n_23), .Y(n_615) );
INVxp67_ASAP7_75t_SL g546 ( .A(n_24), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_24), .A2(n_32), .B1(n_680), .B2(n_683), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_25), .B(n_103), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_26), .A2(n_57), .B1(n_575), .B2(n_578), .Y(n_574) );
INVxp67_ASAP7_75t_L g667 ( .A(n_26), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_27), .B(n_150), .Y(n_149) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_27), .Y(n_737) );
XOR2xp5_ASAP7_75t_L g512 ( .A(n_28), .B(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g619 ( .A(n_29), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_29), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g707 ( .A(n_30), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_31), .B(n_113), .Y(n_112) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_32), .A2(n_49), .B1(n_517), .B2(n_529), .Y(n_516) );
INVx1_ASAP7_75t_L g589 ( .A(n_33), .Y(n_589) );
OAI222xp33_ASAP7_75t_L g636 ( .A1(n_33), .A2(n_49), .B1(n_74), .B2(n_637), .C1(n_642), .C2(n_645), .Y(n_636) );
AND2x4_ASAP7_75t_L g118 ( .A(n_34), .B(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_34), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g563 ( .A1(n_35), .A2(n_564), .B(n_567), .Y(n_563) );
INVxp33_ASAP7_75t_L g627 ( .A(n_35), .Y(n_627) );
NAND2x1_ASAP7_75t_L g257 ( .A(n_36), .B(n_130), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_37), .Y(n_212) );
INVx1_ASAP7_75t_L g253 ( .A(n_38), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_38), .A2(n_253), .B1(n_714), .B2(n_715), .Y(n_713) );
INVx1_ASAP7_75t_L g527 ( .A(n_39), .Y(n_527) );
INVx1_ASAP7_75t_L g538 ( .A(n_39), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_40), .Y(n_226) );
AND2x2_ASAP7_75t_L g128 ( .A(n_41), .B(n_109), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_42), .B(n_102), .Y(n_187) );
INVx1_ASAP7_75t_L g175 ( .A(n_43), .Y(n_175) );
AOI21xp33_ASAP7_75t_L g579 ( .A1(n_44), .A2(n_580), .B(n_582), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_45), .B(n_136), .Y(n_236) );
INVx1_ASAP7_75t_L g94 ( .A(n_46), .Y(n_94) );
BUFx2_ASAP7_75t_L g714 ( .A(n_47), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_48), .B(n_109), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_50), .B(n_121), .Y(n_198) );
OAI22xp33_ASAP7_75t_L g534 ( .A1(n_51), .A2(n_74), .B1(n_535), .B2(n_540), .Y(n_534) );
INVx1_ASAP7_75t_L g676 ( .A(n_51), .Y(n_676) );
INVx1_ASAP7_75t_L g555 ( .A(n_52), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_53), .B(n_190), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g101 ( .A(n_54), .B(n_102), .Y(n_101) );
INVxp67_ASAP7_75t_SL g663 ( .A(n_55), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_56), .B(n_231), .Y(n_230) );
INVxp33_ASAP7_75t_L g609 ( .A(n_57), .Y(n_609) );
AND2x2_ASAP7_75t_L g135 ( .A(n_58), .B(n_136), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_59), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_60), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g97 ( .A(n_61), .B(n_98), .Y(n_97) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_62), .B(n_102), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_63), .Y(n_173) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_63), .A2(n_173), .B1(n_710), .B2(n_711), .Y(n_709) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_64), .B(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_65), .B(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_66), .B(n_122), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g108 ( .A(n_67), .B(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g717 ( .A(n_68), .Y(n_717) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_69), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_70), .B(n_152), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_71), .B(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g106 ( .A(n_72), .Y(n_106) );
BUFx3_ASAP7_75t_L g116 ( .A(n_72), .Y(n_116) );
INVx1_ASAP7_75t_L g133 ( .A(n_72), .Y(n_133) );
INVx2_ASAP7_75t_L g616 ( .A(n_73), .Y(n_616) );
INVxp67_ASAP7_75t_SL g630 ( .A(n_73), .Y(n_630) );
AND2x2_ASAP7_75t_L g635 ( .A(n_73), .B(n_615), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_76), .B(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g521 ( .A(n_77), .Y(n_521) );
AOI21xp33_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_500), .B(n_511), .Y(n_78) );
INVx4_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
AND2x4_ASAP7_75t_L g80 ( .A(n_81), .B(n_381), .Y(n_80) );
NOR4xp75_ASAP7_75t_L g81 ( .A(n_82), .B(n_303), .C(n_334), .D(n_362), .Y(n_81) );
OAI211xp5_ASAP7_75t_SL g82 ( .A1(n_83), .A2(n_163), .B(n_237), .C(n_267), .Y(n_82) );
INVxp67_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
AND2x2_ASAP7_75t_L g84 ( .A(n_85), .B(n_124), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_86), .B(n_440), .Y(n_458) );
NOR2xp67_ASAP7_75t_L g492 ( .A(n_86), .B(n_296), .Y(n_492) );
INVx1_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g238 ( .A(n_87), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g278 ( .A(n_87), .Y(n_278) );
INVx1_ASAP7_75t_L g299 ( .A(n_87), .Y(n_299) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_87), .Y(n_310) );
AND2x2_ASAP7_75t_L g406 ( .A(n_87), .B(n_407), .Y(n_406) );
INVx3_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g323 ( .A(n_88), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g379 ( .A(n_88), .B(n_297), .Y(n_379) );
AND2x2_ASAP7_75t_L g430 ( .A(n_88), .B(n_241), .Y(n_430) );
BUFx3_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g332 ( .A(n_89), .Y(n_332) );
OAI21x1_ASAP7_75t_L g89 ( .A1(n_90), .A2(n_95), .B(n_120), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
BUFx3_ASAP7_75t_L g287 ( .A(n_92), .Y(n_287) );
BUFx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g123 ( .A(n_93), .Y(n_123) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_93), .Y(n_136) );
INVx1_ASAP7_75t_L g177 ( .A(n_94), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g95 ( .A1(n_96), .A2(n_107), .B(n_117), .Y(n_95) );
AOI21xp5_ASAP7_75t_L g96 ( .A1(n_97), .A2(n_101), .B(n_104), .Y(n_96) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_99), .B(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g213 ( .A(n_99), .Y(n_213) );
INVx1_ASAP7_75t_L g223 ( .A(n_99), .Y(n_223) );
INVx2_ASAP7_75t_L g232 ( .A(n_99), .Y(n_232) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx2_ASAP7_75t_L g103 ( .A(n_100), .Y(n_103) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_100), .Y(n_114) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g150 ( .A(n_103), .Y(n_150) );
INVx2_ASAP7_75t_L g190 ( .A(n_103), .Y(n_190) );
INVx2_ASAP7_75t_L g207 ( .A(n_103), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_104), .A2(n_149), .B(n_151), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_104), .A2(n_193), .B(n_195), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_104), .A2(n_230), .B(n_233), .Y(n_229) );
BUFx10_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx3_ASAP7_75t_L g170 ( .A(n_106), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_112), .B(n_115), .Y(n_107) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g158 ( .A(n_110), .Y(n_158) );
INVx2_ASAP7_75t_L g211 ( .A(n_110), .Y(n_211) );
INVx1_ASAP7_75t_L g254 ( .A(n_110), .Y(n_254) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g154 ( .A(n_111), .Y(n_154) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx3_ASAP7_75t_L g130 ( .A(n_114), .Y(n_130) );
INVx3_ASAP7_75t_L g250 ( .A(n_114), .Y(n_250) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g209 ( .A(n_116), .Y(n_209) );
INVx2_ASAP7_75t_L g248 ( .A(n_116), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_116), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g162 ( .A(n_117), .Y(n_162) );
OAI21x1_ASAP7_75t_L g245 ( .A1(n_117), .A2(n_246), .B(n_255), .Y(n_245) );
BUFx6f_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx3_ASAP7_75t_L g144 ( .A(n_118), .Y(n_144) );
INVx2_ASAP7_75t_L g197 ( .A(n_118), .Y(n_197) );
INVx1_ASAP7_75t_L g217 ( .A(n_118), .Y(n_217) );
INVx1_ASAP7_75t_L g505 ( .A(n_118), .Y(n_505) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_119), .Y(n_699) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_122), .B(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g396 ( .A(n_124), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g325 ( .A(n_125), .Y(n_325) );
INVx2_ASAP7_75t_L g333 ( .A(n_125), .Y(n_333) );
AND2x2_ASAP7_75t_L g429 ( .A(n_125), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g483 ( .A(n_125), .Y(n_483) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_145), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_126), .B(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_126), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g293 ( .A(n_126), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g297 ( .A(n_126), .Y(n_297) );
INVx2_ASAP7_75t_L g313 ( .A(n_126), .Y(n_313) );
AO21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_134), .B(n_141), .Y(n_126) );
OAI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_129), .B(n_131), .Y(n_127) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
BUFx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g160 ( .A(n_133), .Y(n_160) );
NOR2xp67_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
AOI21xp33_ASAP7_75t_L g141 ( .A1(n_135), .A2(n_142), .B(n_143), .Y(n_141) );
INVxp33_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
INVx1_ASAP7_75t_L g180 ( .A(n_136), .Y(n_180) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_136), .Y(n_184) );
INVx1_ASAP7_75t_L g244 ( .A(n_136), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_139), .B(n_140), .Y(n_137) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NOR3xp33_ASAP7_75t_L g167 ( .A(n_144), .B(n_168), .C(n_171), .Y(n_167) );
INVx3_ASAP7_75t_L g294 ( .A(n_145), .Y(n_294) );
INVx1_ASAP7_75t_L g308 ( .A(n_145), .Y(n_308) );
AND2x2_ASAP7_75t_L g312 ( .A(n_145), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g407 ( .A(n_145), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g434 ( .A(n_145), .Y(n_434) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
OAI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_155), .B(n_161), .Y(n_147) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx3_ASAP7_75t_L g169 ( .A(n_154), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_159), .Y(n_155) );
INVx2_ASAP7_75t_L g510 ( .A(n_158), .Y(n_510) );
AOI21x1_ASAP7_75t_L g255 ( .A1(n_159), .A2(n_256), .B(n_257), .Y(n_255) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g191 ( .A(n_160), .Y(n_191) );
INVx2_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
AOI32xp33_ASAP7_75t_L g355 ( .A1(n_164), .A2(n_356), .A3(n_358), .B1(n_359), .B2(n_361), .Y(n_355) );
AND2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_199), .Y(n_164) );
INVx1_ASAP7_75t_L g339 ( .A(n_165), .Y(n_339) );
AND2x2_ASAP7_75t_L g444 ( .A(n_165), .B(n_262), .Y(n_444) );
AND2x2_ASAP7_75t_L g497 ( .A(n_165), .B(n_271), .Y(n_497) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_181), .Y(n_165) );
INVx2_ASAP7_75t_L g266 ( .A(n_166), .Y(n_266) );
AND2x2_ASAP7_75t_L g269 ( .A(n_166), .B(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_166), .Y(n_466) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_174), .B(n_178), .Y(n_166) );
NAND2xp33_ASAP7_75t_L g288 ( .A(n_167), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g194 ( .A(n_169), .Y(n_194) );
INVx1_ASAP7_75t_L g215 ( .A(n_170), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_170), .A2(n_222), .B1(n_224), .B2(n_228), .Y(n_221) );
INVx2_ASAP7_75t_SL g227 ( .A(n_170), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_170), .B(n_508), .Y(n_507) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_177), .Y(n_174) );
AOI21x1_ASAP7_75t_L g218 ( .A1(n_175), .A2(n_176), .B(n_177), .Y(n_218) );
NOR2xp33_ASAP7_75t_R g178 ( .A(n_179), .B(n_180), .Y(n_178) );
INVx2_ASAP7_75t_L g265 ( .A(n_181), .Y(n_265) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVxp67_ASAP7_75t_L g390 ( .A(n_182), .Y(n_390) );
OAI21x1_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_185), .B(n_198), .Y(n_182) );
OAI21x1_ASAP7_75t_L g219 ( .A1(n_183), .A2(n_220), .B(n_236), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_183), .A2(n_185), .B(n_198), .Y(n_270) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_183), .A2(n_220), .B(n_236), .Y(n_284) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
OAI21x1_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_192), .B(n_196), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_191), .Y(n_186) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx2_ASAP7_75t_SL g235 ( .A(n_197), .Y(n_235) );
AND2x2_ASAP7_75t_L g375 ( .A(n_199), .B(n_376), .Y(n_375) );
NAND2x1p5_ASAP7_75t_L g413 ( .A(n_199), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g435 ( .A(n_199), .B(n_269), .Y(n_435) );
AND2x4_ASAP7_75t_SL g451 ( .A(n_199), .B(n_264), .Y(n_451) );
AND2x2_ASAP7_75t_L g472 ( .A(n_199), .B(n_301), .Y(n_472) );
AND2x4_ASAP7_75t_L g199 ( .A(n_200), .B(n_219), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g263 ( .A(n_201), .Y(n_263) );
INVx2_ASAP7_75t_L g272 ( .A(n_201), .Y(n_272) );
AND2x2_ASAP7_75t_L g327 ( .A(n_201), .B(n_219), .Y(n_327) );
AND2x2_ASAP7_75t_L g354 ( .A(n_201), .B(n_319), .Y(n_354) );
AND2x4_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
NAND3xp33_ASAP7_75t_L g285 ( .A(n_203), .B(n_286), .C(n_288), .Y(n_285) );
NAND3xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_210), .C(n_216), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_208), .C(n_209), .Y(n_204) );
INVx2_ASAP7_75t_SL g206 ( .A(n_207), .Y(n_206) );
OAI221xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B1(n_213), .B2(n_214), .C(n_215), .Y(n_210) );
INVx2_ASAP7_75t_L g234 ( .A(n_211), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g290 ( .A(n_218), .Y(n_290) );
INVx1_ASAP7_75t_L g273 ( .A(n_219), .Y(n_273) );
OAI21x1_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_229), .B(n_235), .Y(n_220) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_259), .Y(n_237) );
INVxp67_ASAP7_75t_SL g431 ( .A(n_238), .Y(n_431) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g352 ( .A(n_240), .Y(n_352) );
INVx1_ASAP7_75t_L g277 ( .A(n_241), .Y(n_277) );
INVx2_ASAP7_75t_L g324 ( .A(n_241), .Y(n_324) );
INVx1_ASAP7_75t_L g349 ( .A(n_241), .Y(n_349) );
AND2x2_ASAP7_75t_L g361 ( .A(n_241), .B(n_332), .Y(n_361) );
AND2x4_ASAP7_75t_SL g367 ( .A(n_241), .B(n_313), .Y(n_367) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_241), .Y(n_371) );
INVxp67_ASAP7_75t_L g408 ( .A(n_241), .Y(n_408) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_245), .B(n_258), .Y(n_242) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_249), .B(n_251), .Y(n_246) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OAI22xp33_ASAP7_75t_L g455 ( .A1(n_260), .A2(n_456), .B1(n_458), .B2(n_459), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_262), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_262), .B(n_338), .Y(n_479) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g342 ( .A(n_264), .Y(n_342) );
AND2x2_ASAP7_75t_L g380 ( .A(n_264), .B(n_271), .Y(n_380) );
AND2x2_ASAP7_75t_L g499 ( .A(n_264), .B(n_283), .Y(n_499) );
AND2x4_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g280 ( .A(n_265), .Y(n_280) );
AND2x2_ASAP7_75t_L g301 ( .A(n_266), .B(n_302), .Y(n_301) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_266), .Y(n_485) );
AOI222xp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_274), .B1(n_279), .B2(n_291), .C1(n_295), .C2(n_300), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
AND2x2_ASAP7_75t_L g326 ( .A(n_269), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g353 ( .A(n_269), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g358 ( .A(n_269), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_269), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g460 ( .A(n_269), .B(n_404), .Y(n_460) );
INVx1_ASAP7_75t_L g302 ( .A(n_270), .Y(n_302) );
AND2x2_ASAP7_75t_L g343 ( .A(n_271), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_271), .B(n_329), .Y(n_427) );
AND2x2_ASAP7_75t_L g490 ( .A(n_271), .B(n_301), .Y(n_490) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g404 ( .A(n_272), .Y(n_404) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g463 ( .A(n_275), .B(n_341), .Y(n_463) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_277), .Y(n_397) );
NOR2x1p5_ASAP7_75t_SL g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g414 ( .A(n_280), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_280), .B(n_354), .Y(n_469) );
OAI221xp5_ASAP7_75t_L g426 ( .A1(n_281), .A2(n_427), .B1(n_428), .B2(n_431), .C(n_432), .Y(n_426) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_285), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_283), .B(n_299), .Y(n_298) );
INVxp67_ASAP7_75t_SL g401 ( .A(n_283), .Y(n_401) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_283), .Y(n_412) );
OR2x2_ASAP7_75t_L g480 ( .A(n_283), .B(n_285), .Y(n_480) );
BUFx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g319 ( .A(n_284), .Y(n_319) );
INVx1_ASAP7_75t_L g391 ( .A(n_285), .Y(n_391) );
INVx1_ASAP7_75t_L g421 ( .A(n_285), .Y(n_421) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR3xp33_ASAP7_75t_L g304 ( .A(n_291), .B(n_305), .C(n_311), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_291), .A2(n_337), .B1(n_340), .B2(n_342), .Y(n_336) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g369 ( .A(n_293), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_293), .B(n_373), .Y(n_411) );
AND2x2_ASAP7_75t_L g424 ( .A(n_293), .B(n_344), .Y(n_424) );
OR2x2_ASAP7_75t_L g296 ( .A(n_294), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g341 ( .A(n_294), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx3_ASAP7_75t_L g440 ( .A(n_296), .Y(n_440) );
INVx1_ASAP7_75t_L g373 ( .A(n_299), .Y(n_373) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x4_ASAP7_75t_L g317 ( .A(n_301), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_301), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g329 ( .A(n_302), .Y(n_329) );
OAI21xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_314), .B(n_320), .Y(n_303) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g365 ( .A(n_307), .B(n_366), .Y(n_365) );
AND2x4_ASAP7_75t_L g457 ( .A(n_307), .B(n_352), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_307), .B(n_366), .Y(n_493) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g348 ( .A(n_308), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g495 ( .A(n_311), .Y(n_495) );
BUFx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g356 ( .A(n_312), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_312), .B(n_323), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_312), .B(n_331), .Y(n_415) );
BUFx2_ASAP7_75t_L g419 ( .A(n_313), .Y(n_419) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_317), .B(n_406), .Y(n_405) );
INVxp67_ASAP7_75t_L g422 ( .A(n_317), .Y(n_422) );
INVx1_ASAP7_75t_L g392 ( .A(n_318), .Y(n_392) );
AND2x2_ASAP7_75t_L g465 ( .A(n_318), .B(n_466), .Y(n_465) );
BUFx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_326), .B1(n_328), .B2(n_330), .Y(n_320) );
NOR2x1_ASAP7_75t_L g321 ( .A(n_322), .B(n_325), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g454 ( .A(n_323), .B(n_434), .Y(n_454) );
AND2x2_ASAP7_75t_L g331 ( .A(n_324), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g393 ( .A(n_325), .Y(n_393) );
AND2x2_ASAP7_75t_L g328 ( .A(n_327), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g376 ( .A(n_329), .Y(n_376) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
AND2x2_ASAP7_75t_L g418 ( .A(n_331), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_331), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g481 ( .A(n_331), .Y(n_481) );
INVx2_ASAP7_75t_L g344 ( .A(n_332), .Y(n_344) );
NAND2x1_ASAP7_75t_SL g334 ( .A(n_335), .B(n_355), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_343), .B1(n_345), .B2(n_353), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI32xp33_ASAP7_75t_L g410 ( .A1(n_342), .A2(n_411), .A3(n_412), .B1(n_413), .B2(n_415), .Y(n_410) );
NOR2x1_ASAP7_75t_L g347 ( .A(n_344), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g357 ( .A(n_344), .Y(n_357) );
AND2x2_ASAP7_75t_L g449 ( .A(n_344), .B(n_367), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_346), .B(n_350), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g378 ( .A(n_349), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g386 ( .A(n_349), .Y(n_386) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g360 ( .A(n_354), .Y(n_360) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_356), .A2(n_433), .B(n_435), .Y(n_432) );
AND2x2_ASAP7_75t_L g478 ( .A(n_357), .B(n_367), .Y(n_478) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI21xp33_ASAP7_75t_L g377 ( .A1(n_361), .A2(n_378), .B(n_380), .Y(n_377) );
A2O1A1Ixp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_368), .B(n_374), .C(n_377), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2x1_ASAP7_75t_L g368 ( .A(n_369), .B(n_372), .Y(n_368) );
INVx1_ASAP7_75t_L g471 ( .A(n_369), .Y(n_471) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_371), .Y(n_475) );
NAND2x1_ASAP7_75t_L g462 ( .A(n_372), .B(n_457), .Y(n_462) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g438 ( .A(n_378), .Y(n_438) );
NOR2x1_ASAP7_75t_L g381 ( .A(n_382), .B(n_445), .Y(n_381) );
NAND4xp25_ASAP7_75t_L g382 ( .A(n_383), .B(n_409), .C(n_425), .D(n_436), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_393), .B(n_394), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g441 ( .A(n_386), .B(n_434), .Y(n_441) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g452 ( .A(n_389), .Y(n_452) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
NAND2x1p5_ASAP7_75t_L g443 ( .A(n_392), .B(n_444), .Y(n_443) );
OAI21xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_398), .B(n_405), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_401), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_416), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_420), .B1(n_422), .B2(n_423), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g433 ( .A(n_430), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g487 ( .A(n_430), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_441), .B(n_442), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
AND2x4_ASAP7_75t_L g473 ( .A(n_440), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g488 ( .A1(n_444), .A2(n_489), .B1(n_491), .B2(n_493), .C(n_494), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_467), .C(n_488), .Y(n_445) );
NOR3xp33_ASAP7_75t_SL g446 ( .A(n_447), .B(n_455), .C(n_461), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_450), .B1(n_452), .B2(n_453), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_453), .A2(n_495), .B1(n_496), .B2(n_498), .Y(n_494) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B(n_464), .Y(n_461) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_470), .B1(n_472), .B2(n_473), .C(n_476), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVxp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OAI221xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_479), .B1(n_480), .B2(n_481), .C(n_482), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND3xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .C(n_486), .Y(n_482) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx2_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
CKINVDCx6p67_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_506), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVxp67_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AO21x2_ASAP7_75t_L g752 ( .A1(n_507), .A2(n_698), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OAI221xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_695), .B1(n_702), .B2(n_703), .C(n_744), .Y(n_511) );
INVx1_ASAP7_75t_L g702 ( .A(n_513), .Y(n_702) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_606), .Y(n_514) );
OAI31xp33_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_534), .A3(n_544), .B(n_601), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_518), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .Y(n_518) );
NAND2x1_ASAP7_75t_L g540 ( .A(n_519), .B(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OR2x6_ASAP7_75t_SL g530 ( .A(n_520), .B(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_L g535 ( .A(n_520), .B(n_536), .Y(n_535) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
INVx1_ASAP7_75t_L g553 ( .A(n_521), .Y(n_553) );
BUFx2_ASAP7_75t_L g585 ( .A(n_521), .Y(n_585) );
AND2x2_ASAP7_75t_L g552 ( .A(n_522), .B(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g568 ( .A(n_522), .B(n_553), .Y(n_568) );
AND2x4_ASAP7_75t_L g584 ( .A(n_522), .B(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx3_ASAP7_75t_L g562 ( .A(n_524), .Y(n_562) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_525), .Y(n_577) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_528), .Y(n_525) );
AND2x4_ASAP7_75t_L g532 ( .A(n_526), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g599 ( .A(n_526), .Y(n_599) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g550 ( .A(n_527), .B(n_528), .Y(n_550) );
INVx2_ASAP7_75t_L g533 ( .A(n_528), .Y(n_533) );
BUFx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_532), .Y(n_558) );
AND2x4_ASAP7_75t_L g543 ( .A(n_533), .B(n_538), .Y(n_543) );
INVx8_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g593 ( .A(n_539), .Y(n_593) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx3_ASAP7_75t_L g578 ( .A(n_542), .Y(n_578) );
INVx4_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_543), .Y(n_566) );
NAND5xp2_ASAP7_75t_L g544 ( .A(n_545), .B(n_554), .C(n_569), .D(n_586), .E(n_588), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
AND2x4_ASAP7_75t_L g547 ( .A(n_548), .B(n_551), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g560 ( .A(n_549), .Y(n_560) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g581 ( .A(n_550), .Y(n_581) );
INVx3_ASAP7_75t_L g587 ( .A(n_551), .Y(n_587) );
BUFx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g595 ( .A(n_552), .Y(n_595) );
OAI211xp5_ASAP7_75t_SL g554 ( .A1(n_555), .A2(n_556), .B(n_559), .C(n_563), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_555), .A2(n_627), .B1(n_628), .B2(n_632), .Y(n_626) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g572 ( .A(n_558), .Y(n_572) );
BUFx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
NAND3xp33_ASAP7_75t_L g729 ( .A(n_567), .B(n_593), .C(n_730), .Y(n_729) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OAI211xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_573), .B(n_574), .C(n_579), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
OR2x6_ASAP7_75t_L g586 ( .A(n_572), .B(n_587), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_573), .A2(n_609), .B1(n_610), .B2(n_620), .Y(n_608) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
INVx5_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
BUFx6f_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B1(n_596), .B2(n_597), .Y(n_588) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_SL g736 ( .A(n_592), .Y(n_736) );
AND2x4_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g600 ( .A(n_595), .Y(n_600) );
OAI221xp5_ASAP7_75t_SL g673 ( .A1(n_596), .A2(n_674), .B1(n_676), .B2(n_677), .C(n_679), .Y(n_673) );
AND2x4_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx3_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x4_ASAP7_75t_L g617 ( .A(n_605), .B(n_618), .Y(n_617) );
NAND2x1p5_ASAP7_75t_L g640 ( .A(n_605), .B(n_641), .Y(n_640) );
AND2x4_ASAP7_75t_SL g651 ( .A(n_605), .B(n_641), .Y(n_651) );
AND3x1_ASAP7_75t_L g656 ( .A(n_605), .B(n_657), .C(n_659), .Y(n_656) );
INVx2_ASAP7_75t_L g691 ( .A(n_605), .Y(n_691) );
NOR3xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_636), .C(n_652), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_626), .Y(n_607) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x4_ASAP7_75t_L g611 ( .A(n_612), .B(n_617), .Y(n_611) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g672 ( .A(n_613), .Y(n_672) );
INVx5_ASAP7_75t_L g685 ( .A(n_613), .Y(n_685) );
AND2x4_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g631 ( .A(n_614), .Y(n_631) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_614), .Y(n_644) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g624 ( .A(n_615), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_615), .B(n_616), .Y(n_639) );
INVx2_ASAP7_75t_L g625 ( .A(n_616), .Y(n_625) );
AND2x2_ASAP7_75t_L g622 ( .A(n_617), .B(n_623), .Y(n_622) );
AND2x6_ASAP7_75t_L g628 ( .A(n_617), .B(n_629), .Y(n_628) );
AND2x4_ASAP7_75t_L g633 ( .A(n_617), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g658 ( .A(n_619), .Y(n_658) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x4_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g666 ( .A(n_624), .B(n_625), .Y(n_666) );
AND2x4_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g650 ( .A(n_630), .Y(n_650) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_634), .Y(n_670) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
BUFx3_ASAP7_75t_L g682 ( .A(n_635), .Y(n_682) );
OR2x4_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx2_ASAP7_75t_SL g662 ( .A(n_638), .Y(n_662) );
INVx1_ASAP7_75t_L g675 ( .A(n_638), .Y(n_675) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OR2x6_ASAP7_75t_L g642 ( .A(n_640), .B(n_643), .Y(n_642) );
OR2x6_ASAP7_75t_L g694 ( .A(n_640), .B(n_678), .Y(n_694) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
BUFx4f_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x4_ASAP7_75t_L g647 ( .A(n_648), .B(n_651), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_660), .B1(n_673), .B2(n_686), .C(n_692), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OAI221xp5_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_663), .B1(n_664), .B2(n_667), .C(n_668), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
BUFx12f_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_666), .Y(n_678) );
BUFx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
BUFx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx3_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx3_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
BUFx6f_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
BUFx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OR2x6_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_700), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
BUFx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g727 ( .A(n_699), .Y(n_727) );
AND2x2_ASAP7_75t_L g753 ( .A(n_700), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_701), .B(n_727), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_702), .A2(n_745), .B1(n_748), .B2(n_750), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_723), .B1(n_737), .B2(n_738), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_704), .A2(n_737), .B1(n_746), .B2(n_747), .Y(n_745) );
XOR2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_712), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B1(n_708), .B2(n_709), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_710), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_716), .B1(n_721), .B2(n_722), .Y(n_712) );
INVx1_ASAP7_75t_L g721 ( .A(n_713), .Y(n_721) );
INVx1_ASAP7_75t_L g715 ( .A(n_714), .Y(n_715) );
INVx1_ASAP7_75t_L g722 ( .A(n_716), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_716) );
INVx1_ASAP7_75t_SL g719 ( .A(n_717), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_718), .Y(n_720) );
BUFx3_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx3_ASAP7_75t_L g746 ( .A(n_724), .Y(n_746) );
AND2x6_ASAP7_75t_L g724 ( .A(n_725), .B(n_732), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .Y(n_725) );
INVxp67_ASAP7_75t_L g742 ( .A(n_726), .Y(n_742) );
INVx1_ASAP7_75t_L g754 ( .A(n_727), .Y(n_754) );
INVxp67_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_729), .B(n_736), .Y(n_743) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
CKINVDCx11_ASAP7_75t_R g734 ( .A(n_731), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_735), .Y(n_732) );
CKINVDCx5p33_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx4_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
BUFx4f_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
BUFx3_ASAP7_75t_L g747 ( .A(n_740), .Y(n_747) );
INVx4_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
endmodule