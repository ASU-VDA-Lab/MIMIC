module real_jpeg_7941_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_23;
wire n_11;
wire n_14;
wire n_7;
wire n_22;
wire n_18;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

OR2x2_ASAP7_75t_SL g16 ( 
.A(n_1),
.B(n_17),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_2),
.B(n_10),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_10),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_SL g8 ( 
.A1(n_5),
.A2(n_9),
.B(n_11),
.Y(n_8)
);

AOI22xp33_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_15),
.B1(n_22),
.B2(n_23),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_12),
.B(n_14),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_8),
.B(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_13),
.A2(n_16),
.B(n_18),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_19),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);


endmodule