module fake_jpeg_26299_n_141 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_26),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_27),
.A2(n_16),
.B1(n_18),
.B2(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_26),
.A2(n_16),
.B1(n_12),
.B2(n_18),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_11),
.B1(n_26),
.B2(n_25),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_20),
.C(n_17),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_34),
.B1(n_31),
.B2(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_46),
.Y(n_51)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_44),
.B1(n_10),
.B2(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_11),
.B1(n_19),
.B2(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_10),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_24),
.Y(n_46)
);

AO22x1_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_24),
.B1(n_21),
.B2(n_22),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_33),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_31),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_57),
.B(n_37),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_29),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_6),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_47),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_33),
.B(n_30),
.C(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_48),
.B1(n_39),
.B2(n_37),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_22),
.Y(n_62)
);

A2O1A1O1Ixp25_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_56),
.B(n_49),
.C(n_51),
.D(n_47),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_63),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_57),
.C(n_27),
.Y(n_86)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_72),
.B(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_73),
.B(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_43),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_79),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_84),
.B1(n_32),
.B2(n_71),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_50),
.B(n_57),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_78),
.B(n_86),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_6),
.C(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_74),
.B(n_62),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_SL g90 ( 
.A(n_81),
.B(n_20),
.C(n_22),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_57),
.B(n_68),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_32),
.B1(n_21),
.B2(n_28),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_28),
.B1(n_21),
.B2(n_27),
.Y(n_100)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_90),
.B(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_22),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_95),
.C(n_97),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_67),
.C(n_24),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_76),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_100),
.B1(n_76),
.B2(n_78),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_67),
.C(n_27),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_107),
.Y(n_113)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_83),
.A3(n_95),
.B1(n_94),
.B2(n_90),
.C1(n_89),
.C2(n_100),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_106),
.B(n_111),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_99),
.A2(n_83),
.B1(n_87),
.B2(n_2),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

AOI321xp33_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_27),
.A3(n_28),
.B1(n_20),
.B2(n_4),
.C(n_7),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_114),
.B(n_116),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_1),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_108),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_1),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_118),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_2),
.C(n_4),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_124),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_117),
.B(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_125),
.B(n_107),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_122),
.A2(n_112),
.B1(n_109),
.B2(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_128),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_110),
.B1(n_123),
.B2(n_119),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_127),
.B(n_130),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_115),
.C(n_7),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_130),
.B(n_8),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_126),
.B(n_7),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_132),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_135),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_8),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_137),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_140),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_9),
.B(n_0),
.Y(n_140)
);


endmodule