module fake_jpeg_2671_n_88 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_88);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_19),
.B(n_7),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_24),
.B(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_7),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_30),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_18),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_47)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_21),
.B(n_5),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

OR2x2_ASAP7_75t_SL g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_23),
.B(n_22),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_32),
.C(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_35),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_33),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_39),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_56),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_46),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_33),
.C(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_58),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_59),
.B(n_37),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_63),
.B(n_65),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_48),
.B1(n_42),
.B2(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_48),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_56),
.C(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_72),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_70),
.B(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_53),
.B1(n_48),
.B2(n_1),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_64),
.C(n_1),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_74),
.A2(n_78),
.B(n_73),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_79),
.A2(n_76),
.B(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_80),
.A2(n_81),
.B(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_10),
.C(n_11),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_4),
.B(n_8),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_85),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_12),
.Y(n_88)
);


endmodule