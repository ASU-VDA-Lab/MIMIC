module real_jpeg_3751_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_1),
.B(n_42),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_1),
.B(n_54),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_1),
.A2(n_25),
.B(n_26),
.C(n_228),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_1),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_1),
.B(n_31),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_229),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_1),
.B(n_61),
.C(n_64),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_229),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_1),
.B(n_115),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_1),
.B(n_59),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_45),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_45),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_2),
.A2(n_45),
.B1(n_61),
.B2(n_65),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_3),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_4),
.A2(n_38),
.B1(n_61),
.B2(n_65),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_5),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_147),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_147),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_5),
.A2(n_61),
.B1(n_65),
.B2(n_147),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_53),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_53),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_8),
.A2(n_53),
.B1(n_61),
.B2(n_65),
.Y(n_138)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_11),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_179),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_179),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_11),
.A2(n_61),
.B1(n_65),
.B2(n_179),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_13),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_85),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_85),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_13),
.A2(n_61),
.B1(n_65),
.B2(n_85),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_14),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_77),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_77),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_14),
.A2(n_61),
.B1(n_65),
.B2(n_77),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_15),
.A2(n_42),
.B1(n_43),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_15),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_125),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_125),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_15),
.A2(n_61),
.B1(n_65),
.B2(n_125),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_91),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_90),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_21),
.B(n_78),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_57),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_39),
.B1(n_55),
.B2(n_56),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_23),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_31),
.B(n_36),
.Y(n_23)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_24),
.B(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_24),
.A2(n_31),
.B1(n_196),
.B2(n_213),
.Y(n_241)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_30),
.C(n_31),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_26),
.Y(n_30)
);

AO22x2_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_26),
.A2(n_27),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

AOI32xp33_ASAP7_75t_L g199 ( 
.A1(n_26),
.A2(n_43),
.A3(n_48),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp33_ASAP7_75t_SL g201 ( 
.A(n_27),
.B(n_50),
.Y(n_201)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_31),
.B(n_176),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_32),
.A2(n_33),
.B1(n_63),
.B2(n_64),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g228 ( 
.A1(n_32),
.A2(n_35),
.B(n_229),
.Y(n_228)
);

INVx5_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_33),
.B(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_37),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_52),
.B2(n_54),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_47),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_51)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_43),
.A2(n_75),
.B(n_229),
.C(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_46),
.B(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_46),
.A2(n_54),
.B1(n_146),
.B2(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_51),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_75),
.B1(n_76),
.B2(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_47),
.A2(n_84),
.B(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_47),
.B(n_124),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_47),
.A2(n_122),
.B(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_48),
.Y(n_50)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_70),
.C(n_74),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_70),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_SL g86 ( 
.A(n_58),
.B(n_83),
.C(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_58),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_66),
.B(n_68),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_59),
.A2(n_66),
.B1(n_120),
.B2(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_59),
.A2(n_66),
.B1(n_141),
.B2(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_59),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_60),
.A2(n_69),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_60),
.A2(n_101),
.B1(n_102),
.B2(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_60),
.A2(n_244),
.B(n_245),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_60),
.A2(n_245),
.B(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_60),
.A2(n_101),
.B1(n_222),
.B2(n_256),
.Y(n_267)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_61),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_61),
.B(n_285),
.Y(n_284)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_66),
.A2(n_221),
.B(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_66),
.B(n_225),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_71),
.A2(n_73),
.B1(n_89),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_71),
.A2(n_73),
.B1(n_99),
.B2(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_71),
.A2(n_195),
.B(n_197),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_71),
.A2(n_197),
.B(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_73),
.A2(n_143),
.B(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_73),
.A2(n_175),
.B(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_75),
.A2(n_145),
.B(n_148),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.C(n_86),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_79),
.A2(n_83),
.B1(n_104),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_86),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AO21x1_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_155),
.B(n_326),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_150),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_126),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_95),
.B(n_126),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_107),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_103),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_98),
.B(n_100),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_97),
.B(n_103),
.C(n_107),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_101),
.A2(n_224),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B(n_121),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_109),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_118),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_111),
.B1(n_121),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_110),
.A2(n_111),
.B1(n_118),
.B2(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_115),
.B(n_116),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_112),
.A2(n_115),
.B1(n_138),
.B2(n_172),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_112),
.A2(n_229),
.B(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_113),
.A2(n_114),
.B1(n_117),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_113),
.A2(n_114),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_113),
.A2(n_114),
.B1(n_204),
.B2(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_113),
.B(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_113),
.A2(n_260),
.B(n_261),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_113),
.A2(n_114),
.B1(n_260),
.B2(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_114),
.A2(n_219),
.B(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_114),
.B(n_233),
.Y(n_262)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_115),
.A2(n_232),
.B(n_289),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_118),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_132),
.C(n_133),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_128),
.B1(n_132),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_142),
.C(n_144),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_135),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_136),
.A2(n_139),
.B1(n_140),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_142),
.B(n_144),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_149),
.B(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_150),
.A2(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_151),
.B(n_154),
.Y(n_328)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_180),
.B(n_325),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_157),
.B(n_160),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_166),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_173),
.C(n_177),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_168),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_169),
.B(n_171),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_170),
.Y(n_244)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_174),
.B1(n_177),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

OAI21x1_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_206),
.B(n_324),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_182),
.B(n_184),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.C(n_191),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_185),
.B(n_189),
.Y(n_309)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_186),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_191),
.B(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.C(n_198),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_192),
.B(n_194),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_198),
.B(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_199),
.A2(n_202),
.B1(n_203),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_199),
.Y(n_248)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI31xp33_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_306),
.A3(n_316),
.B(n_321),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_250),
.B(n_305),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_234),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_209),
.B(n_234),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_220),
.C(n_226),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_210),
.B(n_302),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_211),
.B(n_215),
.C(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_220),
.B(n_226),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_230),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_246),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_235),
.B(n_247),
.C(n_249),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_236),
.B(n_241),
.C(n_242),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_300),
.B(n_304),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_269),
.B(n_299),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_263),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_253),
.B(n_263),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.C(n_258),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_259),
.B1(n_278),
.B2(n_280),
.Y(n_277)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_267),
.C(n_268),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_281),
.B(n_298),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_277),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_277),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_272),
.A2(n_273),
.B1(n_275),
.B2(n_296),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_292),
.B(n_297),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_287),
.B(n_291),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_290),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_289),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_295),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_303),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI21xp33_ASAP7_75t_L g321 ( 
.A1(n_307),
.A2(n_322),
.B(n_323),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_310),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.C(n_314),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_318),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_313),
.A2(n_314),
.B1(n_315),
.B2(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_320),
.Y(n_322)
);


endmodule