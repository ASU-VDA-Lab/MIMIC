module fake_jpeg_24967_n_75 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_75);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_75;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_67;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_0),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_19),
.A2(n_23),
.B1(n_11),
.B2(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_10),
.B1(n_14),
.B2(n_16),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_11),
.C(n_16),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_12),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_17),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_35),
.B(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_20),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_26),
.C(n_21),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_27),
.B(n_26),
.Y(n_39)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_21),
.Y(n_49)
);

AND2x6_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_45),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_26),
.B1(n_23),
.B2(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_26),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_38),
.C(n_21),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_23),
.B(n_22),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_31),
.A2(n_22),
.B1(n_18),
.B2(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_18),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_46),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_50),
.B(n_53),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_54),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_60),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_48),
.C(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_44),
.B1(n_41),
.B2(n_50),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_61),
.A2(n_64),
.B1(n_4),
.B2(n_7),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_0),
.C(n_1),
.Y(n_67)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_66),
.B(n_67),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_59),
.B(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_68),
.B(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_70),
.B(n_4),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_5),
.C(n_2),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_71),
.C(n_5),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_1),
.Y(n_75)
);


endmodule