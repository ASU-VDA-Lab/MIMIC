module fake_jpeg_13990_n_483 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_483);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_483;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_56),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_22),
.B(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_57),
.B(n_58),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_59),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_60),
.Y(n_164)
);

CKINVDCx9p33_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_22),
.B(n_14),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_63),
.B(n_64),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_13),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_65),
.B(n_67),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_45),
.B(n_0),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_23),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_69),
.B(n_84),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_70),
.Y(n_161)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_72),
.B(n_78),
.Y(n_132)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_74),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_75),
.Y(n_173)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_37),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_80),
.B(n_82),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_83),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_23),
.B(n_0),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_32),
.B(n_12),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_101),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

CKINVDCx6p67_ASAP7_75t_R g196 ( 
.A(n_87),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_88),
.Y(n_193)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_89),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_25),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_90),
.B(n_99),
.Y(n_172)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_91),
.Y(n_174)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_96),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

BUFx2_ASAP7_75t_SL g183 ( 
.A(n_97),
.Y(n_183)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_25),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_100),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_50),
.B(n_1),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_50),
.B(n_1),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_107),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_21),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_104),
.B(n_106),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_32),
.B(n_2),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_105),
.B(n_111),
.Y(n_177)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_47),
.B(n_2),
.Y(n_107)
);

INVxp67_ASAP7_75t_SL g108 ( 
.A(n_19),
.Y(n_108)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_34),
.B(n_2),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_21),
.Y(n_113)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_20),
.Y(n_114)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_30),
.Y(n_115)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_18),
.Y(n_116)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_20),
.Y(n_117)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_117),
.Y(n_202)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_18),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_119),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_20),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_120),
.B(n_3),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_68),
.B(n_53),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_123),
.B(n_132),
.Y(n_214)
);

NAND2x1_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_31),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_125),
.A2(n_179),
.B(n_197),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_31),
.C(n_28),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_127),
.B(n_170),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_114),
.A2(n_31),
.B1(n_28),
.B2(n_27),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_131),
.A2(n_144),
.B1(n_147),
.B2(n_149),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_61),
.A2(n_19),
.B1(n_28),
.B2(n_27),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_108),
.A2(n_27),
.B1(n_26),
.B2(n_52),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_74),
.A2(n_54),
.B1(n_52),
.B2(n_44),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_55),
.A2(n_53),
.B1(n_39),
.B2(n_34),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_151),
.A2(n_155),
.B1(n_157),
.B2(n_160),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_59),
.A2(n_44),
.B1(n_26),
.B2(n_54),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_59),
.A2(n_39),
.B1(n_4),
.B2(n_5),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_60),
.A2(n_97),
.B1(n_102),
.B2(n_94),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_117),
.A2(n_12),
.B1(n_6),
.B2(n_7),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_163),
.A2(n_165),
.B1(n_175),
.B2(n_178),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_66),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_109),
.A2(n_3),
.B1(n_8),
.B2(n_9),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_185),
.B1(n_191),
.B2(n_195),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_56),
.B(n_8),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g227 ( 
.A(n_171),
.B(n_167),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_60),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_97),
.A2(n_11),
.B1(n_12),
.B2(n_91),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_98),
.A2(n_120),
.B(n_87),
.C(n_106),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_179),
.B(n_125),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_85),
.A2(n_88),
.B1(n_83),
.B2(n_81),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_184),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_70),
.A2(n_75),
.B1(n_77),
.B2(n_79),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_113),
.A2(n_100),
.B1(n_96),
.B2(n_71),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_110),
.A2(n_115),
.B1(n_119),
.B2(n_87),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_119),
.A2(n_71),
.B1(n_110),
.B2(n_115),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_106),
.A2(n_107),
.B1(n_103),
.B2(n_101),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_190),
.B(n_199),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_107),
.A2(n_101),
.B1(n_103),
.B2(n_90),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_L g195 ( 
.A1(n_55),
.A2(n_79),
.B1(n_77),
.B2(n_66),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_61),
.A2(n_51),
.B1(n_46),
.B2(n_108),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_69),
.B(n_84),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_90),
.A2(n_99),
.B1(n_107),
.B2(n_33),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_201),
.A2(n_195),
.B1(n_133),
.B2(n_139),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_204),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_205),
.A2(n_243),
.B(n_270),
.Y(n_293)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_206),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_128),
.B(n_122),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_207),
.B(n_211),
.Y(n_289)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_124),
.Y(n_208)
);

INVx6_ASAP7_75t_SL g287 ( 
.A(n_208),
.Y(n_287)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_209),
.Y(n_276)
);

BUFx16f_ASAP7_75t_L g210 ( 
.A(n_124),
.Y(n_210)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_210),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_134),
.B(n_153),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_141),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_212),
.B(n_257),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_214),
.B(n_219),
.Y(n_305)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_146),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_215),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_172),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_216),
.B(n_218),
.Y(n_278)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_140),
.Y(n_217)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_217),
.Y(n_285)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_138),
.C(n_129),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_152),
.B(n_194),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_140),
.Y(n_220)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_220),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_121),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_221),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_168),
.B(n_182),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_222),
.B(n_225),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_121),
.Y(n_223)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_223),
.Y(n_315)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_130),
.Y(n_224)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_224),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_196),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_130),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_226),
.Y(n_281)
);

XOR2x2_ASAP7_75t_SL g301 ( 
.A(n_227),
.B(n_264),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_142),
.Y(n_228)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_228),
.Y(n_302)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_180),
.Y(n_229)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_229),
.Y(n_312)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_158),
.Y(n_230)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_230),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_142),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_233),
.A2(n_238),
.B1(n_240),
.B2(n_254),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_235),
.B(n_242),
.Y(n_282)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_180),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_237),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_161),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_171),
.B(n_164),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_239),
.B(n_244),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_161),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_166),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_241),
.Y(n_272)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_166),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_171),
.B(n_143),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_145),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_245),
.B(n_246),
.Y(n_288)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_196),
.B(n_135),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_247),
.B(n_248),
.Y(n_292)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_126),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g249 ( 
.A(n_192),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_249),
.B(n_250),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_187),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_164),
.B(n_186),
.Y(n_251)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_251),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_136),
.B(n_154),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_252),
.Y(n_295)
);

OA21x2_ASAP7_75t_L g294 ( 
.A1(n_253),
.A2(n_227),
.B(n_270),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_173),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_137),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_255),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_156),
.B(n_155),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_256),
.Y(n_318)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_150),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_203),
.B(n_174),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_260),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_188),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_259),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_192),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_176),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_261),
.B(n_262),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_127),
.B(n_145),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_173),
.Y(n_263)
);

OA22x2_ASAP7_75t_L g310 ( 
.A1(n_263),
.A2(n_238),
.B1(n_254),
.B2(n_240),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_174),
.B(n_162),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_192),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_SL g314 ( 
.A1(n_265),
.A2(n_208),
.B(n_210),
.C(n_261),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_149),
.B(n_160),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_266),
.A2(n_267),
.B1(n_271),
.B2(n_234),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_148),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_176),
.B(n_147),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_198),
.Y(n_286)
);

AND2x6_ASAP7_75t_L g275 ( 
.A(n_212),
.B(n_184),
.Y(n_275)
);

A2O1A1O1Ixp25_ASAP7_75t_L g325 ( 
.A1(n_275),
.A2(n_296),
.B(n_210),
.C(n_265),
.D(n_249),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_253),
.A2(n_193),
.B1(n_159),
.B2(n_144),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_279),
.A2(n_283),
.B1(n_318),
.B2(n_308),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_178),
.C(n_175),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_283),
.B(n_286),
.C(n_321),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_286),
.B(n_293),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_213),
.A2(n_157),
.B1(n_159),
.B2(n_183),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_291),
.A2(n_297),
.B1(n_313),
.B2(n_321),
.Y(n_342)
);

NOR2x1_ASAP7_75t_L g333 ( 
.A(n_294),
.B(n_204),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_L g296 ( 
.A1(n_227),
.A2(n_259),
.B(n_234),
.C(n_232),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_231),
.A2(n_268),
.B(n_236),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_303),
.A2(n_309),
.B(n_220),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_229),
.A2(n_237),
.B(n_224),
.Y(n_309)
);

AO21x2_ASAP7_75t_L g339 ( 
.A1(n_310),
.A2(n_314),
.B(n_287),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_241),
.A2(n_242),
.B1(n_255),
.B2(n_257),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_235),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_322),
.B(n_323),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_305),
.B(n_248),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_324),
.B(n_325),
.Y(n_365)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_290),
.Y(n_326)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_326),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_350),
.C(n_314),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_303),
.A2(n_246),
.B1(n_209),
.B2(n_263),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_328),
.A2(n_329),
.B1(n_331),
.B2(n_346),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_319),
.A2(n_223),
.B1(n_233),
.B2(n_221),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_319),
.A2(n_228),
.B1(n_217),
.B2(n_249),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_290),
.Y(n_332)
);

NOR2x1_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_284),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_280),
.B(n_204),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_334),
.B(n_336),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_318),
.A2(n_206),
.B1(n_291),
.B2(n_281),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_335),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_280),
.B(n_206),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_293),
.B(n_301),
.C(n_294),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_337),
.B(n_344),
.C(n_349),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_295),
.B(n_278),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_338),
.B(n_341),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_339),
.Y(n_376)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_290),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_343),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_295),
.B(n_320),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_342),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_287),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_301),
.B(n_294),
.C(n_300),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_274),
.B(n_300),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_345),
.B(n_348),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_281),
.A2(n_274),
.B(n_298),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_347),
.A2(n_314),
.B(n_299),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_292),
.B(n_298),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_296),
.C(n_279),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_317),
.B(n_288),
.C(n_275),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_304),
.B(n_306),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_351),
.B(n_357),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_277),
.A2(n_309),
.B1(n_310),
.B2(n_272),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_352),
.A2(n_284),
.B1(n_273),
.B2(n_311),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_306),
.A2(n_312),
.B1(n_272),
.B2(n_285),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_353),
.A2(n_273),
.B1(n_311),
.B2(n_352),
.Y(n_378)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_276),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_354),
.B(n_355),
.Y(n_362)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_276),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_282),
.B(n_316),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_356),
.B(n_347),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_304),
.B(n_312),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_314),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_360),
.Y(n_388)
);

OAI32xp33_ASAP7_75t_L g360 ( 
.A1(n_345),
.A2(n_307),
.A3(n_302),
.B1(n_310),
.B2(n_314),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_307),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_364),
.B(n_370),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_367),
.B(n_371),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_330),
.B(n_299),
.C(n_285),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_368),
.B(n_330),
.C(n_343),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_350),
.A2(n_310),
.B1(n_315),
.B2(n_302),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_369),
.A2(n_384),
.B1(n_328),
.B2(n_325),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_357),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_373),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_331),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_378),
.Y(n_403)
);

OAI21xp33_ASAP7_75t_L g399 ( 
.A1(n_380),
.A2(n_356),
.B(n_326),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_330),
.B(n_346),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_333),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_342),
.A2(n_324),
.B1(n_327),
.B2(n_344),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_386),
.B(n_389),
.C(n_405),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_385),
.B(n_337),
.C(n_351),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_372),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_391),
.B(n_394),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_372),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_392),
.B(n_393),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_362),
.Y(n_394)
);

NOR2xp67_ASAP7_75t_SL g395 ( 
.A(n_367),
.B(n_333),
.Y(n_395)
);

AOI21x1_ASAP7_75t_L g421 ( 
.A1(n_395),
.A2(n_359),
.B(n_371),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_366),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_397),
.B(n_379),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_380),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_400),
.Y(n_419)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_382),
.Y(n_401)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_401),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_358),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_402),
.B(n_404),
.Y(n_427)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_382),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_329),
.C(n_355),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_332),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_406),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_381),
.B(n_340),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_407),
.B(n_362),
.C(n_358),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_377),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_408),
.B(n_377),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_354),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_409),
.B(n_374),
.Y(n_422)
);

MAJx2_ASAP7_75t_L g435 ( 
.A(n_410),
.B(n_423),
.C(n_424),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_384),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_411),
.B(n_421),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_403),
.A2(n_361),
.B1(n_369),
.B2(n_365),
.Y(n_414)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_414),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_415),
.B(n_425),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_403),
.A2(n_383),
.B1(n_365),
.B2(n_361),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_416),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_387),
.A2(n_359),
.B(n_365),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_417),
.A2(n_398),
.B(n_373),
.Y(n_445)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_422),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_389),
.B(n_368),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_396),
.B(n_363),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_388),
.A2(n_376),
.B1(n_363),
.B2(n_373),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_387),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_429),
.B(n_405),
.C(n_386),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_L g431 ( 
.A1(n_412),
.A2(n_400),
.B1(n_392),
.B2(n_390),
.Y(n_431)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_431),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_413),
.B(n_401),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_432),
.B(n_443),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_433),
.A2(n_441),
.B1(n_442),
.B2(n_426),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_411),
.C(n_418),
.Y(n_450)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_419),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_439),
.B(n_444),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_420),
.A2(n_388),
.B1(n_404),
.B2(n_400),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_420),
.A2(n_406),
.B1(n_409),
.B2(n_393),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_428),
.B(n_366),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_429),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_445),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_433),
.Y(n_460)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_432),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_SL g463 ( 
.A1(n_449),
.A2(n_451),
.B1(n_453),
.B2(n_455),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_450),
.B(n_452),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_442),
.A2(n_414),
.B1(n_416),
.B2(n_417),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_438),
.B(n_418),
.C(n_423),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_443),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_441),
.A2(n_378),
.B1(n_427),
.B2(n_375),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_435),
.B(n_424),
.C(n_421),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_456),
.B(n_434),
.C(n_435),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_458),
.B(n_465),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_453),
.B(n_430),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_459),
.B(n_462),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_448),
.B(n_430),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_446),
.A2(n_436),
.B1(n_437),
.B2(n_445),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_440),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_450),
.C(n_435),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_466),
.B(n_456),
.Y(n_472)
);

AOI21xp33_ASAP7_75t_L g467 ( 
.A1(n_459),
.A2(n_454),
.B(n_457),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_467),
.B(n_471),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_464),
.A2(n_451),
.B1(n_446),
.B2(n_447),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_463),
.A2(n_440),
.B1(n_449),
.B2(n_436),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_472),
.B(n_466),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_474),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_468),
.B(n_461),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_475),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_473),
.A2(n_472),
.B(n_470),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_478),
.A2(n_470),
.B(n_469),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_477),
.A2(n_476),
.B1(n_460),
.B2(n_454),
.Y(n_479)
);

NOR3xp33_ASAP7_75t_L g481 ( 
.A(n_479),
.B(n_480),
.C(n_419),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_481),
.A2(n_419),
.B(n_395),
.Y(n_482)
);

BUFx24_ASAP7_75t_SL g483 ( 
.A(n_482),
.Y(n_483)
);


endmodule