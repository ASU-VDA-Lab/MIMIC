module fake_jpeg_15760_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_4),
.B(n_3),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_14),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_14),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_17),
.B(n_20),
.Y(n_23)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_18),
.Y(n_30)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_12),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_0),
.C(n_1),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_13),
.A2(n_10),
.B1(n_9),
.B2(n_11),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_22),
.B1(n_6),
.B2(n_12),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_11),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_26),
.B(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_21),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_34),
.B(n_23),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_26),
.A2(n_15),
.B(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

OAI322xp33_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_27),
.A3(n_23),
.B1(n_28),
.B2(n_19),
.C1(n_18),
.C2(n_30),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_34),
.C(n_32),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_35),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_42),
.B1(n_40),
.B2(n_33),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_37),
.B(n_43),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_30),
.C(n_40),
.Y(n_46)
);


endmodule