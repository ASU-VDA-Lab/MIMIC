module fake_jpeg_12920_n_636 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_636);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_636;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_59),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_61),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_25),
.B(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_62),
.B(n_64),
.Y(n_170)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_63),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_8),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_66),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_67),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_69),
.Y(n_190)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

HAxp5_ASAP7_75t_SL g71 ( 
.A(n_45),
.B(n_26),
.CON(n_71),
.SN(n_71)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_71),
.B(n_76),
.Y(n_186)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_73),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_74),
.Y(n_212)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_31),
.Y(n_75)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_75),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_7),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_78),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_79),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_80),
.Y(n_202)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_82),
.Y(n_210)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_21),
.B(n_7),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_84),
.B(n_85),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_21),
.B(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_30),
.B(n_18),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_86),
.B(n_89),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_87),
.Y(n_213)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_88),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_30),
.B(n_7),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_91),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_58),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_92),
.B(n_97),
.Y(n_215)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g162 ( 
.A(n_96),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_32),
.B(n_7),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_99),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_104),
.Y(n_220)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_32),
.B(n_9),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_107),
.B(n_108),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_37),
.B(n_9),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_24),
.Y(n_110)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_37),
.B(n_6),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_119),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_25),
.Y(n_113)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_115),
.Y(n_192)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_36),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_116),
.Y(n_166)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_25),
.Y(n_117)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_40),
.B(n_6),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_25),
.Y(n_121)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_121),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_46),
.Y(n_122)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_122),
.Y(n_211)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_123),
.Y(n_218)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_44),
.Y(n_124)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_38),
.Y(n_126)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_48),
.Y(n_127)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_38),
.Y(n_128)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

BUFx12f_ASAP7_75t_SL g129 ( 
.A(n_48),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_129),
.B(n_54),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_71),
.A2(n_26),
.B1(n_48),
.B2(n_53),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_132),
.A2(n_154),
.B1(n_167),
.B2(n_168),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_62),
.B(n_44),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_134),
.B(n_57),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_26),
.B1(n_48),
.B2(n_113),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_50),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_157),
.B(n_196),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_70),
.B(n_49),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_160),
.B(n_197),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_113),
.A2(n_121),
.B1(n_115),
.B2(n_93),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_63),
.A2(n_34),
.B1(n_22),
.B2(n_19),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_81),
.Y(n_169)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_169),
.Y(n_232)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_73),
.Y(n_172)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_172),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_96),
.A2(n_47),
.B1(n_40),
.B2(n_42),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_174),
.A2(n_185),
.B1(n_58),
.B2(n_1),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_121),
.A2(n_101),
.B1(n_65),
.B2(n_59),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_176),
.A2(n_214),
.B1(n_106),
.B2(n_79),
.Y(n_244)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_60),
.Y(n_177)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_177),
.Y(n_246)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_61),
.Y(n_183)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_183),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_66),
.A2(n_22),
.B1(n_19),
.B2(n_56),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_67),
.Y(n_187)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_187),
.Y(n_265)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_188),
.Y(n_287)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_189),
.Y(n_293)
);

OA22x2_ASAP7_75t_SL g191 ( 
.A1(n_123),
.A2(n_45),
.B1(n_57),
.B2(n_47),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_191),
.A2(n_151),
.B(n_185),
.C(n_192),
.Y(n_270)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_69),
.Y(n_193)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_193),
.Y(n_294)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_74),
.Y(n_195)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_77),
.B(n_49),
.Y(n_197)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_82),
.Y(n_200)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_87),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_90),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_204),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_91),
.B(n_42),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_205),
.B(n_43),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_68),
.B(n_54),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_207),
.B(n_0),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_99),
.A2(n_34),
.B1(n_19),
.B2(n_22),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_104),
.Y(n_216)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_118),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_134),
.B(n_170),
.C(n_159),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_222),
.B(n_227),
.Y(n_321)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_155),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_223),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_224),
.B(n_259),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_154),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_228),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_143),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_230),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_170),
.B(n_198),
.C(n_150),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_231),
.B(n_236),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_139),
.B(n_215),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_233),
.B(n_245),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_186),
.B(n_122),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_235),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_144),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_238),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_131),
.B(n_43),
.C(n_50),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_239),
.B(n_242),
.Y(n_339)
);

OR2x2_ASAP7_75t_SL g338 ( 
.A(n_241),
.B(n_288),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_194),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_244),
.A2(n_247),
.B1(n_252),
.B2(n_261),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_217),
.B(n_55),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_56),
.B1(n_55),
.B2(n_109),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_250),
.Y(n_308)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_130),
.Y(n_251)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_251),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_L g252 ( 
.A1(n_214),
.A2(n_57),
.B1(n_58),
.B2(n_12),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_253),
.B(n_258),
.Y(n_347)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_206),
.Y(n_254)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_142),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_255),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_168),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_256),
.B(n_267),
.Y(n_356)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_137),
.Y(n_257)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_257),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_201),
.B(n_12),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_10),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_143),
.Y(n_260)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_260),
.Y(n_320)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_132),
.A2(n_57),
.B1(n_58),
.B2(n_10),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_186),
.A2(n_58),
.B1(n_1),
.B2(n_2),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_262),
.A2(n_295),
.B1(n_299),
.B2(n_252),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_201),
.B(n_196),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_263),
.B(n_264),
.Y(n_333)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_140),
.Y(n_266)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_266),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_166),
.B(n_10),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_141),
.Y(n_268)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_268),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_171),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_269),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_SL g332 ( 
.A1(n_270),
.A2(n_199),
.B(n_149),
.Y(n_332)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_209),
.Y(n_271)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_271),
.Y(n_331)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_173),
.Y(n_272)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_272),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_166),
.B(n_5),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_273),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_151),
.Y(n_274)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_274),
.Y(n_307)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_161),
.Y(n_275)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_275),
.Y(n_355)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_162),
.Y(n_276)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_276),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_277),
.A2(n_298),
.B1(n_220),
.B2(n_219),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_158),
.B(n_4),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_278),
.Y(n_326)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_178),
.Y(n_279)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_279),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_163),
.B(n_0),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_283),
.Y(n_300)
);

INVx4_ASAP7_75t_SL g281 ( 
.A(n_151),
.Y(n_281)
);

BUFx8_ASAP7_75t_L g353 ( 
.A(n_281),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_218),
.B(n_13),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_282),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_211),
.B(n_0),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_136),
.B(n_13),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_286),
.Y(n_314)
);

BUFx12f_ASAP7_75t_L g285 ( 
.A(n_146),
.Y(n_285)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_285),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_133),
.B(n_14),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_191),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_162),
.A2(n_16),
.B1(n_18),
.B2(n_3),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_289),
.A2(n_277),
.B1(n_292),
.B2(n_249),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_184),
.A2(n_145),
.B1(n_156),
.B2(n_182),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_290),
.A2(n_292),
.B(n_299),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_190),
.Y(n_291)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_291),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_180),
.A2(n_16),
.B1(n_18),
.B2(n_3),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_176),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_153),
.Y(n_296)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_296),
.Y(n_327)
);

BUFx12_ASAP7_75t_L g297 ( 
.A(n_147),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_297),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_180),
.A2(n_1),
.B1(n_2),
.B2(n_179),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_135),
.B(n_148),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_303),
.A2(n_313),
.B1(n_329),
.B2(n_351),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_L g313 ( 
.A1(n_228),
.A2(n_236),
.B1(n_270),
.B2(n_240),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_297),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_324),
.B(n_260),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_332),
.A2(n_287),
.B(n_239),
.Y(n_382)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_251),
.Y(n_334)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_334),
.Y(n_375)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_257),
.Y(n_335)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_335),
.Y(n_376)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_266),
.Y(n_336)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_336),
.Y(n_380)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_268),
.Y(n_337)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_337),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_237),
.B(n_208),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_340),
.B(n_357),
.Y(n_369)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_225),
.Y(n_342)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_342),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_345),
.B(n_281),
.Y(n_388)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_225),
.Y(n_346)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_346),
.Y(n_368)
);

O2A1O1Ixp33_ASAP7_75t_SL g349 ( 
.A1(n_262),
.A2(n_202),
.B(n_2),
.C(n_1),
.Y(n_349)
);

OA22x2_ASAP7_75t_L g365 ( 
.A1(n_349),
.A2(n_289),
.B1(n_274),
.B2(n_254),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_222),
.A2(n_208),
.B1(n_153),
.B2(n_181),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_235),
.A2(n_138),
.B1(n_144),
.B2(n_152),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_352),
.A2(n_238),
.B1(n_229),
.B2(n_250),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_241),
.B(n_152),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_235),
.A2(n_164),
.B1(n_175),
.B2(n_212),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_L g370 ( 
.A1(n_358),
.A2(n_276),
.B1(n_212),
.B2(n_175),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_359),
.Y(n_438)
);

A2O1A1O1Ixp25_ASAP7_75t_L g360 ( 
.A1(n_333),
.A2(n_231),
.B(n_264),
.C(n_283),
.D(n_280),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_360),
.A2(n_362),
.B(n_307),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_313),
.A2(n_290),
.B(n_227),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_303),
.A2(n_299),
.B1(n_223),
.B2(n_296),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_363),
.A2(n_364),
.B1(n_385),
.B2(n_398),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_317),
.A2(n_299),
.B1(n_249),
.B2(n_243),
.Y(n_364)
);

AND2x2_ASAP7_75t_SL g415 ( 
.A(n_365),
.B(n_353),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_356),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_366),
.B(n_367),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_340),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_370),
.A2(n_371),
.B1(n_372),
.B2(n_374),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_312),
.A2(n_345),
.B1(n_357),
.B2(n_338),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_305),
.Y(n_373)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_373),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_312),
.A2(n_164),
.B1(n_165),
.B2(n_210),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_341),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_377),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_304),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_378),
.B(n_381),
.Y(n_412)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_302),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_379),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_319),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_382),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_328),
.A2(n_338),
.B1(n_300),
.B2(n_321),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_383),
.A2(n_387),
.B1(n_388),
.B2(n_390),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_318),
.B(n_272),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_384),
.B(n_389),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_351),
.A2(n_300),
.B1(n_314),
.B2(n_318),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_326),
.A2(n_213),
.B1(n_229),
.B2(n_291),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_339),
.B(n_230),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_352),
.A2(n_265),
.B1(n_294),
.B2(n_246),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_314),
.A2(n_248),
.B1(n_226),
.B2(n_234),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_391),
.A2(n_306),
.B1(n_337),
.B2(n_327),
.Y(n_420)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_308),
.Y(n_392)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_392),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_316),
.B(n_232),
.C(n_293),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_395),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_315),
.B(n_226),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_394),
.B(n_399),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_348),
.B(n_324),
.C(n_335),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_334),
.B(n_255),
.C(n_234),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_397),
.B(n_403),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_344),
.A2(n_279),
.B1(n_275),
.B2(n_271),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_310),
.B(n_285),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_305),
.Y(n_400)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_400),
.Y(n_414)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_305),
.Y(n_401)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_401),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_304),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_402),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_344),
.B(n_285),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_336),
.B(n_202),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_404),
.B(n_353),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_388),
.A2(n_343),
.B1(n_349),
.B2(n_354),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_405),
.A2(n_401),
.B(n_378),
.Y(n_475)
);

NAND3xp33_ASAP7_75t_L g445 ( 
.A(n_407),
.B(n_369),
.C(n_360),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_362),
.A2(n_372),
.B(n_366),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_409),
.A2(n_421),
.B(n_429),
.Y(n_472)
);

O2A1O1Ixp33_ASAP7_75t_L g458 ( 
.A1(n_415),
.A2(n_431),
.B(n_437),
.C(n_405),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_420),
.B(n_440),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_382),
.A2(n_307),
.B(n_349),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_394),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_422),
.B(n_376),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_388),
.A2(n_309),
.B(n_319),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_423),
.A2(n_431),
.B(n_435),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_383),
.B(n_309),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_403),
.C(n_395),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_361),
.A2(n_325),
.B1(n_343),
.B2(n_347),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_426),
.A2(n_427),
.B1(n_440),
.B2(n_371),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_361),
.A2(n_325),
.B1(n_354),
.B2(n_308),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_377),
.A2(n_350),
.B(n_355),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_374),
.A2(n_327),
.B1(n_306),
.B2(n_355),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_430),
.A2(n_439),
.B1(n_380),
.B2(n_375),
.Y(n_450)
);

AO21x1_ASAP7_75t_L g431 ( 
.A1(n_363),
.A2(n_346),
.B(n_342),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_368),
.Y(n_433)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_433),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_SL g435 ( 
.A1(n_404),
.A2(n_302),
.B1(n_350),
.B2(n_330),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_367),
.A2(n_322),
.B1(n_311),
.B2(n_323),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_385),
.A2(n_322),
.B1(n_311),
.B2(n_323),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_368),
.Y(n_441)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_441),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_364),
.Y(n_456)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_443),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_369),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_444),
.B(n_462),
.C(n_470),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_445),
.A2(n_458),
.B(n_474),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_432),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_447),
.B(n_453),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_448),
.B(n_406),
.Y(n_483)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_450),
.Y(n_488)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_451),
.Y(n_497)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_433),
.Y(n_452)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_452),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_413),
.A2(n_365),
.B1(n_390),
.B2(n_391),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_434),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_454),
.Y(n_484)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_441),
.Y(n_455)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_455),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_SL g485 ( 
.A(n_456),
.B(n_476),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_413),
.A2(n_365),
.B1(n_387),
.B2(n_398),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_457),
.B(n_465),
.Y(n_507)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_459),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_432),
.B(n_393),
.Y(n_461)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_461),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_436),
.B(n_397),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_411),
.B(n_396),
.Y(n_463)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_463),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_409),
.A2(n_416),
.B1(n_410),
.B2(n_421),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_464),
.A2(n_466),
.B1(n_467),
.B2(n_477),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_426),
.A2(n_365),
.B1(n_376),
.B2(n_396),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_427),
.A2(n_375),
.B1(n_380),
.B2(n_386),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_410),
.A2(n_386),
.B1(n_381),
.B2(n_402),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_438),
.B(n_301),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_468),
.B(n_471),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_419),
.Y(n_469)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_469),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_436),
.B(n_331),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_419),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_411),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_473),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_407),
.A2(n_373),
.B(n_400),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_475),
.A2(n_423),
.B(n_431),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_418),
.B(n_379),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_415),
.A2(n_392),
.B1(n_320),
.B2(n_331),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_478),
.Y(n_529)
);

NOR2x1_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_418),
.Y(n_480)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_480),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_448),
.B(n_406),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_482),
.B(n_486),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_483),
.B(n_495),
.C(n_496),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_442),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_459),
.Y(n_489)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_489),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_464),
.A2(n_415),
.B1(n_422),
.B2(n_417),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_494),
.A2(n_435),
.B1(n_420),
.B2(n_446),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_470),
.B(n_442),
.C(n_416),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_444),
.B(n_415),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_461),
.B(n_472),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_498),
.B(n_502),
.C(n_504),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_472),
.B(n_463),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_474),
.B(n_476),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_473),
.B(n_412),
.C(n_439),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_505),
.B(n_508),
.C(n_467),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_465),
.B(n_412),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_466),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_509),
.Y(n_526)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_481),
.Y(n_511)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_511),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_486),
.B(n_447),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_514),
.B(n_521),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_487),
.A2(n_457),
.B1(n_453),
.B2(n_443),
.Y(n_515)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_515),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_482),
.B(n_458),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_516),
.B(n_522),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_417),
.Y(n_517)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_517),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_487),
.A2(n_499),
.B1(n_493),
.B2(n_507),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_519),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_SL g521 ( 
.A(n_498),
.B(n_477),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_483),
.B(n_475),
.Y(n_522)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_479),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_524),
.B(n_525),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_499),
.A2(n_451),
.B1(n_460),
.B2(n_430),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_527),
.B(n_533),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_SL g528 ( 
.A(n_485),
.B(n_450),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_528),
.B(n_539),
.Y(n_545)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_510),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_530),
.Y(n_547)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_506),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_531),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_492),
.B(n_460),
.C(n_455),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_532),
.B(n_538),
.C(n_485),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_501),
.B(n_452),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_534),
.A2(n_508),
.B1(n_504),
.B2(n_488),
.Y(n_552)
);

CKINVDCx16_ASAP7_75t_R g535 ( 
.A(n_505),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_535),
.Y(n_544)
);

INVxp33_ASAP7_75t_L g536 ( 
.A(n_484),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_536),
.A2(n_517),
.B(n_512),
.Y(n_549)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_491),
.Y(n_537)
);

BUFx24_ASAP7_75t_SL g555 ( 
.A(n_537),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_492),
.B(n_449),
.C(n_446),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_495),
.B(n_449),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_541),
.B(n_522),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_538),
.B(n_490),
.C(n_502),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_542),
.B(n_546),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_518),
.B(n_520),
.C(n_539),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_527),
.A2(n_493),
.B1(n_507),
.B2(n_488),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_548),
.A2(n_528),
.B1(n_533),
.B2(n_514),
.Y(n_579)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_549),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_552),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_534),
.A2(n_497),
.B1(n_494),
.B2(n_503),
.Y(n_557)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_557),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_529),
.A2(n_478),
.B(n_503),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_558),
.A2(n_554),
.B(n_557),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_518),
.B(n_496),
.C(n_497),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_560),
.B(n_562),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_520),
.B(n_408),
.C(n_480),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_558),
.A2(n_529),
.B(n_526),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_563),
.B(n_575),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_565),
.B(n_568),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_561),
.B(n_513),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_567),
.B(n_578),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_556),
.B(n_511),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_542),
.B(n_532),
.C(n_523),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_571),
.B(n_576),
.C(n_581),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_540),
.B(n_523),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_573),
.B(n_574),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_556),
.B(n_560),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_SL g575 ( 
.A1(n_544),
.A2(n_521),
.B(n_512),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_546),
.B(n_541),
.C(n_562),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_540),
.B(n_516),
.Y(n_577)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_577),
.B(n_579),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_555),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_SL g596 ( 
.A1(n_580),
.A2(n_570),
.B(n_579),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_545),
.B(n_429),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_569),
.A2(n_553),
.B1(n_559),
.B2(n_551),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_582),
.B(n_583),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_564),
.B(n_548),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_569),
.A2(n_559),
.B1(n_544),
.B2(n_552),
.Y(n_584)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_584),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_572),
.A2(n_550),
.B1(n_547),
.B2(n_549),
.Y(n_587)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_587),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_572),
.A2(n_543),
.B1(n_545),
.B2(n_536),
.Y(n_589)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_589),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_574),
.B(n_408),
.Y(n_590)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_590),
.Y(n_604)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_563),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_591),
.B(n_594),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_580),
.B(n_543),
.Y(n_593)
);

CKINVDCx14_ASAP7_75t_R g601 ( 
.A(n_593),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_570),
.B(n_434),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_L g609 ( 
.A1(n_596),
.A2(n_454),
.B(n_414),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_586),
.B(n_576),
.C(n_573),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_600),
.B(n_605),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_595),
.B(n_566),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_L g606 ( 
.A1(n_585),
.A2(n_571),
.B(n_575),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_606),
.B(n_592),
.Y(n_614)
);

OA21x2_ASAP7_75t_L g607 ( 
.A1(n_585),
.A2(n_577),
.B(n_581),
.Y(n_607)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_607),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_596),
.A2(n_565),
.B(n_428),
.Y(n_608)
);

NAND3xp33_ASAP7_75t_SL g620 ( 
.A(n_608),
.B(n_428),
.C(n_424),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_609),
.B(n_414),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_601),
.A2(n_593),
.B1(n_586),
.B2(n_589),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_611),
.A2(n_603),
.B(n_610),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_SL g612 ( 
.A1(n_602),
.A2(n_588),
.B1(n_593),
.B2(n_592),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_612),
.B(n_615),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_SL g626 ( 
.A1(n_614),
.A2(n_598),
.B(n_604),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_600),
.B(n_597),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_599),
.B(n_597),
.Y(n_617)
);

O2A1O1Ixp33_ASAP7_75t_SL g624 ( 
.A1(n_617),
.A2(n_620),
.B(n_608),
.C(n_609),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_618),
.B(n_619),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_605),
.B(n_434),
.Y(n_619)
);

NAND4xp25_ASAP7_75t_L g628 ( 
.A(n_622),
.B(n_624),
.C(n_625),
.D(n_616),
.Y(n_628)
);

INVx6_ASAP7_75t_L g625 ( 
.A(n_613),
.Y(n_625)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_626),
.B(n_611),
.Y(n_627)
);

NOR3xp33_ASAP7_75t_L g632 ( 
.A(n_627),
.B(n_628),
.C(n_630),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_623),
.B(n_617),
.C(n_607),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_SL g631 ( 
.A1(n_629),
.A2(n_424),
.B(n_353),
.Y(n_631)
);

NOR3xp33_ASAP7_75t_SL g630 ( 
.A(n_621),
.B(n_607),
.C(n_620),
.Y(n_630)
);

NOR3xp33_ASAP7_75t_L g633 ( 
.A(n_631),
.B(n_630),
.C(n_320),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_633),
.B(n_632),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_634),
.B(n_297),
.C(n_330),
.Y(n_635)
);

BUFx24_ASAP7_75t_SL g636 ( 
.A(n_635),
.Y(n_636)
);


endmodule