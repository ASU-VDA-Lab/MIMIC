module real_aes_8409_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g106 ( .A(n_0), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_1), .A2(n_129), .B(n_133), .C(n_214), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_2), .A2(n_163), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g508 ( .A(n_3), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_4), .B(n_230), .Y(n_249) );
AOI21xp33_ASAP7_75t_L g473 ( .A1(n_5), .A2(n_163), .B(n_474), .Y(n_473) );
AND2x6_ASAP7_75t_L g129 ( .A(n_6), .B(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g204 ( .A(n_7), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_8), .B(n_42), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_8), .B(n_42), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_9), .A2(n_162), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_10), .B(n_141), .Y(n_216) );
INVx1_ASAP7_75t_L g478 ( .A(n_11), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_12), .B(n_244), .Y(n_533) );
INVx1_ASAP7_75t_L g149 ( .A(n_13), .Y(n_149) );
INVx1_ASAP7_75t_L g545 ( .A(n_14), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_15), .A2(n_139), .B(n_226), .C(n_228), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_16), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_17), .B(n_496), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_18), .B(n_163), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_19), .B(n_175), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_20), .A2(n_244), .B(n_259), .C(n_261), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_21), .B(n_230), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_22), .B(n_141), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_23), .A2(n_171), .B(n_228), .C(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_24), .B(n_141), .Y(n_140) );
CKINVDCx16_ASAP7_75t_R g180 ( .A(n_25), .Y(n_180) );
INVx1_ASAP7_75t_L g137 ( .A(n_26), .Y(n_137) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_27), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_28), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_29), .B(n_141), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_30), .A2(n_31), .B1(n_740), .B2(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_30), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_31), .Y(n_740) );
INVx1_ASAP7_75t_L g169 ( .A(n_32), .Y(n_169) );
INVx1_ASAP7_75t_L g487 ( .A(n_33), .Y(n_487) );
AOI222xp33_ASAP7_75t_L g456 ( .A1(n_34), .A2(n_457), .B1(n_739), .B2(n_742), .C1(n_745), .C2(n_746), .Y(n_456) );
INVx2_ASAP7_75t_L g127 ( .A(n_35), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_36), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_37), .A2(n_244), .B(n_245), .C(n_247), .Y(n_243) );
INVxp67_ASAP7_75t_L g170 ( .A(n_38), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g132 ( .A1(n_39), .A2(n_133), .B(n_136), .C(n_144), .Y(n_132) );
CKINVDCx14_ASAP7_75t_R g242 ( .A(n_40), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_41), .A2(n_129), .B(n_133), .C(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g486 ( .A(n_43), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_44), .A2(n_188), .B(n_202), .C(n_203), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_45), .B(n_141), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_46), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_47), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_48), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g257 ( .A(n_49), .Y(n_257) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_50), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_51), .A2(n_102), .B1(n_110), .B2(n_751), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_52), .B(n_163), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_53), .A2(n_133), .B1(n_261), .B2(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_54), .Y(n_524) );
CKINVDCx16_ASAP7_75t_R g505 ( .A(n_55), .Y(n_505) );
CKINVDCx14_ASAP7_75t_R g200 ( .A(n_56), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_57), .A2(n_202), .B(n_247), .C(n_477), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_58), .Y(n_561) );
INVx1_ASAP7_75t_L g475 ( .A(n_59), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_60), .A2(n_88), .B1(n_443), .B2(n_444), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_60), .Y(n_444) );
INVx1_ASAP7_75t_L g130 ( .A(n_61), .Y(n_130) );
INVx1_ASAP7_75t_L g148 ( .A(n_62), .Y(n_148) );
INVx1_ASAP7_75t_SL g246 ( .A(n_63), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_64), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_65), .B(n_230), .Y(n_263) );
INVx1_ASAP7_75t_L g183 ( .A(n_66), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_SL g495 ( .A1(n_67), .A2(n_247), .B(n_496), .C(n_497), .Y(n_495) );
INVxp67_ASAP7_75t_L g498 ( .A(n_68), .Y(n_498) );
INVx1_ASAP7_75t_L g109 ( .A(n_69), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_70), .A2(n_163), .B(n_199), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_71), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_72), .A2(n_163), .B(n_223), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_73), .Y(n_490) );
INVx1_ASAP7_75t_L g555 ( .A(n_74), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_75), .A2(n_162), .B(n_164), .Y(n_161) );
CKINVDCx16_ASAP7_75t_R g131 ( .A(n_76), .Y(n_131) );
INVx1_ASAP7_75t_L g224 ( .A(n_77), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g556 ( .A1(n_78), .A2(n_129), .B(n_133), .C(n_557), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_79), .A2(n_163), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g227 ( .A(n_80), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_81), .B(n_138), .Y(n_521) );
INVx2_ASAP7_75t_L g146 ( .A(n_82), .Y(n_146) );
INVx1_ASAP7_75t_L g215 ( .A(n_83), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_84), .B(n_496), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_85), .A2(n_129), .B(n_133), .C(n_507), .Y(n_506) );
NAND3xp33_ASAP7_75t_SL g105 ( .A(n_86), .B(n_106), .C(n_107), .Y(n_105) );
OR2x2_ASAP7_75t_L g447 ( .A(n_86), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g460 ( .A(n_86), .B(n_449), .Y(n_460) );
INVx2_ASAP7_75t_L g464 ( .A(n_86), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_87), .A2(n_133), .B(n_182), .C(n_190), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_88), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_89), .B(n_145), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_90), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_91), .A2(n_129), .B(n_133), .C(n_531), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_92), .Y(n_537) );
INVx1_ASAP7_75t_L g494 ( .A(n_93), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g542 ( .A(n_94), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_95), .B(n_138), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_96), .B(n_153), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_97), .B(n_153), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_98), .B(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g260 ( .A(n_99), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_100), .A2(n_163), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
BUFx2_ASAP7_75t_L g751 ( .A(n_103), .Y(n_751) );
OR2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
AND2x2_ASAP7_75t_L g449 ( .A(n_106), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
AO21x2_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_115), .B(n_455), .Y(n_110) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g750 ( .A(n_114), .Y(n_750) );
OAI21xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_445), .B(n_451), .Y(n_115) );
XOR2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_442), .Y(n_116) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_117), .A2(n_458), .B1(n_461), .B2(n_465), .Y(n_457) );
INVx1_ASAP7_75t_L g743 ( .A(n_117), .Y(n_743) );
OR4x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_332), .C(n_379), .D(n_419), .Y(n_117) );
NAND3xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_278), .C(n_307), .Y(n_118) );
AOI211xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_193), .B(n_231), .C(n_271), .Y(n_119) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_120), .A2(n_291), .B(n_308), .C(n_312), .Y(n_307) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_155), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_122), .B(n_270), .Y(n_269) );
INVx3_ASAP7_75t_SL g274 ( .A(n_122), .Y(n_274) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_122), .Y(n_286) );
AND2x4_ASAP7_75t_L g290 ( .A(n_122), .B(n_238), .Y(n_290) );
AND2x2_ASAP7_75t_L g301 ( .A(n_122), .B(n_178), .Y(n_301) );
OR2x2_ASAP7_75t_L g325 ( .A(n_122), .B(n_234), .Y(n_325) );
AND2x2_ASAP7_75t_L g338 ( .A(n_122), .B(n_239), .Y(n_338) );
AND2x2_ASAP7_75t_L g378 ( .A(n_122), .B(n_364), .Y(n_378) );
AND2x2_ASAP7_75t_L g385 ( .A(n_122), .B(n_348), .Y(n_385) );
AND2x2_ASAP7_75t_L g415 ( .A(n_122), .B(n_156), .Y(n_415) );
OR2x6_ASAP7_75t_L g122 ( .A(n_123), .B(n_150), .Y(n_122) );
O2A1O1Ixp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_131), .B(n_132), .C(n_145), .Y(n_123) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_124), .A2(n_180), .B(n_181), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_124), .A2(n_212), .B(n_213), .Y(n_211) );
OAI22xp33_ASAP7_75t_L g483 ( .A1(n_124), .A2(n_173), .B1(n_484), .B2(n_488), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_124), .A2(n_505), .B(n_506), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_124), .A2(n_555), .B(n_556), .Y(n_554) );
NAND2x1p5_ASAP7_75t_L g124 ( .A(n_125), .B(n_129), .Y(n_124) );
AND2x4_ASAP7_75t_L g163 ( .A(n_125), .B(n_129), .Y(n_163) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_128), .Y(n_125) );
INVx1_ASAP7_75t_L g143 ( .A(n_126), .Y(n_143) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g134 ( .A(n_127), .Y(n_134) );
INVx1_ASAP7_75t_L g262 ( .A(n_127), .Y(n_262) );
INVx1_ASAP7_75t_L g135 ( .A(n_128), .Y(n_135) );
INVx3_ASAP7_75t_L g139 ( .A(n_128), .Y(n_139) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_128), .Y(n_141) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_128), .Y(n_172) );
INVx1_ASAP7_75t_L g496 ( .A(n_128), .Y(n_496) );
BUFx3_ASAP7_75t_L g144 ( .A(n_129), .Y(n_144) );
INVx4_ASAP7_75t_SL g173 ( .A(n_129), .Y(n_173) );
INVx5_ASAP7_75t_L g166 ( .A(n_133), .Y(n_166) );
AND2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
BUFx3_ASAP7_75t_L g189 ( .A(n_134), .Y(n_189) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_134), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B(n_140), .C(n_142), .Y(n_136) );
OAI22xp33_ASAP7_75t_L g168 ( .A1(n_138), .A2(n_169), .B1(n_170), .B2(n_171), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_138), .A2(n_508), .B(n_509), .C(n_510), .Y(n_507) );
INVx5_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_139), .B(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_139), .B(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_139), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g202 ( .A(n_141), .Y(n_202) );
INVx4_ASAP7_75t_L g244 ( .A(n_141), .Y(n_244) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_143), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g176 ( .A(n_145), .Y(n_176) );
OA21x2_ASAP7_75t_L g197 ( .A1(n_145), .A2(n_198), .B(n_205), .Y(n_197) );
INVx1_ASAP7_75t_L g210 ( .A(n_145), .Y(n_210) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_145), .A2(n_540), .B(n_546), .Y(n_539) );
AND2x2_ASAP7_75t_SL g145 ( .A(n_146), .B(n_147), .Y(n_145) );
AND2x2_ASAP7_75t_L g154 ( .A(n_146), .B(n_147), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_152), .A2(n_179), .B(n_191), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_152), .B(n_218), .Y(n_217) );
INVx3_ASAP7_75t_L g230 ( .A(n_152), .Y(n_230) );
NOR2xp33_ASAP7_75t_SL g523 ( .A(n_152), .B(n_524), .Y(n_523) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_153), .Y(n_221) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_153), .A2(n_492), .B(n_499), .Y(n_491) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g160 ( .A(n_154), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_155), .B(n_342), .Y(n_354) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_177), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_156), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g292 ( .A(n_156), .B(n_177), .Y(n_292) );
BUFx3_ASAP7_75t_L g300 ( .A(n_156), .Y(n_300) );
OR2x2_ASAP7_75t_L g321 ( .A(n_156), .B(n_196), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_156), .B(n_342), .Y(n_432) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_161), .B(n_174), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_158), .A2(n_235), .B(n_236), .Y(n_234) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_158), .A2(n_554), .B(n_560), .Y(n_553) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_SL g517 ( .A1(n_159), .A2(n_518), .B(n_519), .Y(n_517) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_160), .A2(n_483), .B(n_489), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_160), .B(n_490), .Y(n_489) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_160), .A2(n_504), .B(n_511), .Y(n_503) );
INVx1_ASAP7_75t_L g235 ( .A(n_161), .Y(n_235) );
BUFx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_SL g164 ( .A1(n_165), .A2(n_166), .B(n_167), .C(n_173), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_SL g199 ( .A1(n_166), .A2(n_173), .B(n_200), .C(n_201), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_SL g223 ( .A1(n_166), .A2(n_173), .B(n_224), .C(n_225), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_166), .A2(n_173), .B(n_242), .C(n_243), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_SL g256 ( .A1(n_166), .A2(n_173), .B(n_257), .C(n_258), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_L g474 ( .A1(n_166), .A2(n_173), .B(n_475), .C(n_476), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_166), .A2(n_173), .B(n_494), .C(n_495), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_166), .A2(n_173), .B(n_542), .C(n_543), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_171), .B(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_171), .B(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_171), .B(n_545), .Y(n_544) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g185 ( .A(n_172), .Y(n_185) );
OAI22xp5_ASAP7_75t_SL g485 ( .A1(n_172), .A2(n_185), .B1(n_486), .B2(n_487), .Y(n_485) );
INVx1_ASAP7_75t_L g190 ( .A(n_173), .Y(n_190) );
INVx1_ASAP7_75t_L g236 ( .A(n_174), .Y(n_236) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_176), .B(n_192), .Y(n_191) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_176), .A2(n_529), .B(n_536), .Y(n_528) );
AND2x2_ASAP7_75t_L g237 ( .A(n_177), .B(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g285 ( .A(n_177), .Y(n_285) );
AND2x2_ASAP7_75t_L g348 ( .A(n_177), .B(n_239), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g350 ( .A1(n_177), .A2(n_351), .B1(n_353), .B2(n_355), .C(n_356), .Y(n_350) );
AND2x2_ASAP7_75t_L g364 ( .A(n_177), .B(n_234), .Y(n_364) );
AND2x2_ASAP7_75t_L g390 ( .A(n_177), .B(n_274), .Y(n_390) );
INVx2_ASAP7_75t_SL g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g270 ( .A(n_178), .B(n_239), .Y(n_270) );
BUFx2_ASAP7_75t_L g404 ( .A(n_178), .Y(n_404) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_186), .C(n_187), .Y(n_182) );
O2A1O1Ixp5_ASAP7_75t_L g214 ( .A1(n_184), .A2(n_187), .B(n_215), .C(n_216), .Y(n_214) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_187), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_187), .A2(n_558), .B(n_559), .Y(n_557) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g228 ( .A(n_189), .Y(n_228) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
OAI32xp33_ASAP7_75t_L g370 ( .A1(n_194), .A2(n_331), .A3(n_345), .B1(n_371), .B2(n_372), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_195), .B(n_206), .Y(n_194) );
AND2x2_ASAP7_75t_L g311 ( .A(n_195), .B(n_253), .Y(n_311) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
OR2x2_ASAP7_75t_L g293 ( .A(n_196), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_196), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g365 ( .A(n_196), .B(n_253), .Y(n_365) );
AND2x2_ASAP7_75t_L g376 ( .A(n_196), .B(n_268), .Y(n_376) );
BUFx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OR2x2_ASAP7_75t_L g277 ( .A(n_197), .B(n_254), .Y(n_277) );
AND2x2_ASAP7_75t_L g281 ( .A(n_197), .B(n_254), .Y(n_281) );
AND2x2_ASAP7_75t_L g316 ( .A(n_197), .B(n_267), .Y(n_316) );
AND2x2_ASAP7_75t_L g323 ( .A(n_197), .B(n_219), .Y(n_323) );
OAI211xp5_ASAP7_75t_L g328 ( .A1(n_197), .A2(n_274), .B(n_285), .C(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g382 ( .A(n_197), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_197), .B(n_208), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_206), .B(n_265), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_206), .B(n_281), .Y(n_371) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OR2x2_ASAP7_75t_L g276 ( .A(n_207), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_219), .Y(n_207) );
AND2x2_ASAP7_75t_L g268 ( .A(n_208), .B(n_220), .Y(n_268) );
OR2x2_ASAP7_75t_L g283 ( .A(n_208), .B(n_220), .Y(n_283) );
AND2x2_ASAP7_75t_L g306 ( .A(n_208), .B(n_267), .Y(n_306) );
INVx1_ASAP7_75t_L g310 ( .A(n_208), .Y(n_310) );
AND2x2_ASAP7_75t_L g329 ( .A(n_208), .B(n_266), .Y(n_329) );
OAI22xp33_ASAP7_75t_L g339 ( .A1(n_208), .A2(n_294), .B1(n_340), .B2(n_341), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_208), .B(n_382), .Y(n_406) );
AND2x2_ASAP7_75t_L g421 ( .A(n_208), .B(n_281), .Y(n_421) );
INVx4_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
BUFx3_ASAP7_75t_L g251 ( .A(n_209), .Y(n_251) );
AND2x2_ASAP7_75t_L g295 ( .A(n_209), .B(n_220), .Y(n_295) );
AND2x2_ASAP7_75t_L g297 ( .A(n_209), .B(n_253), .Y(n_297) );
AND3x2_ASAP7_75t_L g359 ( .A(n_209), .B(n_323), .C(n_360), .Y(n_359) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_217), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_210), .B(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_210), .B(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_210), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g394 ( .A(n_219), .B(n_266), .Y(n_394) );
INVx1_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g253 ( .A(n_220), .B(n_254), .Y(n_253) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_220), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_220), .B(n_265), .Y(n_327) );
NAND3xp33_ASAP7_75t_L g434 ( .A(n_220), .B(n_306), .C(n_382), .Y(n_434) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_229), .Y(n_220) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_221), .A2(n_240), .B(n_249), .Y(n_239) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_221), .A2(n_255), .B(n_263), .Y(n_254) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_230), .A2(n_473), .B(n_479), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_250), .B1(n_264), .B2(n_269), .Y(n_231) );
INVx1_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_237), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_234), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_SL g346 ( .A(n_234), .Y(n_346) );
OAI31xp33_ASAP7_75t_L g362 ( .A1(n_237), .A2(n_363), .A3(n_364), .B(n_365), .Y(n_362) );
AND2x2_ASAP7_75t_L g387 ( .A(n_237), .B(n_274), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_237), .B(n_300), .Y(n_433) );
AND2x2_ASAP7_75t_L g342 ( .A(n_238), .B(n_274), .Y(n_342) );
AND2x2_ASAP7_75t_L g403 ( .A(n_238), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g273 ( .A(n_239), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g331 ( .A(n_239), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_244), .B(n_246), .Y(n_245) );
INVx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_248), .Y(n_534) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
CKINVDCx16_ASAP7_75t_R g352 ( .A(n_251), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_252), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
AOI221x1_ASAP7_75t_SL g319 ( .A1(n_253), .A2(n_320), .B1(n_322), .B2(n_324), .C(n_326), .Y(n_319) );
INVx2_ASAP7_75t_L g267 ( .A(n_254), .Y(n_267) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_254), .Y(n_361) );
INVx2_ASAP7_75t_L g510 ( .A(n_261), .Y(n_510) );
INVx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g349 ( .A(n_264), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_265), .B(n_282), .Y(n_374) );
INVx1_ASAP7_75t_SL g437 ( .A(n_265), .Y(n_437) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g355 ( .A(n_268), .B(n_281), .Y(n_355) );
INVx1_ASAP7_75t_L g423 ( .A(n_269), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_269), .B(n_352), .Y(n_436) );
INVx2_ASAP7_75t_SL g275 ( .A(n_270), .Y(n_275) );
AND2x2_ASAP7_75t_L g318 ( .A(n_270), .B(n_274), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_270), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_270), .B(n_345), .Y(n_372) );
AOI21xp33_ASAP7_75t_SL g271 ( .A1(n_272), .A2(n_275), .B(n_276), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_273), .B(n_345), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_273), .B(n_300), .Y(n_441) );
OR2x2_ASAP7_75t_L g313 ( .A(n_274), .B(n_292), .Y(n_313) );
AND2x2_ASAP7_75t_L g412 ( .A(n_274), .B(n_403), .Y(n_412) );
OAI22xp5_ASAP7_75t_SL g287 ( .A1(n_275), .A2(n_288), .B1(n_293), .B2(n_296), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_275), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g335 ( .A(n_277), .B(n_283), .Y(n_335) );
INVx1_ASAP7_75t_L g399 ( .A(n_277), .Y(n_399) );
AOI311xp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_284), .A3(n_286), .B(n_287), .C(n_298), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_282), .A2(n_414), .B1(n_426), .B2(n_429), .C(n_431), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_282), .B(n_437), .Y(n_439) );
INVx2_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g336 ( .A(n_284), .Y(n_336) );
AOI211xp5_ASAP7_75t_L g326 ( .A1(n_285), .A2(n_327), .B(n_328), .C(n_330), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_SL g395 ( .A1(n_289), .A2(n_291), .B(n_396), .C(n_397), .Y(n_395) );
INVx3_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_290), .B(n_364), .Y(n_430) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
OAI221xp5_ASAP7_75t_L g312 ( .A1(n_293), .A2(n_313), .B1(n_314), .B2(n_317), .C(n_319), .Y(n_312) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g315 ( .A(n_295), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g398 ( .A(n_295), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_302), .Y(n_298) );
A2O1A1Ixp33_ASAP7_75t_L g356 ( .A1(n_299), .A2(n_357), .B(n_358), .C(n_362), .Y(n_356) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_300), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_300), .B(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g322 ( .A(n_306), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_310), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g424 ( .A(n_313), .Y(n_424) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_316), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g351 ( .A(n_316), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_SL g428 ( .A(n_316), .Y(n_428) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g369 ( .A(n_318), .B(n_345), .Y(n_369) );
INVx1_ASAP7_75t_SL g363 ( .A(n_325), .Y(n_363) );
INVx1_ASAP7_75t_L g340 ( .A(n_331), .Y(n_340) );
NAND3xp33_ASAP7_75t_SL g332 ( .A(n_333), .B(n_350), .C(n_366), .Y(n_332) );
AOI322xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .A3(n_337), .B1(n_339), .B2(n_343), .C1(n_347), .C2(n_349), .Y(n_333) );
AOI211xp5_ASAP7_75t_L g386 ( .A1(n_334), .A2(n_387), .B(n_388), .C(n_395), .Y(n_386) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_337), .A2(n_358), .B1(n_389), .B2(n_391), .Y(n_388) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g347 ( .A(n_345), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g384 ( .A(n_345), .B(n_385), .Y(n_384) );
AOI32xp33_ASAP7_75t_L g435 ( .A1(n_345), .A2(n_436), .A3(n_437), .B1(n_438), .B2(n_440), .Y(n_435) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g357 ( .A(n_348), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_348), .A2(n_401), .B1(n_405), .B2(n_407), .C(n_410), .Y(n_400) );
AND2x2_ASAP7_75t_L g414 ( .A(n_348), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g417 ( .A(n_352), .B(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g427 ( .A(n_352), .B(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g418 ( .A(n_361), .B(n_382), .Y(n_418) );
AOI211xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B(n_370), .C(n_373), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI21xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B(n_377), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI211xp5_ASAP7_75t_SL g379 ( .A1(n_380), .A2(n_383), .B(n_386), .C(n_400), .Y(n_379) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_394), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g409 ( .A(n_406), .Y(n_409) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AOI21xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .B(n_416), .Y(n_410) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI211xp5_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_422), .B(n_425), .C(n_435), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_421), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx2_ASAP7_75t_L g454 ( .A(n_447), .Y(n_454) );
NOR2x2_ASAP7_75t_L g748 ( .A(n_448), .B(n_464), .Y(n_748) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g463 ( .A(n_449), .B(n_464), .Y(n_463) );
AOI21xp33_ASAP7_75t_L g455 ( .A1(n_451), .A2(n_456), .B(n_749), .Y(n_455) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI22x1_ASAP7_75t_L g742 ( .A1(n_458), .A2(n_461), .B1(n_743), .B2(n_744), .Y(n_742) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVxp67_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g744 ( .A(n_466), .Y(n_744) );
BUFx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND3x1_ASAP7_75t_L g467 ( .A(n_468), .B(n_661), .C(n_706), .Y(n_467) );
NOR4xp25_ASAP7_75t_L g468 ( .A(n_469), .B(n_584), .C(n_625), .D(n_642), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_500), .B(n_514), .C(n_547), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_480), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_471), .B(n_501), .Y(n_500) );
NOR4xp25_ASAP7_75t_L g608 ( .A(n_471), .B(n_602), .C(n_609), .D(n_615), .Y(n_608) );
AND2x2_ASAP7_75t_L g681 ( .A(n_471), .B(n_570), .Y(n_681) );
AND2x2_ASAP7_75t_L g700 ( .A(n_471), .B(n_646), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_471), .B(n_695), .Y(n_709) );
AND2x2_ASAP7_75t_L g722 ( .A(n_471), .B(n_513), .Y(n_722) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_SL g567 ( .A(n_472), .Y(n_567) );
AND2x2_ASAP7_75t_L g574 ( .A(n_472), .B(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g624 ( .A(n_472), .B(n_481), .Y(n_624) );
AND2x2_ASAP7_75t_SL g635 ( .A(n_472), .B(n_570), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_472), .B(n_481), .Y(n_639) );
AND2x2_ASAP7_75t_L g648 ( .A(n_472), .B(n_573), .Y(n_648) );
BUFx2_ASAP7_75t_L g671 ( .A(n_472), .Y(n_671) );
AND2x2_ASAP7_75t_L g675 ( .A(n_472), .B(n_491), .Y(n_675) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_491), .Y(n_480) );
AND2x2_ASAP7_75t_L g513 ( .A(n_481), .B(n_491), .Y(n_513) );
BUFx2_ASAP7_75t_L g577 ( .A(n_481), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_481), .A2(n_610), .B1(n_612), .B2(n_613), .Y(n_609) );
OR2x2_ASAP7_75t_L g631 ( .A(n_481), .B(n_503), .Y(n_631) );
AND2x2_ASAP7_75t_L g695 ( .A(n_481), .B(n_573), .Y(n_695) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g563 ( .A(n_482), .B(n_503), .Y(n_563) );
AND2x2_ASAP7_75t_L g570 ( .A(n_482), .B(n_491), .Y(n_570) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_482), .Y(n_612) );
OR2x2_ASAP7_75t_L g647 ( .A(n_482), .B(n_502), .Y(n_647) );
INVx1_ASAP7_75t_L g566 ( .A(n_491), .Y(n_566) );
INVx3_ASAP7_75t_L g575 ( .A(n_491), .Y(n_575) );
BUFx2_ASAP7_75t_L g599 ( .A(n_491), .Y(n_599) );
AND2x2_ASAP7_75t_L g632 ( .A(n_491), .B(n_567), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_500), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_717) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_513), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_502), .B(n_575), .Y(n_579) );
INVx1_ASAP7_75t_L g607 ( .A(n_502), .Y(n_607) );
INVx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx3_ASAP7_75t_L g573 ( .A(n_503), .Y(n_573) );
INVx1_ASAP7_75t_L g585 ( .A(n_513), .Y(n_585) );
NAND2x1_ASAP7_75t_SL g514 ( .A(n_515), .B(n_525), .Y(n_514) );
AND2x2_ASAP7_75t_L g583 ( .A(n_515), .B(n_538), .Y(n_583) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_515), .Y(n_657) );
AND2x2_ASAP7_75t_L g684 ( .A(n_515), .B(n_604), .Y(n_684) );
AND2x2_ASAP7_75t_L g692 ( .A(n_515), .B(n_654), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_515), .B(n_550), .Y(n_719) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g551 ( .A(n_516), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g568 ( .A(n_516), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g589 ( .A(n_516), .Y(n_589) );
INVx1_ASAP7_75t_L g595 ( .A(n_516), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_516), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g628 ( .A(n_516), .B(n_553), .Y(n_628) );
OR2x2_ASAP7_75t_L g666 ( .A(n_516), .B(n_621), .Y(n_666) );
AOI32xp33_ASAP7_75t_L g678 ( .A1(n_516), .A2(n_679), .A3(n_682), .B1(n_683), .B2(n_684), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_516), .B(n_654), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_516), .B(n_614), .Y(n_729) );
OR2x6_ASAP7_75t_L g516 ( .A(n_517), .B(n_523), .Y(n_516) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g640 ( .A(n_526), .B(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_538), .Y(n_526) );
INVx1_ASAP7_75t_L g602 ( .A(n_527), .Y(n_602) );
AND2x2_ASAP7_75t_L g604 ( .A(n_527), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_527), .B(n_552), .Y(n_621) );
AND2x2_ASAP7_75t_L g654 ( .A(n_527), .B(n_630), .Y(n_654) );
AND2x2_ASAP7_75t_L g691 ( .A(n_527), .B(n_553), .Y(n_691) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g550 ( .A(n_528), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_528), .B(n_552), .Y(n_581) );
AND2x2_ASAP7_75t_L g588 ( .A(n_528), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g629 ( .A(n_528), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_535), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B(n_534), .Y(n_531) );
INVx2_ASAP7_75t_L g605 ( .A(n_538), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_538), .B(n_552), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_538), .B(n_596), .Y(n_677) );
INVx1_ASAP7_75t_L g699 ( .A(n_538), .Y(n_699) );
INVx1_ASAP7_75t_L g716 ( .A(n_538), .Y(n_716) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g569 ( .A(n_539), .B(n_552), .Y(n_569) );
AND2x2_ASAP7_75t_L g591 ( .A(n_539), .B(n_553), .Y(n_591) );
INVx1_ASAP7_75t_L g630 ( .A(n_539), .Y(n_630) );
AOI221x1_ASAP7_75t_SL g547 ( .A1(n_548), .A2(n_562), .B1(n_568), .B2(n_570), .C(n_571), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_548), .A2(n_635), .B1(n_702), .B2(n_703), .Y(n_701) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_551), .Y(n_548) );
AND2x2_ASAP7_75t_L g593 ( .A(n_549), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g688 ( .A(n_549), .B(n_568), .Y(n_688) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g644 ( .A(n_550), .B(n_569), .Y(n_644) );
INVx1_ASAP7_75t_L g656 ( .A(n_551), .Y(n_656) );
AND2x2_ASAP7_75t_L g667 ( .A(n_551), .B(n_654), .Y(n_667) );
AND2x2_ASAP7_75t_L g734 ( .A(n_551), .B(n_629), .Y(n_734) );
INVx2_ASAP7_75t_L g596 ( .A(n_552), .Y(n_596) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_563), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g686 ( .A(n_563), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_564), .B(n_647), .Y(n_650) );
INVx3_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_565), .A2(n_686), .B(n_731), .Y(n_730) );
AND2x4_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NOR2xp33_ASAP7_75t_SL g708 ( .A(n_568), .B(n_594), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_569), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g660 ( .A(n_569), .B(n_588), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_569), .B(n_595), .Y(n_737) );
AND2x2_ASAP7_75t_L g606 ( .A(n_570), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g673 ( .A(n_570), .Y(n_673) );
AOI21xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_576), .B(n_580), .Y(n_571) );
NAND2x1_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_573), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g622 ( .A(n_573), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_SL g634 ( .A(n_573), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_573), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g658 ( .A(n_574), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_574), .B(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_574), .B(n_577), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
AOI211xp5_ASAP7_75t_L g645 ( .A1(n_577), .A2(n_616), .B(n_646), .C(n_648), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_577), .A2(n_664), .B1(n_667), .B2(n_668), .C(n_672), .Y(n_663) );
AND2x2_ASAP7_75t_L g659 ( .A(n_578), .B(n_612), .Y(n_659) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g619 ( .A(n_583), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g690 ( .A(n_583), .B(n_691), .Y(n_690) );
OAI211xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_586), .B(n_592), .C(n_617), .Y(n_584) );
NAND3xp33_ASAP7_75t_SL g703 ( .A(n_585), .B(n_704), .C(n_705), .Y(n_703) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .Y(n_586) );
OR2x2_ASAP7_75t_L g676 ( .A(n_587), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_597), .B1(n_600), .B2(n_606), .C(n_608), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_594), .B(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_594), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g616 ( .A(n_599), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_599), .A2(n_656), .B1(n_657), .B2(n_658), .Y(n_655) );
OR2x2_ASAP7_75t_L g736 ( .A(n_599), .B(n_647), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVxp67_ASAP7_75t_L g710 ( .A(n_602), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_604), .B(n_725), .Y(n_724) );
INVxp67_ASAP7_75t_L g611 ( .A(n_605), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_607), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_607), .B(n_654), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_607), .B(n_674), .Y(n_713) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_611), .Y(n_637) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g727 ( .A(n_616), .B(n_647), .Y(n_727) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_622), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g705 ( .A(n_622), .Y(n_705) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI322xp33_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_631), .A3(n_632), .B1(n_633), .B2(n_636), .C1(n_638), .C2(n_640), .Y(n_625) );
OAI322xp33_ASAP7_75t_L g707 ( .A1(n_626), .A2(n_708), .A3(n_709), .B1(n_710), .B2(n_711), .C1(n_712), .C2(n_714), .Y(n_707) );
CKINVDCx16_ASAP7_75t_R g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx4_ASAP7_75t_L g641 ( .A(n_628), .Y(n_641) );
AND2x2_ASAP7_75t_L g702 ( .A(n_628), .B(n_654), .Y(n_702) );
AND2x2_ASAP7_75t_L g715 ( .A(n_628), .B(n_716), .Y(n_715) );
CKINVDCx16_ASAP7_75t_R g726 ( .A(n_631), .Y(n_726) );
INVx1_ASAP7_75t_L g704 ( .A(n_632), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
OR2x2_ASAP7_75t_L g638 ( .A(n_634), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g721 ( .A(n_634), .B(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_634), .B(n_675), .Y(n_732) );
OR2x2_ASAP7_75t_L g665 ( .A(n_637), .B(n_666), .Y(n_665) );
INVxp33_ASAP7_75t_L g682 ( .A(n_637), .Y(n_682) );
OAI221xp5_ASAP7_75t_SL g642 ( .A1(n_641), .A2(n_643), .B1(n_645), .B2(n_649), .C(n_651), .Y(n_642) );
NOR2xp67_ASAP7_75t_L g698 ( .A(n_641), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g725 ( .A(n_641), .Y(n_725) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
INVx3_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
AOI322xp5_ASAP7_75t_L g689 ( .A1(n_648), .A2(n_673), .A3(n_690), .B1(n_692), .B2(n_693), .C1(n_696), .C2(n_700), .Y(n_689) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_655), .B1(n_659), .B2(n_660), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_685), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_663), .B(n_678), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_666), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
NAND2xp33_ASAP7_75t_SL g683 ( .A(n_669), .B(n_680), .Y(n_683) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
OAI322xp33_ASAP7_75t_L g723 ( .A1(n_671), .A2(n_724), .A3(n_726), .B1(n_727), .B2(n_728), .C1(n_730), .C2(n_733), .Y(n_723) );
AOI21xp33_ASAP7_75t_SL g672 ( .A1(n_673), .A2(n_674), .B(n_676), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_681), .B(n_729), .Y(n_738) );
OAI211xp5_ASAP7_75t_SL g685 ( .A1(n_686), .A2(n_687), .B(n_689), .C(n_701), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NOR4xp25_ASAP7_75t_L g706 ( .A(n_707), .B(n_717), .C(n_723), .D(n_735), .Y(n_706) );
INVxp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
CKINVDCx14_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
OAI21xp5_ASAP7_75t_SL g735 ( .A1(n_736), .A2(n_737), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g745 ( .A(n_739), .Y(n_745) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
endmodule