module real_jpeg_7225_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_0),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_0),
.B(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_0),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_0),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_0),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_0),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_0),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_1),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_1),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_1),
.B(n_186),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_1),
.B(n_339),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_1),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_1),
.B(n_389),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_1),
.B(n_62),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_2),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_2),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_2),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_2),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_3),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_3),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_3),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_3),
.B(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_3),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_3),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_3),
.B(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_4),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_4),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_4),
.Y(n_170)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_4),
.Y(n_180)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_4),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_5),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_5),
.B(n_80),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_5),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_5),
.B(n_312),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_5),
.B(n_325),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_5),
.B(n_70),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_5),
.B(n_384),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_5),
.B(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_6),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_6),
.B(n_192),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_6),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_6),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_6),
.B(n_293),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_6),
.B(n_186),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_6),
.B(n_376),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_6),
.B(n_188),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_7),
.Y(n_104)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_7),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_7),
.Y(n_142)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_9),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_9),
.Y(n_296)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_11),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_11),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_11),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_11),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g185 ( 
.A(n_11),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_11),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_11),
.B(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_12),
.Y(n_162)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_12),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_12),
.Y(n_328)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_14),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_14),
.B(n_142),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_14),
.B(n_310),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_14),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_14),
.B(n_74),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_14),
.B(n_392),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_14),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_15),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_15),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_15),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_15),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_15),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_15),
.B(n_183),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_15),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_15),
.B(n_373),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_16),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_16),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_16),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_16),
.B(n_172),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_16),
.B(n_330),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_16),
.B(n_347),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_16),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_17),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_17),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_17),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_17),
.B(n_117),
.Y(n_231)
);

AND2x2_ASAP7_75t_SL g289 ( 
.A(n_17),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_17),
.B(n_373),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_17),
.B(n_420),
.Y(n_419)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_125),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_123),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_105),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_28),
.B(n_105),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_90),
.C(n_91),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_29),
.A2(n_30),
.B1(n_528),
.B2(n_529),
.Y(n_527)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_60),
.C(n_77),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_31),
.A2(n_32),
.B1(n_508),
.B2(n_510),
.Y(n_507)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_43),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_34),
.B(n_38),
.C(n_43),
.Y(n_90)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_37),
.Y(n_147)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_41),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g390 ( 
.A(n_42),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_49),
.C(n_55),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_44),
.B(n_498),
.Y(n_497)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_49),
.A2(n_50),
.B1(n_55),
.B2(n_56),
.Y(n_498)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_54),
.Y(n_138)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_54),
.Y(n_226)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_59),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_59),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_60),
.A2(n_77),
.B1(n_78),
.B2(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_60),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.C(n_72),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_61),
.B(n_504),
.Y(n_503)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_65),
.A2(n_66),
.B1(n_202),
.B2(n_207),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_65),
.A2(n_66),
.B1(n_72),
.B2(n_73),
.Y(n_504)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_66),
.B(n_197),
.C(n_202),
.Y(n_505)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_71),
.Y(n_290)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_71),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_73),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_85),
.C(n_89),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_76),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_76),
.Y(n_340)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_76),
.Y(n_386)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_83),
.B1(n_84),
.B2(n_89),
.Y(n_78)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_82),
.Y(n_245)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_86),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_98),
.C(n_100),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_90),
.B(n_91),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_94),
.C(n_95),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_98),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_122),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_120),
.B2(n_121),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_526),
.B(n_531),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_491),
.B(n_523),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_298),
.B(n_490),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_253),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_129),
.B(n_253),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_194),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_130),
.B(n_195),
.C(n_232),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_167),
.C(n_176),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_131),
.B(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_143),
.C(n_157),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_132),
.B(n_476),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_136),
.C(n_139),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_138),
.B(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_SL g240 ( 
.A(n_142),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_143),
.A2(n_144),
.B1(n_157),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.C(n_153),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_145),
.B(n_153),
.Y(n_466)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_148),
.B(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_152),
.Y(n_415)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_156),
.Y(n_358)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_157),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_158),
.B(n_160),
.C(n_164),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_160),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g310 ( 
.A(n_162),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_162),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_163),
.B(n_202),
.C(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_163),
.A2(n_164),
.B1(n_202),
.B2(n_207),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_167),
.B(n_176),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_175),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_171),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_171),
.B(n_173),
.C(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_171),
.A2(n_174),
.B1(n_242),
.B2(n_246),
.Y(n_241)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_174),
.B(n_237),
.C(n_246),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_187),
.C(n_191),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_177),
.B(n_282),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.C(n_185),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_178),
.B(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_182),
.B(n_185),
.Y(n_265)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_187),
.B(n_191),
.Y(n_282)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_189),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_232),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_208),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_196),
.B(n_209),
.C(n_220),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_202),
.Y(n_207)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_206),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_220),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.C(n_216),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_210),
.B(n_216),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx24_ASAP7_75t_SL g532 ( 
.A(n_220),
.Y(n_532)
);

FAx1_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_227),
.CI(n_231),
.CON(n_220),
.SN(n_220)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_221),
.B(n_227),
.C(n_231),
.Y(n_506)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx8_ASAP7_75t_L g412 ( 
.A(n_225),
.Y(n_412)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_226),
.Y(n_393)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_230),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_247),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_234),
.B(n_236),
.C(n_247),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_238),
.B(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.C(n_251),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_251),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.C(n_260),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_255),
.B(n_258),
.Y(n_486)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_260),
.B(n_486),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_280),
.C(n_283),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_262),
.B(n_479),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.C(n_273),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_263),
.A2(n_264),
.B1(n_457),
.B2(n_458),
.Y(n_456)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_266),
.A2(n_267),
.B(n_269),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_266),
.B(n_273),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_268),
.Y(n_313)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_268),
.Y(n_331)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.C(n_278),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_434)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_278),
.B(n_434),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_279),
.B(n_370),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_280),
.A2(n_281),
.B1(n_283),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_283),
.Y(n_480)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_294),
.C(n_297),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_285),
.B(n_468),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.C(n_291),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_286),
.B(n_446),
.Y(n_445)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_289),
.A2(n_291),
.B1(n_292),
.B2(n_447),
.Y(n_446)
);

CKINVDCx14_ASAP7_75t_R g447 ( 
.A(n_289),
.Y(n_447)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_294),
.B(n_297),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_296),
.Y(n_370)
);

AOI21x1_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_484),
.B(n_489),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_471),
.B(n_483),
.Y(n_299)
);

AOI21x1_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_453),
.B(n_470),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_427),
.B(n_452),
.Y(n_301)
);

AOI21x1_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_397),
.B(n_426),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_362),
.B(n_396),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_342),
.B(n_361),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_319),
.B(n_341),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_316),
.B(n_318),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_314),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_314),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_317),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_311),
.Y(n_320)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_320),
.B(n_321),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_332),
.B2(n_333),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_322),
.B(n_335),
.C(n_337),
.Y(n_360)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_329),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_324),
.B(n_329),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_337),
.B2(n_338),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_360),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_360),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_352),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_351),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_351),
.C(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_350),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_350),
.Y(n_367)
);

INVx6_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_352),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_380),
.C(n_381),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_359),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_355),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_359),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_365),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_363),
.B(n_365),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_378),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_366),
.B(n_379),
.C(n_382),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_367),
.B(n_369),
.C(n_371),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_371),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_374),
.B1(n_375),
.B2(n_377),
.Y(n_371)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_372),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_374),
.B(n_377),
.Y(n_407)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_SL g421 ( 
.A(n_376),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_382),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_387),
.Y(n_382)
);

MAJx2_ASAP7_75t_L g424 ( 
.A(n_383),
.B(n_391),
.C(n_394),
.Y(n_424)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_388),
.A2(n_391),
.B1(n_394),
.B2(n_395),
.Y(n_387)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_388),
.Y(n_394)
);

INVx5_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_390),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_391),
.Y(n_395)
);

INVx6_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_425),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_425),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_409),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_408),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_400),
.B(n_408),
.C(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_407),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_406),
.Y(n_401)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_402),
.Y(n_441)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_406),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_407),
.B(n_441),
.C(n_442),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_409),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_416),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_410),
.B(n_418),
.C(n_423),
.Y(n_430)
);

BUFx24_ASAP7_75t_SL g533 ( 
.A(n_410),
.Y(n_533)
);

FAx1_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_413),
.CI(n_414),
.CON(n_410),
.SN(n_410)
);

MAJx2_ASAP7_75t_L g438 ( 
.A(n_411),
.B(n_413),
.C(n_414),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_418),
.B1(n_423),
.B2(n_424),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_422),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_419),
.B(n_422),
.Y(n_437)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_424),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_428),
.B(n_450),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_450),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_439),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_431),
.C(n_439),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_432),
.A2(n_433),
.B1(n_435),
.B2(n_436),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_432),
.B(n_462),
.C(n_463),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_438),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_443),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_440),
.B(n_444),
.C(n_449),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_445),
.B1(n_448),
.B2(n_449),
.Y(n_443)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_444),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_445),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_454),
.B(n_469),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_469),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_455),
.B(n_460),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_459),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_456),
.B(n_459),
.C(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_457),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_460),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_461),
.B(n_464),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_461),
.B(n_465),
.C(n_467),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_467),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_481),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_481),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_473),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_478),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_475),
.B(n_478),
.C(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_485),
.B(n_487),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_485),
.B(n_487),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_519),
.Y(n_491)
);

OAI21xp33_ASAP7_75t_L g523 ( 
.A1(n_492),
.A2(n_524),
.B(n_525),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_493),
.B(n_512),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_493),
.B(n_512),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_494),
.A2(n_495),
.B1(n_501),
.B2(n_511),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_494),
.B(n_502),
.C(n_507),
.Y(n_530)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_497),
.C(n_499),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_514),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_497),
.A2(n_499),
.B1(n_500),
.B2(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_497),
.Y(n_515)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_501),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_507),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_505),
.C(n_506),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_503),
.B(n_517),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_505),
.B(n_506),
.Y(n_517)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_508),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_516),
.C(n_518),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_516),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_518),
.B(n_521),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_520),
.B(n_522),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_522),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_530),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_527),
.B(n_530),
.Y(n_531)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_528),
.Y(n_529)
);


endmodule