module real_aes_118_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_404;
wire n_147;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_0), .B(n_494), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_1), .A2(n_496), .B(n_497), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_2), .B(n_813), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_3), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g782 ( .A1(n_3), .A2(n_783), .B(n_787), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_4), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_5), .B(n_205), .Y(n_531) );
INVx1_ASAP7_75t_L g137 ( .A(n_6), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_7), .B(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_8), .B(n_205), .Y(n_580) );
INVx1_ASAP7_75t_L g175 ( .A(n_9), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g813 ( .A(n_10), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_11), .Y(n_143) );
NAND2xp33_ASAP7_75t_L g572 ( .A(n_12), .B(n_202), .Y(n_572) );
INVx2_ASAP7_75t_L g119 ( .A(n_13), .Y(n_119) );
AOI221x1_ASAP7_75t_L g516 ( .A1(n_14), .A2(n_26), .B1(n_494), .B2(n_496), .C(n_517), .Y(n_516) );
CKINVDCx16_ASAP7_75t_R g477 ( .A(n_15), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_16), .B(n_494), .Y(n_568) );
INVx1_ASAP7_75t_L g203 ( .A(n_17), .Y(n_203) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_18), .A2(n_172), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_19), .B(n_167), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_20), .B(n_205), .Y(n_505) );
AO21x1_ASAP7_75t_L g526 ( .A1(n_21), .A2(n_494), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g481 ( .A(n_22), .Y(n_481) );
INVx1_ASAP7_75t_L g200 ( .A(n_23), .Y(n_200) );
INVx1_ASAP7_75t_SL g187 ( .A(n_24), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_25), .B(n_130), .Y(n_245) );
AOI33xp33_ASAP7_75t_L g225 ( .A1(n_27), .A2(n_53), .A3(n_123), .B1(n_148), .B2(n_226), .B3(n_227), .Y(n_225) );
NAND2x1_ASAP7_75t_L g547 ( .A(n_28), .B(n_205), .Y(n_547) );
NAND2x1_ASAP7_75t_L g579 ( .A(n_29), .B(n_202), .Y(n_579) );
INVx1_ASAP7_75t_L g128 ( .A(n_30), .Y(n_128) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_31), .A2(n_86), .B(n_119), .Y(n_118) );
OR2x2_ASAP7_75t_L g169 ( .A(n_31), .B(n_86), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_32), .B(n_152), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_33), .B(n_202), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_34), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_35), .B(n_205), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_36), .B(n_202), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_37), .A2(n_496), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g136 ( .A(n_38), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g147 ( .A(n_38), .Y(n_147) );
AND2x2_ASAP7_75t_L g156 ( .A(n_38), .B(n_126), .Y(n_156) );
OR2x6_ASAP7_75t_L g479 ( .A(n_39), .B(n_480), .Y(n_479) );
NOR3xp33_ASAP7_75t_L g811 ( .A(n_39), .B(n_477), .C(n_812), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_40), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_41), .B(n_494), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_42), .B(n_152), .Y(n_160) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_43), .A2(n_117), .B1(n_194), .B2(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_44), .B(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_45), .B(n_130), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_46), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_47), .B(n_202), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_48), .B(n_172), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_49), .B(n_130), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_50), .A2(n_496), .B(n_578), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_51), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_52), .B(n_202), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_54), .B(n_130), .Y(n_164) );
INVx1_ASAP7_75t_L g124 ( .A(n_55), .Y(n_124) );
INVx1_ASAP7_75t_L g132 ( .A(n_55), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_56), .Y(n_794) );
AND2x2_ASAP7_75t_L g166 ( .A(n_57), .B(n_167), .Y(n_166) );
AOI221xp5_ASAP7_75t_L g173 ( .A1(n_58), .A2(n_74), .B1(n_145), .B2(n_152), .C(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_59), .B(n_152), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_60), .B(n_205), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_61), .B(n_117), .Y(n_150) );
AOI21xp5_ASAP7_75t_SL g212 ( .A1(n_62), .A2(n_145), .B(n_213), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_63), .A2(n_496), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g197 ( .A(n_64), .Y(n_197) );
AO21x1_ASAP7_75t_L g528 ( .A1(n_65), .A2(n_496), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_66), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g163 ( .A(n_67), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_68), .B(n_494), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_69), .A2(n_145), .B(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g541 ( .A(n_70), .B(n_168), .Y(n_541) );
INVx1_ASAP7_75t_L g126 ( .A(n_71), .Y(n_126) );
INVx1_ASAP7_75t_L g134 ( .A(n_71), .Y(n_134) );
AND2x2_ASAP7_75t_L g582 ( .A(n_72), .B(n_116), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_73), .B(n_152), .Y(n_228) );
AND2x2_ASAP7_75t_L g189 ( .A(n_75), .B(n_116), .Y(n_189) );
INVx1_ASAP7_75t_L g198 ( .A(n_76), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_77), .A2(n_145), .B(n_186), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_78), .A2(n_145), .B(n_220), .C(n_244), .Y(n_243) );
OAI22xp33_ASAP7_75t_SL g802 ( .A1(n_79), .A2(n_483), .B1(n_785), .B2(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_79), .Y(n_803) );
INVx1_ASAP7_75t_L g482 ( .A(n_80), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_80), .B(n_481), .Y(n_810) );
AND2x2_ASAP7_75t_L g491 ( .A(n_81), .B(n_116), .Y(n_491) );
AND2x2_ASAP7_75t_SL g210 ( .A(n_82), .B(n_116), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_83), .B(n_494), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_84), .A2(n_145), .B1(n_223), .B2(n_224), .Y(n_222) );
AND2x2_ASAP7_75t_L g527 ( .A(n_85), .B(n_194), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_87), .B(n_202), .Y(n_506) );
AND2x2_ASAP7_75t_L g550 ( .A(n_88), .B(n_116), .Y(n_550) );
INVx1_ASAP7_75t_L g214 ( .A(n_89), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_90), .B(n_205), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_91), .A2(n_496), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_92), .B(n_202), .Y(n_518) );
AND2x2_ASAP7_75t_L g229 ( .A(n_93), .B(n_116), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_94), .B(n_205), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g120 ( .A1(n_95), .A2(n_121), .B(n_127), .C(n_135), .Y(n_120) );
BUFx2_ASAP7_75t_L g799 ( .A(n_96), .Y(n_799) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_97), .A2(n_496), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_98), .B(n_130), .Y(n_215) );
AOI21xp33_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_807), .B(n_814), .Y(n_99) );
AO21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_797), .B(n_800), .Y(n_100) );
OAI211xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_104), .B(n_782), .C(n_792), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
OAI22x1_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_474), .B1(n_483), .B2(n_778), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
OAI22xp5_ASAP7_75t_SL g783 ( .A1(n_107), .A2(n_784), .B1(n_785), .B2(n_786), .Y(n_783) );
NAND3x1_ASAP7_75t_L g107 ( .A(n_108), .B(n_353), .C(n_420), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_313), .Y(n_108) );
NOR3x1_ASAP7_75t_L g109 ( .A(n_110), .B(n_264), .C(n_293), .Y(n_109) );
OAI221xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_178), .B1(n_217), .B2(n_232), .C(n_249), .Y(n_110) );
A2O1A1Ixp33_ASAP7_75t_SL g427 ( .A1(n_111), .A2(n_191), .B(n_428), .C(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_112), .A2(n_399), .B1(n_402), .B2(n_404), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_112), .B(n_218), .Y(n_473) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_157), .Y(n_112) );
BUFx2_ASAP7_75t_L g392 ( .A(n_113), .Y(n_392) );
INVx1_ASAP7_75t_SL g405 ( .A(n_113), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_113), .B(n_260), .Y(n_447) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g230 ( .A(n_114), .B(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g275 ( .A(n_114), .B(n_171), .Y(n_275) );
INVx1_ASAP7_75t_L g286 ( .A(n_114), .Y(n_286) );
INVx2_ASAP7_75t_L g290 ( .A(n_114), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_114), .B(n_261), .Y(n_417) );
OR2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_140), .Y(n_114) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_120), .B1(n_138), .B2(n_139), .Y(n_115) );
INVx3_ASAP7_75t_L g139 ( .A(n_116), .Y(n_139) );
INVx4_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_117), .B(n_142), .Y(n_141) );
INVx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx4f_ASAP7_75t_L g172 ( .A(n_118), .Y(n_172) );
AND2x2_ASAP7_75t_SL g168 ( .A(n_119), .B(n_169), .Y(n_168) );
AND2x4_ASAP7_75t_L g194 ( .A(n_119), .B(n_169), .Y(n_194) );
INVxp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
O2A1O1Ixp33_ASAP7_75t_L g162 ( .A1(n_122), .A2(n_163), .B(n_164), .C(n_165), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_SL g174 ( .A1(n_122), .A2(n_165), .B(n_175), .C(n_176), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_SL g186 ( .A1(n_122), .A2(n_165), .B(n_187), .C(n_188), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_122), .A2(n_129), .B1(n_197), .B2(n_198), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_122), .A2(n_165), .B(n_214), .C(n_215), .Y(n_213) );
INVx2_ASAP7_75t_L g247 ( .A(n_122), .Y(n_247) );
OR2x6_ASAP7_75t_L g122 ( .A(n_123), .B(n_125), .Y(n_122) );
AND2x2_ASAP7_75t_L g153 ( .A(n_123), .B(n_154), .Y(n_153) );
INVxp33_ASAP7_75t_L g226 ( .A(n_123), .Y(n_226) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g149 ( .A(n_124), .B(n_137), .Y(n_149) );
AND2x4_ASAP7_75t_L g205 ( .A(n_124), .B(n_133), .Y(n_205) );
INVx3_ASAP7_75t_L g148 ( .A(n_125), .Y(n_148) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x6_ASAP7_75t_L g202 ( .A(n_126), .B(n_131), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g494 ( .A(n_130), .B(n_136), .Y(n_494) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx5_ASAP7_75t_L g165 ( .A(n_136), .Y(n_165) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_137), .Y(n_154) );
AO21x2_ASAP7_75t_L g158 ( .A1(n_139), .A2(n_159), .B(n_166), .Y(n_158) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_139), .A2(n_159), .B(n_166), .Y(n_261) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_139), .A2(n_535), .B(n_541), .Y(n_534) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_139), .A2(n_544), .B(n_550), .Y(n_543) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_139), .A2(n_544), .B(n_550), .Y(n_556) );
AO21x2_ASAP7_75t_L g559 ( .A1(n_139), .A2(n_535), .B(n_541), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_144), .B1(n_150), .B2(n_151), .Y(n_140) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVxp67_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_149), .Y(n_145) );
NOR2x1p5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
INVx1_ASAP7_75t_L g227 ( .A(n_148), .Y(n_227) );
AND2x6_ASAP7_75t_L g496 ( .A(n_149), .B(n_156), .Y(n_496) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
INVx1_ASAP7_75t_L g240 ( .A(n_153), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_155), .Y(n_241) );
BUFx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g366 ( .A(n_157), .B(n_367), .Y(n_366) );
NOR2x1_ASAP7_75t_L g157 ( .A(n_158), .B(n_170), .Y(n_157) );
INVx2_ASAP7_75t_L g269 ( .A(n_158), .Y(n_269) );
AND2x2_ASAP7_75t_L g289 ( .A(n_158), .B(n_290), .Y(n_289) );
NOR2xp67_ASAP7_75t_L g414 ( .A(n_158), .B(n_290), .Y(n_414) );
AND2x2_ASAP7_75t_L g439 ( .A(n_158), .B(n_282), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_165), .B(n_194), .Y(n_206) );
INVx1_ASAP7_75t_L g223 ( .A(n_165), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_165), .A2(n_245), .B(n_246), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_165), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_165), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_165), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_165), .A2(n_530), .B(n_531), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_165), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_165), .A2(n_547), .B(n_548), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_165), .A2(n_571), .B(n_572), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_165), .A2(n_579), .B(n_580), .Y(n_578) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_167), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_167), .A2(n_493), .B(n_495), .Y(n_492) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_167), .A2(n_516), .B(n_520), .Y(n_515) );
OA21x2_ASAP7_75t_L g586 ( .A1(n_167), .A2(n_516), .B(n_520), .Y(n_586) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g231 ( .A(n_171), .Y(n_231) );
INVx1_ASAP7_75t_L g253 ( .A(n_171), .Y(n_253) );
INVxp67_ASAP7_75t_L g292 ( .A(n_171), .Y(n_292) );
AND2x4_ASAP7_75t_L g332 ( .A(n_171), .B(n_333), .Y(n_332) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_171), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_171), .B(n_283), .Y(n_418) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_177), .Y(n_171) );
INVx2_ASAP7_75t_SL g220 ( .A(n_172), .Y(n_220) );
INVx1_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_190), .Y(n_179) );
AND2x2_ASAP7_75t_L g306 ( .A(n_180), .B(n_278), .Y(n_306) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_181), .Y(n_234) );
AND2x2_ASAP7_75t_L g262 ( .A(n_181), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g273 ( .A(n_181), .Y(n_273) );
INVx1_ASAP7_75t_L g297 ( .A(n_181), .Y(n_297) );
AND2x2_ASAP7_75t_L g300 ( .A(n_181), .B(n_192), .Y(n_300) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_181), .Y(n_322) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_189), .Y(n_181) );
AO21x2_ASAP7_75t_L g575 ( .A1(n_182), .A2(n_576), .B(n_582), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
NOR2x1_ASAP7_75t_L g190 ( .A(n_191), .B(n_207), .Y(n_190) );
AND2x2_ASAP7_75t_L g287 ( .A(n_191), .B(n_209), .Y(n_287) );
NAND2x1_ASAP7_75t_L g320 ( .A(n_191), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g423 ( .A(n_191), .Y(n_423) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx3_ASAP7_75t_L g263 ( .A(n_192), .Y(n_263) );
AND2x2_ASAP7_75t_L g278 ( .A(n_192), .B(n_237), .Y(n_278) );
NOR2x1_ASAP7_75t_SL g347 ( .A(n_192), .B(n_209), .Y(n_347) );
AND2x4_ASAP7_75t_L g192 ( .A(n_193), .B(n_195), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_194), .A2(n_212), .B(n_216), .Y(n_211) );
INVx1_ASAP7_75t_SL g501 ( .A(n_194), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_194), .B(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_194), .A2(n_568), .B(n_569), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_199), .B(n_206), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B1(n_203), .B2(n_204), .Y(n_199) );
INVxp67_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVxp67_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2x1_ASAP7_75t_L g384 ( .A(n_207), .B(n_371), .Y(n_384) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g309 ( .A(n_208), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx4_ASAP7_75t_L g248 ( .A(n_209), .Y(n_248) );
AND2x4_ASAP7_75t_L g255 ( .A(n_209), .B(n_256), .Y(n_255) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_209), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_209), .B(n_272), .Y(n_372) );
AND2x2_ASAP7_75t_L g400 ( .A(n_209), .B(n_237), .Y(n_400) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
NAND2x1_ASAP7_75t_SL g217 ( .A(n_218), .B(n_230), .Y(n_217) );
OR2x2_ASAP7_75t_L g428 ( .A(n_218), .B(n_340), .Y(n_428) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x4_ASAP7_75t_L g268 ( .A(n_219), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g333 ( .A(n_219), .Y(n_333) );
AND2x2_ASAP7_75t_L g367 ( .A(n_219), .B(n_290), .Y(n_367) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_229), .Y(n_219) );
AO21x2_ASAP7_75t_L g283 ( .A1(n_220), .A2(n_221), .B(n_229), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_222), .B(n_228), .Y(n_221) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx3_ASAP7_75t_L g340 ( .A(n_230), .Y(n_340) );
AND2x2_ASAP7_75t_L g348 ( .A(n_230), .B(n_281), .Y(n_348) );
AND2x2_ASAP7_75t_L g465 ( .A(n_230), .B(n_268), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
BUFx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g419 ( .A(n_234), .B(n_360), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_234), .B(n_259), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_235), .A2(n_296), .B(n_299), .Y(n_295) );
AND2x2_ASAP7_75t_L g365 ( .A(n_235), .B(n_271), .Y(n_365) );
INVx2_ASAP7_75t_SL g452 ( .A(n_235), .Y(n_452) );
AND2x4_ASAP7_75t_SL g235 ( .A(n_236), .B(n_248), .Y(n_235) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g256 ( .A(n_237), .Y(n_256) );
INVx2_ASAP7_75t_L g303 ( .A(n_237), .Y(n_303) );
AND2x4_ASAP7_75t_L g310 ( .A(n_237), .B(n_263), .Y(n_310) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_243), .Y(n_237) );
NOR3xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .C(n_242), .Y(n_239) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_248), .Y(n_266) );
AND2x4_ASAP7_75t_L g342 ( .A(n_248), .B(n_256), .Y(n_342) );
OR2x2_ASAP7_75t_L g468 ( .A(n_248), .B(n_469), .Y(n_468) );
NAND4xp25_ASAP7_75t_L g249 ( .A(n_250), .B(n_254), .C(n_257), .D(n_262), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g315 ( .A(n_251), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g412 ( .A(n_251), .Y(n_412) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2x1p5_ASAP7_75t_L g312 ( .A(n_252), .B(n_260), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_252), .B(n_317), .Y(n_446) );
BUFx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_255), .B(n_271), .Y(n_324) );
INVx2_ASAP7_75t_L g426 ( .A(n_255), .Y(n_426) );
AND2x2_ASAP7_75t_SL g436 ( .A(n_255), .B(n_296), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_255), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g328 ( .A(n_259), .B(n_275), .Y(n_328) );
AND2x2_ASAP7_75t_L g396 ( .A(n_259), .B(n_332), .Y(n_396) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x4_ASAP7_75t_L g281 ( .A(n_260), .B(n_282), .Y(n_281) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_261), .Y(n_335) );
AND2x2_ASAP7_75t_L g386 ( .A(n_261), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_261), .B(n_283), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_262), .B(n_426), .Y(n_433) );
INVx1_ASAP7_75t_SL g469 ( .A(n_262), .Y(n_469) );
INVx1_ASAP7_75t_L g298 ( .A(n_263), .Y(n_298) );
AND2x2_ASAP7_75t_L g360 ( .A(n_263), .B(n_303), .Y(n_360) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_274), .B(n_276), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
AND2x2_ASAP7_75t_L g326 ( .A(n_268), .B(n_275), .Y(n_326) );
AND2x2_ASAP7_75t_L g434 ( .A(n_268), .B(n_285), .Y(n_434) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g308 ( .A(n_271), .Y(n_308) );
AND2x2_ASAP7_75t_L g341 ( .A(n_271), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g346 ( .A(n_271), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_271), .B(n_310), .Y(n_395) );
NOR3xp33_ASAP7_75t_L g445 ( .A(n_271), .B(n_446), .C(n_447), .Y(n_445) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVxp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_280), .B1(n_287), .B2(n_288), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx2_ASAP7_75t_L g371 ( .A(n_278), .Y(n_371) );
AND2x2_ASAP7_75t_L g305 ( .A(n_279), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g327 ( .A(n_279), .B(n_300), .Y(n_327) );
AND2x2_ASAP7_75t_SL g359 ( .A(n_279), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_284), .Y(n_280) );
INVx1_ASAP7_75t_L g338 ( .A(n_281), .Y(n_338) );
AND2x2_ASAP7_75t_L g291 ( .A(n_282), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g317 ( .A(n_282), .Y(n_317) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g380 ( .A(n_286), .B(n_332), .Y(n_380) );
INVx1_ASAP7_75t_L g438 ( .A(n_286), .Y(n_438) );
INVx1_ASAP7_75t_L g294 ( .A(n_288), .Y(n_294) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_289), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g425 ( .A(n_289), .B(n_332), .Y(n_425) );
AND2x2_ASAP7_75t_L g391 ( .A(n_291), .B(n_392), .Y(n_391) );
NAND2x1p5_ASAP7_75t_L g459 ( .A(n_291), .B(n_460), .Y(n_459) );
OAI21xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_295), .B(n_304), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_296), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g352 ( .A(n_296), .B(n_301), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_296), .B(n_342), .Y(n_403) );
AND2x4_ASAP7_75t_SL g296 ( .A(n_297), .B(n_298), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_297), .B(n_360), .Y(n_390) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_297), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_299), .A2(n_326), .B1(n_327), .B2(n_328), .Y(n_325) );
AND2x2_ASAP7_75t_SL g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_300), .B(n_342), .Y(n_361) );
INVx1_ASAP7_75t_L g462 ( .A(n_300), .Y(n_462) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI21xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_307), .B(n_311), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_306), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g443 ( .A(n_309), .Y(n_443) );
INVx4_ASAP7_75t_L g345 ( .A(n_310), .Y(n_345) );
INVxp33_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g373 ( .A(n_312), .B(n_374), .Y(n_373) );
NOR2x1_ASAP7_75t_L g313 ( .A(n_314), .B(n_329), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_318), .B(n_325), .Y(n_314) );
INVx1_ASAP7_75t_L g363 ( .A(n_316), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_323), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g368 ( .A(n_320), .Y(n_368) );
INVx1_ASAP7_75t_L g401 ( .A(n_321), .Y(n_401) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_326), .A2(n_365), .B1(n_366), .B2(n_368), .Y(n_364) );
INVx1_ASAP7_75t_L g378 ( .A(n_327), .Y(n_378) );
NAND4xp25_ASAP7_75t_SL g329 ( .A(n_330), .B(n_336), .C(n_343), .D(n_349), .Y(n_329) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
INVx1_ASAP7_75t_L g351 ( .A(n_332), .Y(n_351) );
AND2x2_ASAP7_75t_L g463 ( .A(n_332), .B(n_460), .Y(n_463) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_341), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g470 ( .A(n_340), .B(n_407), .Y(n_470) );
INVx1_ASAP7_75t_L g467 ( .A(n_341), .Y(n_467) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_342), .Y(n_376) );
OAI21xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_346), .B(n_348), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_381), .Y(n_353) );
NOR3xp33_ASAP7_75t_L g354 ( .A(n_355), .B(n_369), .C(n_377), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_362), .B(n_364), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_361), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_359), .A2(n_391), .B1(n_394), .B2(n_396), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g369 ( .A1(n_362), .A2(n_370), .B1(n_373), .B2(n_375), .Y(n_369) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g374 ( .A(n_367), .Y(n_374) );
AND2x4_ASAP7_75t_L g385 ( .A(n_367), .B(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_372), .Y(n_472) );
AOI31xp33_ASAP7_75t_L g471 ( .A1(n_375), .A2(n_448), .A3(n_472), .B(n_473), .Y(n_471) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_382), .B(n_397), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_383), .B(n_393), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_388), .B2(n_391), .Y(n_383) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_387), .Y(n_451) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_395), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_398), .B(n_408), .Y(n_397) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
AND2x2_ASAP7_75t_L g409 ( .A(n_400), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g448 ( .A(n_400), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g457 ( .A1(n_400), .A2(n_458), .B1(n_461), .B2(n_463), .Y(n_457) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_405), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_411), .B1(n_415), .B2(n_419), .Y(n_408) );
NOR2xp33_ASAP7_75t_SL g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx2_ASAP7_75t_SL g460 ( .A(n_417), .Y(n_460) );
INVx2_ASAP7_75t_L g441 ( .A(n_418), .Y(n_441) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_455), .Y(n_420) );
AOI211xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_427), .B(n_430), .C(n_444), .Y(n_421) );
OAI21xp33_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B(n_426), .Y(n_422) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g429 ( .A(n_426), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_431), .B(n_435), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_437), .B1(n_440), .B2(n_442), .Y(n_435) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
AND2x2_ASAP7_75t_L g440 ( .A(n_438), .B(n_441), .Y(n_440) );
AO22x1_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_448), .B1(n_449), .B2(n_453), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_466), .C(n_471), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_457), .B(n_464), .Y(n_456) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AOI21xp33_ASAP7_75t_R g466 ( .A1(n_467), .A2(n_468), .B(n_470), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_475), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_475), .Y(n_784) );
CKINVDCx11_ASAP7_75t_R g475 ( .A(n_476), .Y(n_475) );
OR2x6_ASAP7_75t_SL g476 ( .A(n_477), .B(n_478), .Y(n_476) );
AND2x6_ASAP7_75t_SL g781 ( .A(n_477), .B(n_479), .Y(n_781) );
OR2x2_ASAP7_75t_L g791 ( .A(n_477), .B(n_479), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_477), .B(n_478), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
BUFx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx3_ASAP7_75t_SL g785 ( .A(n_484), .Y(n_785) );
NOR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_665), .Y(n_484) );
AO211x2_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_510), .B(n_560), .C(n_633), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVxp67_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
AND3x2_ASAP7_75t_L g714 ( .A(n_488), .B(n_595), .C(n_611), .Y(n_714) );
AND2x4_ASAP7_75t_L g717 ( .A(n_488), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_500), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g573 ( .A(n_489), .B(n_574), .Y(n_573) );
INVx4_ASAP7_75t_L g626 ( .A(n_489), .Y(n_626) );
AND2x2_ASAP7_75t_SL g711 ( .A(n_489), .B(n_620), .Y(n_711) );
AND2x2_ASAP7_75t_L g754 ( .A(n_489), .B(n_575), .Y(n_754) );
INVx5_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx2_ASAP7_75t_L g603 ( .A(n_490), .Y(n_603) );
AND2x2_ASAP7_75t_L g622 ( .A(n_490), .B(n_566), .Y(n_622) );
AND2x2_ASAP7_75t_L g640 ( .A(n_490), .B(n_575), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_490), .B(n_574), .Y(n_700) );
NOR2x1_ASAP7_75t_SL g727 ( .A(n_490), .B(n_500), .Y(n_727) );
OR2x6_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_500), .B(n_566), .Y(n_565) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B(n_508), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_501), .B(n_509), .Y(n_508) );
AO21x2_ASAP7_75t_L g599 ( .A1(n_501), .A2(n_502), .B(n_508), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_507), .Y(n_502) );
AO21x1_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_542), .B(n_551), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OAI22xp33_ASAP7_75t_L g608 ( .A1(n_512), .A2(n_609), .B1(n_613), .B2(n_614), .Y(n_608) );
OR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_521), .Y(n_512) );
AND2x2_ASAP7_75t_L g669 ( .A(n_513), .B(n_557), .Y(n_669) );
BUFx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x4_ASAP7_75t_L g602 ( .A(n_514), .B(n_585), .Y(n_602) );
AND2x2_ASAP7_75t_L g674 ( .A(n_514), .B(n_559), .Y(n_674) );
AND2x2_ASAP7_75t_L g693 ( .A(n_514), .B(n_659), .Y(n_693) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g552 ( .A(n_515), .Y(n_552) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_515), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_521), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g653 ( .A(n_522), .B(n_554), .Y(n_653) );
AND2x4_ASAP7_75t_L g522 ( .A(n_523), .B(n_534), .Y(n_522) );
AND2x2_ASAP7_75t_L g557 ( .A(n_523), .B(n_558), .Y(n_557) );
OR2x2_ASAP7_75t_L g590 ( .A(n_523), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_SL g650 ( .A(n_523), .B(n_586), .Y(n_650) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx2_ASAP7_75t_L g743 ( .A(n_524), .Y(n_743) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g585 ( .A(n_525), .Y(n_585) );
OAI21x1_ASAP7_75t_SL g525 ( .A1(n_526), .A2(n_528), .B(n_532), .Y(n_525) );
INVx1_ASAP7_75t_L g533 ( .A(n_527), .Y(n_533) );
INVx2_ASAP7_75t_L g591 ( .A(n_534), .Y(n_591) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_534), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_536), .B(n_540), .Y(n_535) );
INVx2_ASAP7_75t_L g587 ( .A(n_542), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_542), .B(n_719), .Y(n_745) );
AND2x2_ASAP7_75t_L g764 ( .A(n_542), .B(n_754), .Y(n_764) );
BUFx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x4_ASAP7_75t_SL g632 ( .A(n_543), .B(n_591), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_549), .Y(n_544) );
AND2x2_ASAP7_75t_SL g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AND2x2_ASAP7_75t_L g631 ( .A(n_552), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_552), .B(n_601), .Y(n_636) );
INVx1_ASAP7_75t_SL g763 ( .A(n_552), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_553), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
INVx1_ASAP7_75t_L g589 ( .A(n_554), .Y(n_589) );
AND2x2_ASAP7_75t_L g775 ( .A(n_554), .B(n_776), .Y(n_775) );
BUFx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g651 ( .A(n_555), .B(n_558), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_555), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g705 ( .A(n_555), .B(n_559), .Y(n_705) );
AND2x2_ASAP7_75t_L g736 ( .A(n_555), .B(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g601 ( .A(n_556), .B(n_559), .Y(n_601) );
INVxp67_ASAP7_75t_L g618 ( .A(n_556), .Y(n_618) );
BUFx3_ASAP7_75t_L g659 ( .A(n_556), .Y(n_659) );
AND2x2_ASAP7_75t_L g679 ( .A(n_557), .B(n_680), .Y(n_679) );
NAND2xp33_ASAP7_75t_L g692 ( .A(n_557), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_558), .B(n_585), .Y(n_648) );
AND2x2_ASAP7_75t_L g737 ( .A(n_558), .B(n_586), .Y(n_737) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g664 ( .A(n_559), .B(n_586), .Y(n_664) );
OR3x1_ASAP7_75t_L g560 ( .A(n_561), .B(n_608), .C(n_623), .Y(n_560) );
OAI321xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_573), .A3(n_583), .B1(n_588), .B2(n_592), .C(n_600), .Y(n_561) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_565), .Y(n_639) );
INVxp67_ASAP7_75t_SL g657 ( .A(n_565), .Y(n_657) );
OR2x2_ASAP7_75t_L g661 ( .A(n_565), .B(n_573), .Y(n_661) );
BUFx3_ASAP7_75t_L g595 ( .A(n_566), .Y(n_595) );
AND2x2_ASAP7_75t_L g612 ( .A(n_566), .B(n_598), .Y(n_612) );
INVx1_ASAP7_75t_L g629 ( .A(n_566), .Y(n_629) );
INVx2_ASAP7_75t_L g645 ( .A(n_566), .Y(n_645) );
OR2x2_ASAP7_75t_L g684 ( .A(n_566), .B(n_574), .Y(n_684) );
INVx2_ASAP7_75t_L g672 ( .A(n_573), .Y(n_672) );
AND2x2_ASAP7_75t_L g596 ( .A(n_574), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g611 ( .A(n_574), .Y(n_611) );
AND2x4_ASAP7_75t_L g620 ( .A(n_574), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_574), .B(n_597), .Y(n_643) );
AND2x2_ASAP7_75t_L g750 ( .A(n_574), .B(n_645), .Y(n_750) );
INVx4_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_575), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_581), .Y(n_576) );
INVx1_ASAP7_75t_L g637 ( .A(n_583), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_584), .B(n_587), .Y(n_583) );
AND2x2_ASAP7_75t_L g724 ( .A(n_584), .B(n_651), .Y(n_724) );
INVx1_ASAP7_75t_SL g741 ( .A(n_584), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_584), .B(n_717), .Y(n_770) );
AND2x4_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
OR2x2_ASAP7_75t_L g613 ( .A(n_585), .B(n_586), .Y(n_613) );
AND2x2_ASAP7_75t_L g706 ( .A(n_587), .B(n_602), .Y(n_706) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g729 ( .A(n_591), .B(n_602), .Y(n_729) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_593), .A2(n_742), .B1(n_747), .B2(n_749), .Y(n_746) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
AND2x2_ASAP7_75t_L g671 ( .A(n_594), .B(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g766 ( .A(n_594), .B(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g722 ( .A(n_595), .B(n_640), .Y(n_722) );
AND2x4_ASAP7_75t_L g676 ( .A(n_596), .B(n_622), .Y(n_676) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_598), .Y(n_774) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g607 ( .A(n_599), .Y(n_607) );
INVx1_ASAP7_75t_L g621 ( .A(n_599), .Y(n_621) );
NAND4xp25_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .C(n_603), .D(n_604), .Y(n_600) );
AND2x2_ASAP7_75t_L g758 ( .A(n_601), .B(n_743), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_601), .B(n_769), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_602), .B(n_678), .Y(n_677) );
OAI322xp33_ASAP7_75t_L g685 ( .A1(n_602), .A2(n_686), .A3(n_690), .B1(n_692), .B2(n_694), .C1(n_696), .C2(n_701), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_602), .B(n_651), .Y(n_701) );
INVx1_ASAP7_75t_L g769 ( .A(n_602), .Y(n_769) );
INVx2_ASAP7_75t_L g615 ( .A(n_603), .Y(n_615) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_606), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_607), .B(n_626), .Y(n_683) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_610), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g656 ( .A(n_611), .Y(n_656) );
AND2x2_ASAP7_75t_L g728 ( .A(n_611), .B(n_639), .Y(n_728) );
AOI31xp33_ASAP7_75t_L g614 ( .A1(n_612), .A2(n_615), .A3(n_616), .B(n_619), .Y(n_614) );
AND2x2_ASAP7_75t_L g625 ( .A(n_612), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g753 ( .A(n_612), .B(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_SL g760 ( .A(n_612), .B(n_640), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_612), .Y(n_761) );
INVx1_ASAP7_75t_SL g719 ( .A(n_613), .Y(n_719) );
NAND3xp33_ASAP7_75t_SL g747 ( .A(n_613), .B(n_741), .C(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g647 ( .A(n_618), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
AND2x2_ASAP7_75t_L g628 ( .A(n_620), .B(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g689 ( .A(n_620), .Y(n_689) );
AOI322xp5_ASAP7_75t_L g771 ( .A1(n_620), .A2(n_650), .A3(n_653), .B1(n_772), .B2(n_773), .C1(n_775), .C2(n_777), .Y(n_771) );
AND2x2_ASAP7_75t_L g777 ( .A(n_620), .B(n_626), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_627), .B(n_630), .Y(n_623) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_626), .B(n_645), .Y(n_644) );
AND2x4_ASAP7_75t_L g772 ( .A(n_626), .B(n_659), .Y(n_772) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g698 ( .A(n_629), .Y(n_698) );
AND2x2_ASAP7_75t_L g726 ( .A(n_629), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g773 ( .A(n_629), .B(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g678 ( .A(n_632), .Y(n_678) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
O2A1O1Ixp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_637), .B(n_638), .C(n_641), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
AND2x2_ASAP7_75t_L g695 ( .A(n_640), .B(n_645), .Y(n_695) );
OAI211xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_646), .B(n_652), .C(n_654), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g667 ( .A1(n_642), .A2(n_668), .B1(n_670), .B2(n_673), .C(n_675), .Y(n_667) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g687 ( .A(n_644), .Y(n_687) );
OR2x2_ASAP7_75t_L g707 ( .A(n_644), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
INVx1_ASAP7_75t_L g752 ( .A(n_647), .Y(n_752) );
INVx1_ASAP7_75t_L g776 ( .A(n_648), .Y(n_776) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_650), .B(n_651), .Y(n_649) );
AND2x2_ASAP7_75t_L g658 ( .A(n_650), .B(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_650), .B(n_720), .Y(n_732) );
INVx1_ASAP7_75t_L g712 ( .A(n_651), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_658), .B1(n_660), .B2(n_662), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx1_ASAP7_75t_SL g720 ( .A(n_659), .Y(n_720) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND4xp75_ASAP7_75t_L g665 ( .A(n_666), .B(n_702), .C(n_730), .D(n_755), .Y(n_665) );
NOR2xp67_ASAP7_75t_L g666 ( .A(n_667), .B(n_685), .Y(n_666) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_SL g742 ( .A(n_674), .B(n_743), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B1(n_679), .B2(n_681), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_678), .B(n_741), .Y(n_740) );
INVx2_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
OR2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx2_ASAP7_75t_L g718 ( .A(n_684), .Y(n_718) );
OR2x2_ASAP7_75t_L g733 ( .A(n_684), .B(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_687), .B(n_688), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g748 ( .A(n_693), .Y(n_748) );
INVx1_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
OAI21xp5_ASAP7_75t_SL g739 ( .A1(n_695), .A2(n_740), .B(n_742), .Y(n_739) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NOR2x1_ASAP7_75t_L g702 ( .A(n_703), .B(n_715), .Y(n_702) );
OAI221xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_707), .B1(n_710), .B2(n_712), .C(n_713), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
OAI21xp33_ASAP7_75t_L g751 ( .A1(n_705), .A2(n_752), .B(n_753), .Y(n_751) );
INVx3_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
OAI322xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_719), .A3(n_720), .B1(n_721), .B2(n_723), .C1(n_725), .C2(n_729), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
NOR2x1_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .Y(n_725) );
INVx1_ASAP7_75t_L g738 ( .A(n_726), .Y(n_738) );
INVx1_ASAP7_75t_L g734 ( .A(n_727), .Y(n_734) );
AND2x2_ASAP7_75t_L g749 ( .A(n_727), .B(n_750), .Y(n_749) );
NOR2x1_ASAP7_75t_L g730 ( .A(n_731), .B(n_744), .Y(n_730) );
OAI221xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B1(n_735), .B2(n_738), .C(n_739), .Y(n_731) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
OAI211xp5_ASAP7_75t_SL g744 ( .A1(n_738), .A2(n_745), .B(n_746), .C(n_751), .Y(n_744) );
INVx2_ASAP7_75t_SL g767 ( .A(n_754), .Y(n_767) );
NOR2x1_ASAP7_75t_L g755 ( .A(n_756), .B(n_765), .Y(n_755) );
OAI22xp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_759), .B1(n_761), .B2(n_762), .Y(n_756) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
OAI211xp5_ASAP7_75t_SL g765 ( .A1(n_766), .A2(n_768), .B(n_770), .C(n_771), .Y(n_765) );
CKINVDCx11_ASAP7_75t_R g778 ( .A(n_779), .Y(n_778) );
INVx3_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_781), .Y(n_780) );
CKINVDCx11_ASAP7_75t_R g786 ( .A(n_781), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_790), .Y(n_789) );
INVx3_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g800 ( .A1(n_792), .A2(n_801), .B(n_804), .Y(n_800) );
CKINVDCx14_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_795), .B(n_802), .Y(n_801) );
BUFx3_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_798), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_799), .Y(n_798) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_799), .Y(n_806) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx2_ASAP7_75t_L g816 ( .A(n_808), .Y(n_816) );
INVx3_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
AND2x2_ASAP7_75t_SL g809 ( .A(n_810), .B(n_811), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
endmodule