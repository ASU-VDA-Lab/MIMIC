module fake_aes_1429_n_18 (n_1, n_2, n_0, n_18);
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
BUFx2_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
NOR2xp33_ASAP7_75t_L g4 ( .A(n_0), .B(n_1), .Y(n_4) );
INVx3_ASAP7_75t_L g5 ( .A(n_1), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g6 ( .A(n_3), .B(n_0), .Y(n_6) );
OAI22xp5_ASAP7_75t_L g7 ( .A1(n_3), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_7) );
OAI22xp5_ASAP7_75t_L g8 ( .A1(n_4), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_8) );
AND2x4_ASAP7_75t_L g9 ( .A(n_6), .B(n_5), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_7), .B(n_5), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_9), .B(n_5), .Y(n_12) );
AOI221xp5_ASAP7_75t_L g13 ( .A1(n_11), .A2(n_10), .B1(n_8), .B2(n_9), .C(n_5), .Y(n_13) );
NAND4xp25_ASAP7_75t_SL g14 ( .A(n_12), .B(n_0), .C(n_2), .D(n_11), .Y(n_14) );
NOR4xp75_ASAP7_75t_SL g15 ( .A(n_14), .B(n_2), .C(n_0), .D(n_12), .Y(n_15) );
NOR2xp33_ASAP7_75t_R g16 ( .A(n_13), .B(n_11), .Y(n_16) );
OAI22xp5_ASAP7_75t_L g17 ( .A1(n_15), .A2(n_2), .B1(n_12), .B2(n_16), .Y(n_17) );
OAI21xp33_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_12), .B(n_15), .Y(n_18) );
endmodule