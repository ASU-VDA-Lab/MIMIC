module fake_jpeg_2272_n_535 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_535);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_535;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_293;
wire n_38;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_46),
.B(n_54),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_51),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_52),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_53),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_7),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

AND2x4_ASAP7_75t_SL g56 ( 
.A(n_29),
.B(n_16),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_56),
.B(n_61),
.Y(n_110)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_58),
.Y(n_134)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_7),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_78),
.Y(n_120)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_7),
.B(n_13),
.Y(n_71)
);

OR2x2_ASAP7_75t_SL g130 ( 
.A(n_71),
.B(n_24),
.Y(n_130)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_25),
.B(n_14),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_98),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_34),
.B(n_36),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_17),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_81),
.Y(n_131)
);

BUFx16f_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

INVx5_ASAP7_75t_SL g84 ( 
.A(n_17),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_84),
.B(n_24),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_36),
.B(n_14),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_88),
.Y(n_121)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_41),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_94),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_41),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_82),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_102),
.B(n_158),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_25),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_103),
.B(n_104),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_58),
.B(n_37),
.Y(n_104)
);

BUFx2_ASAP7_75t_SL g111 ( 
.A(n_82),
.Y(n_111)
);

CKINVDCx6p67_ASAP7_75t_R g208 ( 
.A(n_111),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_45),
.B1(n_42),
.B2(n_32),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_114),
.A2(n_22),
.B1(n_32),
.B2(n_45),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_60),
.B(n_37),
.C(n_43),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_115),
.B(n_13),
.Y(n_178)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_42),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_119),
.B(n_130),
.Y(n_187)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_122),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_80),
.B(n_42),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_132),
.B(n_140),
.Y(n_206)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_135),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_42),
.Y(n_140)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_147),
.Y(n_204)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_52),
.Y(n_157)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_56),
.A2(n_24),
.B(n_28),
.Y(n_158)
);

NAND2x1_ASAP7_75t_SL g176 ( 
.A(n_160),
.B(n_26),
.Y(n_176)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_161),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_162),
.Y(n_214)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_110),
.A2(n_56),
.B1(n_97),
.B2(n_89),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_164),
.A2(n_193),
.B1(n_194),
.B2(n_196),
.Y(n_229)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_121),
.B(n_72),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_168),
.B(n_173),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_110),
.A2(n_19),
.B1(n_131),
.B2(n_73),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_99),
.A2(n_49),
.B1(n_91),
.B2(n_48),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_170),
.A2(n_200),
.B1(n_32),
.B2(n_118),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_171),
.Y(n_238)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_172),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_69),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_108),
.A2(n_84),
.B(n_66),
.C(n_24),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_174),
.B(n_188),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_108),
.B(n_59),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_175),
.B(n_178),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_177),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_70),
.B(n_85),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_120),
.B(n_55),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_101),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_95),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_181),
.Y(n_232)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_145),
.A2(n_19),
.B1(n_45),
.B2(n_32),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_184),
.A2(n_190),
.B1(n_207),
.B2(n_209),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_128),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

CKINVDCx12_ASAP7_75t_R g190 ( 
.A(n_134),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_134),
.Y(n_191)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_120),
.B(n_95),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_133),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_126),
.B(n_52),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_127),
.B(n_22),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_201),
.Y(n_230)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_113),
.Y(n_198)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_129),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_125),
.Y(n_203)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_146),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_166),
.A2(n_67),
.B1(n_51),
.B2(n_53),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_217),
.B(n_245),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_136),
.B1(n_150),
.B2(n_148),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_221),
.A2(n_236),
.B1(n_237),
.B2(n_244),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_153),
.C(n_156),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_228),
.C(n_240),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_154),
.C(n_152),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_112),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_177),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_192),
.A2(n_109),
.B1(n_146),
.B2(n_124),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_174),
.A2(n_124),
.B1(n_133),
.B2(n_129),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_185),
.B(n_66),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_200),
.A2(n_136),
.B1(n_113),
.B2(n_150),
.Y(n_245)
);

NOR2x1_ASAP7_75t_SL g246 ( 
.A(n_176),
.B(n_106),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_212),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_247),
.B(n_253),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_218),
.A2(n_178),
.B1(n_170),
.B2(n_144),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_248),
.A2(n_138),
.B1(n_144),
.B2(n_148),
.Y(n_307)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_249),
.Y(n_294)
);

NOR3xp33_ASAP7_75t_L g304 ( 
.A(n_250),
.B(n_263),
.C(n_273),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_202),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_251),
.B(n_255),
.Y(n_281)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_178),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_213),
.B(n_195),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_180),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_260),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_212),
.A2(n_218),
.B(n_210),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_259),
.A2(n_270),
.B(n_208),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_163),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_181),
.C(n_167),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_225),
.C(n_234),
.Y(n_290)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_211),
.Y(n_262)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_243),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_240),
.B(n_181),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_264),
.B(n_224),
.Y(n_298)
);

OAI32xp33_ASAP7_75t_L g265 ( 
.A1(n_239),
.A2(n_172),
.A3(n_207),
.B1(n_203),
.B2(n_208),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_268),
.Y(n_300)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_227),
.Y(n_266)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_225),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_165),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_228),
.B(n_208),
.CI(n_165),
.CON(n_270),
.SN(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_191),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_271),
.B(n_274),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_231),
.B(n_208),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_230),
.B(n_204),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_230),
.B(n_198),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_275),
.B(n_276),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_219),
.B(n_204),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_221),
.B(n_183),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_277),
.B(n_241),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_277),
.B1(n_275),
.B2(n_247),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_295),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_248),
.A2(n_212),
.B1(n_210),
.B2(n_217),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_283),
.A2(n_291),
.B1(n_293),
.B2(n_303),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_250),
.A2(n_246),
.B(n_229),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_284),
.A2(n_287),
.B(n_288),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_259),
.A2(n_229),
.B(n_232),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_259),
.A2(n_220),
.B(n_215),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_290),
.B(n_257),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_277),
.A2(n_244),
.B1(n_245),
.B2(n_227),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_269),
.A2(n_224),
.B1(n_171),
.B2(n_118),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_296),
.B(n_299),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_298),
.B(n_257),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_270),
.A2(n_219),
.B(n_216),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_265),
.A2(n_214),
.B(n_216),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_301),
.A2(n_305),
.B(n_274),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_269),
.A2(n_238),
.B1(n_242),
.B2(n_241),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_265),
.A2(n_105),
.B(n_209),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_266),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_269),
.A2(n_238),
.B1(n_242),
.B2(n_138),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_308),
.A2(n_272),
.B1(n_269),
.B2(n_248),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_253),
.B(n_223),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_309),
.B(n_252),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_326),
.Y(n_343)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_311),
.Y(n_355)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_279),
.Y(n_312)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_312),
.Y(n_357)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_313),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_281),
.B(n_273),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_315),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_281),
.B(n_268),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_316),
.B(n_318),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_292),
.B(n_260),
.Y(n_317)
);

NOR3xp33_ASAP7_75t_L g354 ( 
.A(n_317),
.B(n_323),
.C(n_325),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_258),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_SL g320 ( 
.A(n_283),
.B(n_257),
.C(n_287),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_320),
.A2(n_328),
.B(n_336),
.Y(n_356)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_321),
.Y(n_368)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_280),
.Y(n_322)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_322),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_286),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_292),
.B(n_251),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_324),
.B(n_263),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_282),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_280),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_327),
.Y(n_374)
);

AND2x6_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_270),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_330),
.Y(n_365)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_285),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_331),
.B(n_298),
.C(n_261),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_282),
.B(n_254),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_332),
.B(n_334),
.Y(n_349)
);

CKINVDCx10_ASAP7_75t_R g333 ( 
.A(n_294),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_333),
.Y(n_359)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_285),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_296),
.A2(n_270),
.B(n_271),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_297),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_337),
.B(n_341),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_339),
.Y(n_363)
);

OAI32xp33_ASAP7_75t_L g340 ( 
.A1(n_300),
.A2(n_255),
.A3(n_256),
.B1(n_262),
.B2(n_267),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_340),
.A2(n_306),
.B(n_297),
.Y(n_366)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_289),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_342),
.B(n_290),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_290),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_344),
.B(n_346),
.C(n_361),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_314),
.A2(n_300),
.B1(n_301),
.B2(n_305),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_348),
.A2(n_351),
.B1(n_327),
.B2(n_322),
.Y(n_396)
);

BUFx24_ASAP7_75t_SL g350 ( 
.A(n_337),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_350),
.B(n_352),
.Y(n_391)
);

OAI21xp33_ASAP7_75t_L g351 ( 
.A1(n_336),
.A2(n_335),
.B(n_299),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_304),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_335),
.A2(n_284),
.B(n_287),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_358),
.A2(n_288),
.B(n_278),
.Y(n_389)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_360),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_342),
.B(n_298),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_364),
.B(n_373),
.C(n_264),
.Y(n_392)
);

XOR2x1_ASAP7_75t_L g397 ( 
.A(n_366),
.B(n_375),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_325),
.B(n_306),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_367),
.B(n_369),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_323),
.B(n_309),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_332),
.B(n_276),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_371),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_311),
.B(n_289),
.Y(n_372)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_372),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_320),
.B(n_261),
.C(n_264),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_338),
.B(n_288),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_344),
.B(n_346),
.Y(n_376)
);

MAJx2_ASAP7_75t_L g429 ( 
.A(n_376),
.B(n_381),
.C(n_392),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_343),
.A2(n_314),
.B1(n_338),
.B2(n_329),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_380),
.A2(n_388),
.B1(n_359),
.B2(n_368),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_364),
.B(n_340),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_345),
.Y(n_382)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_382),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_349),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_385),
.Y(n_420)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_349),
.Y(n_384)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_384),
.Y(n_414)
);

AO22x1_ASAP7_75t_SL g385 ( 
.A1(n_343),
.A2(n_328),
.B1(n_310),
.B2(n_291),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_374),
.Y(n_386)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_386),
.Y(n_415)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_374),
.Y(n_387)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_387),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_366),
.A2(n_319),
.B1(n_301),
.B2(n_305),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_389),
.A2(n_395),
.B(n_358),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_354),
.B(n_339),
.Y(n_390)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_390),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_348),
.A2(n_319),
.B1(n_326),
.B2(n_307),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_393),
.A2(n_357),
.B1(n_308),
.B2(n_293),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_361),
.B(n_341),
.C(n_334),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_394),
.B(n_401),
.C(n_370),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_365),
.A2(n_333),
.B(n_330),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_396),
.A2(n_343),
.B1(n_363),
.B2(n_365),
.Y(n_412)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_355),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_400),
.Y(n_431)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_362),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_321),
.C(n_312),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_356),
.B(n_307),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_402),
.B(n_375),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_355),
.B(n_313),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_404),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_362),
.B(n_302),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_405),
.B(n_303),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_378),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_406),
.B(n_407),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_377),
.B(n_347),
.Y(n_407)
);

XNOR2x1_ASAP7_75t_L g434 ( 
.A(n_409),
.B(n_411),
.Y(n_434)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_410),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_412),
.A2(n_427),
.B1(n_385),
.B2(n_404),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_401),
.B(n_356),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_421),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_388),
.A2(n_363),
.B1(n_353),
.B2(n_357),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_417),
.A2(n_428),
.B1(n_386),
.B2(n_387),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_391),
.B(n_359),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_418),
.B(n_205),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_379),
.B(n_370),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_422),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_379),
.B(n_368),
.Y(n_422)
);

XNOR2x1_ASAP7_75t_L g456 ( 
.A(n_424),
.B(n_155),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_376),
.B(n_380),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_425),
.B(n_430),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_384),
.A2(n_362),
.B1(n_294),
.B2(n_266),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_394),
.B(n_223),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_392),
.B(n_249),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_249),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_426),
.A2(n_395),
.B(n_390),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_433),
.A2(n_445),
.B1(n_447),
.B2(n_416),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_419),
.B(n_402),
.C(n_381),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_435),
.B(n_440),
.Y(n_467)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_437),
.Y(n_463)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_431),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_428),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_441),
.B(n_444),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_417),
.A2(n_393),
.B1(n_398),
.B2(n_403),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_442),
.A2(n_427),
.B1(n_406),
.B2(n_409),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_451),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_420),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_408),
.A2(n_400),
.B1(n_405),
.B2(n_397),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_422),
.B(n_397),
.C(n_385),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_446),
.B(n_453),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_SL g447 ( 
.A1(n_414),
.A2(n_389),
.B1(n_106),
.B2(n_186),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_415),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_452),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_410),
.B(n_47),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_189),
.C(n_186),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_423),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_454),
.B(n_455),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_162),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_442),
.A2(n_411),
.B(n_412),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_459),
.A2(n_469),
.B(n_434),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_460),
.A2(n_465),
.B1(n_472),
.B2(n_161),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_434),
.B(n_425),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_461),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_430),
.C(n_413),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_468),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_432),
.C(n_429),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_437),
.A2(n_429),
.B(n_151),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_436),
.B(n_205),
.C(n_143),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_473),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_162),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_439),
.A2(n_79),
.B1(n_75),
.B2(n_62),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_436),
.B(n_199),
.C(n_100),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_448),
.A2(n_199),
.B1(n_19),
.B2(n_162),
.Y(n_474)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_474),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_438),
.B(n_12),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_475),
.B(n_13),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_479),
.B(n_487),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_457),
.A2(n_446),
.B1(n_435),
.B2(n_452),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_480),
.A2(n_485),
.B1(n_28),
.B2(n_11),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_450),
.C(n_453),
.Y(n_481)
);

NOR2xp67_ASAP7_75t_SL g496 ( 
.A(n_481),
.B(n_490),
.Y(n_496)
);

FAx1_ASAP7_75t_SL g482 ( 
.A(n_465),
.B(n_450),
.CI(n_451),
.CON(n_482),
.SN(n_482)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_482),
.B(n_483),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_467),
.B(n_456),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_484),
.B(n_486),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_462),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_458),
.B(n_452),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_489),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_463),
.B(n_468),
.C(n_464),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g491 ( 
.A(n_459),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_471),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_469),
.A2(n_10),
.B(n_12),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_492),
.A2(n_11),
.B(n_1),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_493),
.A2(n_476),
.B1(n_472),
.B2(n_464),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_494),
.B(n_497),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_478),
.A2(n_476),
.B(n_461),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_495),
.A2(n_499),
.B(n_2),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_490),
.B(n_470),
.C(n_473),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_498),
.B(n_503),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_493),
.A2(n_28),
.B(n_10),
.Y(n_499)
);

MAJx2_ASAP7_75t_L g501 ( 
.A(n_481),
.B(n_10),
.C(n_12),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_501),
.B(n_0),
.C(n_2),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_477),
.B(n_9),
.Y(n_503)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_504),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_507),
.B(n_0),
.Y(n_513)
);

AOI322xp5_ASAP7_75t_L g510 ( 
.A1(n_505),
.A2(n_488),
.A3(n_482),
.B1(n_487),
.B2(n_492),
.C1(n_38),
.C2(n_20),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_510),
.A2(n_26),
.B1(n_38),
.B2(n_20),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_506),
.B(n_11),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_511),
.B(n_512),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_496),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_513),
.Y(n_523)
);

INVxp33_ASAP7_75t_L g525 ( 
.A(n_514),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_515),
.A2(n_516),
.B(n_518),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_500),
.B(n_2),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_500),
.A2(n_20),
.B(n_38),
.Y(n_518)
);

AO21x1_ASAP7_75t_L g527 ( 
.A1(n_519),
.A2(n_522),
.B(n_524),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_502),
.C(n_501),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_509),
.B(n_502),
.C(n_508),
.Y(n_524)
);

AOI322xp5_ASAP7_75t_L g526 ( 
.A1(n_520),
.A2(n_513),
.A3(n_38),
.B1(n_26),
.B2(n_33),
.C1(n_27),
.C2(n_4),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_526),
.Y(n_531)
);

AOI322xp5_ASAP7_75t_L g528 ( 
.A1(n_521),
.A2(n_38),
.A3(n_26),
.B1(n_33),
.B2(n_5),
.C1(n_2),
.C2(n_4),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_528),
.A2(n_529),
.B(n_523),
.Y(n_530)
);

AOI322xp5_ASAP7_75t_L g529 ( 
.A1(n_525),
.A2(n_3),
.A3(n_4),
.B1(n_6),
.B2(n_26),
.C1(n_33),
.C2(n_523),
.Y(n_529)
);

AOI322xp5_ASAP7_75t_L g532 ( 
.A1(n_530),
.A2(n_527),
.A3(n_26),
.B1(n_33),
.B2(n_4),
.C1(n_6),
.C2(n_3),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_532),
.A2(n_531),
.B(n_6),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_3),
.B(n_33),
.Y(n_534)
);

BUFx24_ASAP7_75t_SL g535 ( 
.A(n_534),
.Y(n_535)
);


endmodule