module fake_jpeg_865_n_88 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_22),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_17),
.B(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_28),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_30),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_44),
.B(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_37),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_40),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_49),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_31),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_43),
.Y(n_54)
);

FAx1_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_27),
.CI(n_1),
.CON(n_53),
.SN(n_53)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_0),
.C(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_55),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_39),
.B1(n_40),
.B2(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_4),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_40),
.C(n_24),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_3),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_53),
.B1(n_50),
.B2(n_6),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_5),
.C(n_7),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_53),
.B(n_46),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_7),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_4),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_12),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_74),
.C(n_75),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_72),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_69),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_15),
.C(n_19),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_63),
.B1(n_62),
.B2(n_10),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_79),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_11),
.C(n_16),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_76),
.C(n_18),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_81),
.B(n_82),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_83),
.A2(n_78),
.B1(n_9),
.B2(n_10),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_8),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_23),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_8),
.Y(n_88)
);


endmodule