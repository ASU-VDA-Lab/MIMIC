module fake_netlist_5_2322_n_1123 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1123);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1123;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_718;
wire n_671;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_936;
wire n_757;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_1063;
wire n_556;
wire n_1107;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_1016;
wire n_724;
wire n_856;
wire n_546;
wire n_900;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_1096;
wire n_976;
wire n_1095;
wire n_234;
wire n_343;
wire n_428;
wire n_379;
wire n_308;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_223;
wire n_1114;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_1020;
wire n_662;
wire n_459;
wire n_1062;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_962;
wire n_436;
wire n_930;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_974;
wire n_395;
wire n_553;
wire n_432;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_482;
wire n_517;
wire n_342;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_1069;
wire n_236;
wire n_1075;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1101;
wire n_1053;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_1052;
wire n_1116;
wire n_954;
wire n_627;
wire n_767;
wire n_206;
wire n_993;
wire n_217;
wire n_440;
wire n_793;
wire n_478;
wire n_726;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_607;
wire n_237;
wire n_513;
wire n_425;
wire n_407;
wire n_527;
wire n_679;
wire n_710;
wire n_707;
wire n_832;
wire n_695;
wire n_795;
wire n_857;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_1027;
wire n_490;
wire n_805;
wire n_971;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_895;
wire n_644;
wire n_728;
wire n_1037;
wire n_202;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_1038;
wire n_409;
wire n_797;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_536;
wire n_531;
wire n_1004;
wire n_935;
wire n_242;
wire n_817;
wire n_1032;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_189),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_116),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_104),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_56),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_187),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_152),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_67),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_105),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_24),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_2),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_33),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_44),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_45),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_98),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_35),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_22),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_148),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_28),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_115),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_27),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_23),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_5),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_191),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_97),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_142),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_165),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_72),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_136),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_188),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_80),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_192),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_122),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_195),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_39),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_17),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_55),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_111),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_38),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_163),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_144),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_194),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_46),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_124),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_26),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_181),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_0),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_183),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_10),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_184),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_153),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_156),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_43),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_39),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_130),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_157),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_42),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_66),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_85),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_6),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_77),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_128),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_93),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_50),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_186),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_190),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_54),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

INVxp67_ASAP7_75t_SL g267 ( 
.A(n_200),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_216),
.Y(n_269)
);

INVxp33_ASAP7_75t_SL g270 ( 
.A(n_206),
.Y(n_270)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_253),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_232),
.Y(n_272)
);

BUFx2_ASAP7_75t_SL g273 ( 
.A(n_229),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_237),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_241),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_212),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_215),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_198),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_204),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_233),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_209),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_223),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_228),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_217),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_230),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_197),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_234),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_250),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_236),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_206),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_221),
.Y(n_294)
);

INVxp33_ASAP7_75t_SL g295 ( 
.A(n_207),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_207),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_238),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_239),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_222),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_248),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_249),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_224),
.Y(n_302)
);

INVxp33_ASAP7_75t_SL g303 ( 
.A(n_208),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_208),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_248),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_259),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_261),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_225),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_248),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_248),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_205),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_211),
.Y(n_314)
);

INVxp33_ASAP7_75t_SL g315 ( 
.A(n_210),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_280),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_311),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

NAND2x1p5_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_220),
.Y(n_319)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_305),
.A2(n_227),
.B(n_226),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_280),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_298),
.B(n_245),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_305),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_305),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_273),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_292),
.B(n_199),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_289),
.A2(n_218),
.B1(n_247),
.B2(n_219),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_312),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_312),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_300),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_312),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_301),
.B(n_199),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_300),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_267),
.A2(n_258),
.B1(n_210),
.B2(n_255),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_278),
.B(n_279),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_266),
.Y(n_337)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_300),
.Y(n_338)
);

AND2x4_ASAP7_75t_L g339 ( 
.A(n_281),
.B(n_201),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_300),
.Y(n_340)
);

AND2x2_ASAP7_75t_SL g341 ( 
.A(n_289),
.B(n_52),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_300),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_287),
.B(n_201),
.Y(n_343)
);

INVxp33_ASAP7_75t_SL g344 ( 
.A(n_294),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_266),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_282),
.B(n_202),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_300),
.Y(n_347)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_313),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_282),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_284),
.Y(n_350)
);

INVx6_ASAP7_75t_L g351 ( 
.A(n_313),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_284),
.B(n_202),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_299),
.B(n_240),
.Y(n_354)
);

AND2x6_ASAP7_75t_L g355 ( 
.A(n_285),
.B(n_53),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_291),
.B(n_203),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_302),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_285),
.Y(n_358)
);

OA21x2_ASAP7_75t_L g359 ( 
.A1(n_286),
.A2(n_258),
.B(n_231),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_268),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_271),
.B(n_203),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_268),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_309),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_272),
.Y(n_364)
);

AND2x6_ASAP7_75t_L g365 ( 
.A(n_286),
.B(n_57),
.Y(n_365)
);

AND2x2_ASAP7_75t_SL g366 ( 
.A(n_288),
.B(n_58),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_270),
.A2(n_303),
.B1(n_315),
.B2(n_295),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_288),
.B(n_242),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_290),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_290),
.B(n_231),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_332),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_297),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_369),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_316),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_369),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_297),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_348),
.B(n_304),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_316),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_369),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_343),
.B(n_306),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_369),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_369),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_354),
.B(n_306),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_322),
.B(n_252),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_348),
.B(n_319),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_361),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_317),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_317),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_321),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_341),
.A2(n_262),
.B1(n_296),
.B2(n_293),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_318),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_341),
.A2(n_296),
.B1(n_314),
.B2(n_273),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_318),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_349),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_349),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_350),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_339),
.B(n_307),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_350),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_321),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_323),
.Y(n_404)
);

AND2x6_ASAP7_75t_L g405 ( 
.A(n_333),
.B(n_307),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_326),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_341),
.A2(n_314),
.B1(n_269),
.B2(n_264),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_337),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_330),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g410 ( 
.A(n_333),
.B(n_308),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_358),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_361),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_358),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_337),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_323),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_345),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_345),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_324),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_324),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_360),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_360),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_362),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_328),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_328),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_362),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_329),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_322),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_364),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_364),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_329),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_331),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_331),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_330),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_339),
.B(n_272),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_319),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_330),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_334),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_334),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_327),
.A2(n_263),
.B1(n_257),
.B2(n_260),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_326),
.A2(n_263),
.B1(n_257),
.B2(n_260),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_334),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_338),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_340),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_340),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_387),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_385),
.B(n_366),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_382),
.B(n_366),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_414),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_406),
.B(n_366),
.Y(n_450)
);

NAND2xp33_ASAP7_75t_SL g451 ( 
.A(n_407),
.B(n_325),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_371),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_371),
.B(n_344),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_414),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_375),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_L g456 ( 
.A(n_405),
.B(n_355),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_405),
.B(n_326),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_405),
.B(n_336),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_375),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_374),
.B(n_357),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_405),
.A2(n_365),
.B1(n_355),
.B2(n_359),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_380),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_405),
.B(n_368),
.Y(n_463)
);

INVxp33_ASAP7_75t_L g464 ( 
.A(n_377),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_405),
.B(n_359),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_405),
.B(n_359),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_410),
.B(n_359),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_380),
.Y(n_468)
);

NOR3xp33_ASAP7_75t_L g469 ( 
.A(n_393),
.B(n_367),
.C(n_335),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_410),
.B(n_357),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_410),
.B(n_357),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_406),
.B(n_348),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_392),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_392),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_372),
.B(n_348),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_410),
.B(n_339),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_410),
.B(n_346),
.Y(n_477)
);

NAND2x1_ASAP7_75t_L g478 ( 
.A(n_410),
.B(n_355),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_372),
.B(n_348),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_387),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_L g481 ( 
.A(n_389),
.B(n_353),
.C(n_346),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_412),
.B(n_344),
.Y(n_482)
);

BUFx5_ASAP7_75t_L g483 ( 
.A(n_410),
.Y(n_483)
);

INVx8_ASAP7_75t_L g484 ( 
.A(n_435),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_L g485 ( 
.A(n_436),
.B(n_355),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_403),
.Y(n_486)
);

NAND3xp33_ASAP7_75t_L g487 ( 
.A(n_441),
.B(n_353),
.C(n_346),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_377),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_386),
.B(n_325),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_417),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_440),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_378),
.B(n_353),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_378),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_403),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_435),
.B(n_348),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_417),
.B(n_370),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_435),
.B(n_363),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_401),
.B(n_319),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_431),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_401),
.B(n_370),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_408),
.B(n_351),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_418),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_387),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_418),
.B(n_421),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_421),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_431),
.Y(n_506)
);

BUFx4_ASAP7_75t_L g507 ( 
.A(n_386),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_422),
.B(n_351),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_422),
.B(n_370),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_423),
.B(n_426),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_423),
.B(n_351),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_404),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_426),
.Y(n_513)
);

OR2x2_ASAP7_75t_SL g514 ( 
.A(n_395),
.B(n_351),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_429),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_429),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_397),
.B(n_320),
.Y(n_517)
);

NOR3xp33_ASAP7_75t_L g518 ( 
.A(n_428),
.B(n_310),
.C(n_308),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_L g519 ( 
.A(n_430),
.B(n_355),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_388),
.B(n_310),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_430),
.B(n_235),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_397),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_398),
.B(n_320),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_398),
.B(n_355),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_399),
.B(n_355),
.Y(n_525)
);

NOR3xp33_ASAP7_75t_L g526 ( 
.A(n_379),
.B(n_275),
.C(n_274),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_400),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_399),
.B(n_365),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_390),
.B(n_365),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_390),
.B(n_365),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_391),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_484),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_499),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_391),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_452),
.Y(n_535)
);

AND2x6_ASAP7_75t_L g536 ( 
.A(n_465),
.B(n_373),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_499),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_448),
.A2(n_396),
.B1(n_394),
.B2(n_373),
.Y(n_538)
);

OR2x6_ASAP7_75t_L g539 ( 
.A(n_488),
.B(n_274),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_493),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_482),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_506),
.Y(n_542)
);

AO22x2_ASAP7_75t_L g543 ( 
.A1(n_469),
.A2(n_396),
.B1(n_394),
.B2(n_276),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_491),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_506),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_527),
.B(n_400),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_516),
.Y(n_547)
);

OAI221xp5_ASAP7_75t_L g548 ( 
.A1(n_492),
.A2(n_411),
.B1(n_402),
.B2(n_413),
.C(n_277),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_512),
.Y(n_549)
);

AO22x2_ASAP7_75t_L g550 ( 
.A1(n_450),
.A2(n_276),
.B1(n_277),
.B2(n_275),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_516),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_522),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_449),
.Y(n_553)
);

AO22x2_ASAP7_75t_L g554 ( 
.A1(n_450),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_512),
.Y(n_555)
);

AO22x2_ASAP7_75t_L g556 ( 
.A1(n_447),
.A2(n_489),
.B1(n_487),
.B2(n_481),
.Y(n_556)
);

NAND2x1p5_ASAP7_75t_L g557 ( 
.A(n_495),
.B(n_402),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_464),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_454),
.Y(n_559)
);

NOR2xp67_ASAP7_75t_L g560 ( 
.A(n_482),
.B(n_411),
.Y(n_560)
);

OAI221xp5_ASAP7_75t_L g561 ( 
.A1(n_496),
.A2(n_413),
.B1(n_235),
.B2(n_264),
.C(n_433),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_510),
.B(n_376),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_531),
.B(n_443),
.Y(n_563)
);

OAI221xp5_ASAP7_75t_L g564 ( 
.A1(n_509),
.A2(n_244),
.B1(n_246),
.B2(n_256),
.C(n_416),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_510),
.B(n_376),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_453),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_490),
.B(n_381),
.Y(n_567)
);

AO22x2_ASAP7_75t_L g568 ( 
.A1(n_498),
.A2(n_4),
.B1(n_1),
.B2(n_3),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_497),
.B(n_404),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_484),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_455),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_497),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_484),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_475),
.A2(n_365),
.B1(n_383),
.B2(n_381),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_502),
.B(n_505),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_513),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_455),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_515),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_462),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_462),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_508),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_468),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_468),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_460),
.B(n_443),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_473),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_473),
.Y(n_586)
);

NOR2x1p5_ASAP7_75t_L g587 ( 
.A(n_470),
.B(n_383),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_518),
.Y(n_588)
);

BUFx4f_ASAP7_75t_L g589 ( 
.A(n_446),
.Y(n_589)
);

AO22x2_ASAP7_75t_L g590 ( 
.A1(n_475),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_590)
);

NAND2x1p5_ASAP7_75t_L g591 ( 
.A(n_495),
.B(n_384),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_474),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_479),
.A2(n_384),
.B1(n_438),
.B2(n_442),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_474),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_457),
.A2(n_442),
.B1(n_439),
.B2(n_365),
.Y(n_595)
);

AO22x2_ASAP7_75t_L g596 ( 
.A1(n_507),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_596)
);

AO22x2_ASAP7_75t_L g597 ( 
.A1(n_472),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_486),
.Y(n_598)
);

OAI221xp5_ASAP7_75t_L g599 ( 
.A1(n_526),
.A2(n_424),
.B1(n_416),
.B2(n_425),
.C(n_419),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_504),
.B(n_439),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_569),
.B(n_508),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_558),
.Y(n_602)
);

BUFx8_ASAP7_75t_L g603 ( 
.A(n_544),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_581),
.B(n_458),
.Y(n_604)
);

NOR2xp67_ASAP7_75t_L g605 ( 
.A(n_535),
.B(n_501),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_532),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_532),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_534),
.B(n_511),
.Y(n_608)
);

AOI221xp5_ASAP7_75t_L g609 ( 
.A1(n_588),
.A2(n_451),
.B1(n_521),
.B2(n_501),
.C(n_511),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_589),
.A2(n_456),
.B(n_461),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_560),
.B(n_471),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_542),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_589),
.A2(n_461),
.B(n_485),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_545),
.Y(n_614)
);

AO21x1_ASAP7_75t_L g615 ( 
.A1(n_562),
.A2(n_523),
.B(n_517),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_572),
.B(n_520),
.Y(n_616)
);

O2A1O1Ixp5_ASAP7_75t_L g617 ( 
.A1(n_565),
.A2(n_523),
.B(n_517),
.C(n_467),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_533),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_600),
.A2(n_519),
.B(n_466),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_537),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_534),
.B(n_486),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_541),
.B(n_483),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_566),
.B(n_514),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_575),
.A2(n_463),
.B(n_478),
.Y(n_624)
);

O2A1O1Ixp33_ASAP7_75t_SL g625 ( 
.A1(n_547),
.A2(n_477),
.B(n_476),
.C(n_529),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_551),
.B(n_494),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_546),
.B(n_483),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_595),
.A2(n_480),
.B(n_446),
.Y(n_628)
);

A2O1A1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_553),
.A2(n_530),
.B(n_528),
.C(n_525),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_550),
.B(n_494),
.Y(n_630)
);

NAND2x1p5_ASAP7_75t_L g631 ( 
.A(n_570),
.B(n_446),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_532),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_540),
.B(n_459),
.Y(n_633)
);

NOR2xp67_ASAP7_75t_L g634 ( 
.A(n_561),
.B(n_524),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_550),
.B(n_459),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_567),
.A2(n_480),
.B(n_446),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_574),
.A2(n_480),
.B(n_503),
.Y(n_637)
);

OA22x2_ASAP7_75t_L g638 ( 
.A1(n_539),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_571),
.Y(n_639)
);

OA22x2_ASAP7_75t_L g640 ( 
.A1(n_539),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_546),
.B(n_480),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_559),
.B(n_576),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_571),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_549),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_543),
.B(n_419),
.Y(n_645)
);

NOR3xp33_ASAP7_75t_L g646 ( 
.A(n_564),
.B(n_424),
.C(n_420),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_549),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_578),
.B(n_552),
.Y(n_648)
);

BUFx4f_ASAP7_75t_L g649 ( 
.A(n_563),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_543),
.B(n_420),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_584),
.A2(n_483),
.B(n_409),
.Y(n_651)
);

O2A1O1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_548),
.A2(n_599),
.B(n_555),
.C(n_582),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_584),
.A2(n_483),
.B(n_409),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_556),
.A2(n_483),
.B1(n_365),
.B2(n_437),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_555),
.Y(n_655)
);

NAND2x1p5_ASAP7_75t_L g656 ( 
.A(n_570),
.B(n_437),
.Y(n_656)
);

OAI21x1_ASAP7_75t_SL g657 ( 
.A1(n_573),
.A2(n_445),
.B(n_434),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g658 ( 
.A1(n_538),
.A2(n_445),
.B(n_434),
.Y(n_658)
);

O2A1O1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_580),
.A2(n_425),
.B(n_427),
.C(n_432),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_577),
.A2(n_483),
.B(n_594),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_563),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_556),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_596),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_583),
.B(n_437),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_601),
.B(n_577),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_648),
.B(n_594),
.Y(n_666)
);

BUFx12f_ASAP7_75t_L g667 ( 
.A(n_603),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_605),
.B(n_573),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_604),
.B(n_642),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_644),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_604),
.B(n_598),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_609),
.B(n_598),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_647),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_655),
.Y(n_674)
);

BUFx8_ASAP7_75t_L g675 ( 
.A(n_606),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_649),
.B(n_557),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_645),
.B(n_554),
.Y(n_677)
);

INVxp33_ASAP7_75t_SL g678 ( 
.A(n_623),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_602),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_616),
.B(n_579),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_641),
.B(n_608),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_606),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_650),
.B(n_554),
.Y(n_683)
);

AND3x1_ASAP7_75t_SL g684 ( 
.A(n_663),
.B(n_596),
.C(n_568),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_603),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_639),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_662),
.B(n_590),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_649),
.A2(n_591),
.B1(n_587),
.B2(n_593),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_633),
.B(n_592),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_606),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_612),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_661),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_643),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_607),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_626),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_621),
.B(n_585),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_627),
.A2(n_634),
.B1(n_622),
.B2(n_614),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_618),
.B(n_586),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_607),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_626),
.Y(n_700)
);

NAND2x1p5_ASAP7_75t_L g701 ( 
.A(n_613),
.B(n_427),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_607),
.B(n_387),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_611),
.B(n_387),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_619),
.A2(n_536),
.B(n_432),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_620),
.B(n_590),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_L g706 ( 
.A(n_610),
.B(n_536),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_632),
.B(n_597),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_632),
.B(n_597),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_630),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_630),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_635),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_635),
.B(n_568),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_652),
.B(n_536),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_638),
.B(n_536),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_631),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_617),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_631),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_654),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_624),
.B(n_409),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_629),
.B(n_12),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_664),
.B(n_646),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_638),
.A2(n_415),
.B1(n_409),
.B2(n_444),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_720),
.A2(n_640),
.B1(n_615),
.B2(n_658),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_679),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_717),
.Y(n_725)
);

AOI21x1_ASAP7_75t_SL g726 ( 
.A1(n_721),
.A2(n_640),
.B(n_625),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_669),
.B(n_636),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_670),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_681),
.B(n_659),
.Y(n_729)
);

NAND3xp33_ASAP7_75t_L g730 ( 
.A(n_680),
.B(n_658),
.C(n_628),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_682),
.Y(n_731)
);

AOI21x1_ASAP7_75t_L g732 ( 
.A1(n_719),
.A2(n_703),
.B(n_713),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_670),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_667),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_673),
.Y(n_735)
);

INVx5_ASAP7_75t_L g736 ( 
.A(n_717),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_673),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_666),
.B(n_637),
.Y(n_738)
);

O2A1O1Ixp5_ASAP7_75t_L g739 ( 
.A1(n_716),
.A2(n_660),
.B(n_653),
.C(n_651),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_678),
.A2(n_656),
.B1(n_409),
.B2(n_444),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_706),
.A2(n_704),
.B(n_672),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_717),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_689),
.B(n_656),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_SL g744 ( 
.A1(n_718),
.A2(n_657),
.B1(n_14),
.B2(n_15),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_693),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_675),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_SL g747 ( 
.A(n_685),
.B(n_415),
.Y(n_747)
);

INVx5_ASAP7_75t_L g748 ( 
.A(n_717),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_678),
.B(n_13),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_687),
.B(n_14),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_696),
.B(n_15),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_674),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_675),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_674),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_693),
.Y(n_755)
);

INVx6_ASAP7_75t_L g756 ( 
.A(n_675),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_718),
.B(n_16),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_687),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_691),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_706),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_686),
.B(n_59),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_686),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_682),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_677),
.B(n_19),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_698),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_717),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_677),
.B(n_20),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_R g768 ( 
.A(n_685),
.B(n_60),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_665),
.B(n_21),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_700),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_711),
.B(n_21),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_711),
.B(n_22),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_682),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_716),
.A2(n_444),
.B(n_415),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_683),
.B(n_23),
.Y(n_775)
);

O2A1O1Ixp5_ASAP7_75t_SL g776 ( 
.A1(n_710),
.A2(n_712),
.B(n_702),
.C(n_695),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_683),
.B(n_692),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_671),
.A2(n_676),
.B(n_688),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_695),
.B(n_24),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_682),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_709),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_714),
.B(n_61),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_707),
.B(n_25),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_667),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_700),
.B(n_25),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_709),
.Y(n_786)
);

OAI21x1_ASAP7_75t_L g787 ( 
.A1(n_701),
.A2(n_444),
.B(n_415),
.Y(n_787)
);

AOI21x1_ASAP7_75t_L g788 ( 
.A1(n_708),
.A2(n_444),
.B(n_415),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_710),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_705),
.B(n_26),
.Y(n_790)
);

CKINVDCx11_ASAP7_75t_R g791 ( 
.A(n_682),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_728),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_777),
.B(n_764),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_741),
.A2(n_727),
.B(n_738),
.Y(n_794)
);

OA21x2_ASAP7_75t_L g795 ( 
.A1(n_774),
.A2(n_697),
.B(n_714),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_778),
.A2(n_701),
.B(n_722),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_733),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_730),
.A2(n_701),
.B(n_668),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_767),
.B(n_705),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_760),
.B(n_715),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_770),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_765),
.B(n_715),
.Y(n_802)
);

O2A1O1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_760),
.A2(n_694),
.B(n_684),
.C(n_29),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_739),
.A2(n_699),
.B(n_690),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_SL g805 ( 
.A1(n_758),
.A2(n_690),
.B(n_694),
.C(n_699),
.Y(n_805)
);

BUFx10_ASAP7_75t_L g806 ( 
.A(n_756),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_734),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_791),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_724),
.B(n_690),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_770),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_751),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_811)
);

INVxp33_ASAP7_75t_L g812 ( 
.A(n_749),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_736),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_SL g814 ( 
.A1(n_757),
.A2(n_699),
.B1(n_31),
.B2(n_32),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_791),
.Y(n_815)
);

OA21x2_ASAP7_75t_L g816 ( 
.A1(n_787),
.A2(n_338),
.B(n_30),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_723),
.A2(n_699),
.B(n_31),
.C(n_32),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_735),
.Y(n_818)
);

OA21x2_ASAP7_75t_L g819 ( 
.A1(n_787),
.A2(n_338),
.B(n_30),
.Y(n_819)
);

A2O1A1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_723),
.A2(n_699),
.B(n_34),
.C(n_35),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_729),
.A2(n_342),
.B(n_340),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_769),
.B(n_33),
.Y(n_822)
);

INVxp33_ASAP7_75t_L g823 ( 
.A(n_743),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_758),
.A2(n_338),
.B1(n_36),
.B2(n_37),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_775),
.B(n_750),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_779),
.B(n_34),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_736),
.A2(n_342),
.B(n_340),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_761),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_786),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_790),
.B(n_62),
.Y(n_830)
);

OA21x2_ASAP7_75t_L g831 ( 
.A1(n_732),
.A2(n_40),
.B(n_41),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_786),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_789),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_780),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_737),
.B(n_40),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_757),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_836)
);

NAND3xp33_ASAP7_75t_L g837 ( 
.A(n_744),
.B(n_347),
.C(n_342),
.Y(n_837)
);

AOI221xp5_ASAP7_75t_L g838 ( 
.A1(n_771),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.C(n_47),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_752),
.B(n_47),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_785),
.B(n_48),
.Y(n_840)
);

OAI21x1_ASAP7_75t_SL g841 ( 
.A1(n_772),
.A2(n_48),
.B(n_49),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_782),
.B(n_63),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_SL g843 ( 
.A(n_734),
.B(n_340),
.Y(n_843)
);

A2O1A1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_761),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_725),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_781),
.B(n_51),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_761),
.A2(n_64),
.B(n_65),
.C(n_68),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_756),
.A2(n_347),
.B1(n_342),
.B2(n_71),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_782),
.B(n_69),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_783),
.B(n_759),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_754),
.B(n_70),
.Y(n_851)
);

CKINVDCx6p67_ASAP7_75t_R g852 ( 
.A(n_753),
.Y(n_852)
);

AND2x2_ASAP7_75t_SL g853 ( 
.A(n_747),
.B(n_73),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_814),
.A2(n_824),
.B1(n_838),
.B2(n_837),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_792),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_SL g856 ( 
.A1(n_853),
.A2(n_768),
.B1(n_756),
.B2(n_753),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_806),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_833),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_797),
.Y(n_859)
);

BUFx12f_ASAP7_75t_L g860 ( 
.A(n_807),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_822),
.A2(n_768),
.B1(n_746),
.B2(n_762),
.Y(n_861)
);

OAI22x1_ASAP7_75t_L g862 ( 
.A1(n_800),
.A2(n_746),
.B1(n_784),
.B2(n_788),
.Y(n_862)
);

INVx5_ASAP7_75t_L g863 ( 
.A(n_806),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_793),
.B(n_725),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_812),
.A2(n_784),
.B1(n_745),
.B2(n_755),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_818),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_810),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_817),
.A2(n_748),
.B1(n_736),
.B2(n_740),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_829),
.Y(n_869)
);

HB1xp67_ASAP7_75t_SL g870 ( 
.A(n_807),
.Y(n_870)
);

BUFx4f_ASAP7_75t_L g871 ( 
.A(n_853),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_850),
.B(n_745),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_812),
.A2(n_755),
.B1(n_742),
.B2(n_725),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_832),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_799),
.B(n_742),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_823),
.B(n_742),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_808),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_826),
.A2(n_841),
.B1(n_840),
.B2(n_800),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_SL g879 ( 
.A1(n_808),
.A2(n_736),
.B1(n_748),
.B2(n_766),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_817),
.A2(n_748),
.B1(n_736),
.B2(n_766),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_SL g881 ( 
.A1(n_815),
.A2(n_748),
.B1(n_766),
.B2(n_763),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_825),
.A2(n_780),
.B1(n_763),
.B2(n_731),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_SL g883 ( 
.A1(n_836),
.A2(n_726),
.B(n_773),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_852),
.Y(n_884)
);

INVx4_ASAP7_75t_L g885 ( 
.A(n_806),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_801),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_SL g887 ( 
.A1(n_811),
.A2(n_773),
.B(n_776),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_SL g888 ( 
.A(n_809),
.B(n_731),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_823),
.A2(n_763),
.B1(n_731),
.B2(n_748),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_SL g890 ( 
.A1(n_803),
.A2(n_773),
.B(n_75),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_796),
.A2(n_773),
.B1(n_76),
.B2(n_78),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_801),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_834),
.B(n_74),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_802),
.B(n_79),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_852),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_820),
.A2(n_347),
.B1(n_342),
.B2(n_83),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_835),
.A2(n_81),
.B1(n_82),
.B2(n_84),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_801),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_835),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_899)
);

INVx5_ASAP7_75t_SL g900 ( 
.A(n_843),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_845),
.B(n_89),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_820),
.A2(n_347),
.B1(n_91),
.B2(n_92),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_858),
.B(n_794),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_890),
.A2(n_828),
.B1(n_844),
.B2(n_848),
.Y(n_904)
);

AND2x2_ASAP7_75t_SL g905 ( 
.A(n_871),
.B(n_831),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_876),
.B(n_846),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_855),
.Y(n_907)
);

A2O1A1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_871),
.A2(n_844),
.B(n_828),
.C(n_902),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_855),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_878),
.A2(n_847),
.B(n_798),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_859),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_877),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_854),
.A2(n_849),
.B1(n_842),
.B2(n_830),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_896),
.A2(n_805),
.B(n_847),
.C(n_839),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_887),
.A2(n_805),
.B(n_839),
.C(n_821),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_864),
.B(n_815),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_867),
.B(n_845),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_877),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_869),
.Y(n_919)
);

NOR2x1_ASAP7_75t_SL g920 ( 
.A(n_863),
.B(n_813),
.Y(n_920)
);

OR2x6_ASAP7_75t_L g921 ( 
.A(n_862),
.B(n_804),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_870),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_875),
.B(n_845),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_854),
.A2(n_813),
.B1(n_795),
.B2(n_851),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_874),
.B(n_851),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_857),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_860),
.Y(n_927)
);

OA21x2_ASAP7_75t_L g928 ( 
.A1(n_889),
.A2(n_827),
.B(n_831),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_SL g929 ( 
.A1(n_880),
.A2(n_831),
.B(n_795),
.C(n_816),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_SL g930 ( 
.A1(n_891),
.A2(n_795),
.B(n_819),
.C(n_816),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_878),
.A2(n_819),
.B(n_816),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_866),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_883),
.A2(n_819),
.B(n_94),
.C(n_95),
.Y(n_933)
);

INVx5_ASAP7_75t_SL g934 ( 
.A(n_860),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_919),
.B(n_886),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_906),
.B(n_876),
.Y(n_936)
);

INVxp67_ASAP7_75t_SL g937 ( 
.A(n_903),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_919),
.B(n_892),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_907),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_909),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_917),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_923),
.B(n_898),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_922),
.B(n_888),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_932),
.Y(n_944)
);

NOR2x1p5_ASAP7_75t_L g945 ( 
.A(n_927),
.B(n_884),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_917),
.Y(n_946)
);

AOI221xp5_ASAP7_75t_L g947 ( 
.A1(n_910),
.A2(n_861),
.B1(n_865),
.B2(n_897),
.C(n_899),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_912),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_906),
.B(n_872),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_911),
.B(n_873),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_926),
.B(n_882),
.Y(n_951)
);

INVx4_ASAP7_75t_L g952 ( 
.A(n_918),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_918),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_921),
.B(n_873),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_921),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_925),
.B(n_865),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_916),
.B(n_882),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_939),
.Y(n_958)
);

INVx1_ASAP7_75t_SL g959 ( 
.A(n_948),
.Y(n_959)
);

NAND3xp33_ASAP7_75t_L g960 ( 
.A(n_947),
.B(n_908),
.C(n_904),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_937),
.B(n_921),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_936),
.B(n_934),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_939),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_940),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_946),
.B(n_905),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_948),
.Y(n_966)
);

OAI21x1_ASAP7_75t_L g967 ( 
.A1(n_955),
.A2(n_931),
.B(n_928),
.Y(n_967)
);

INVx4_ASAP7_75t_SL g968 ( 
.A(n_951),
.Y(n_968)
);

INVxp67_ASAP7_75t_SL g969 ( 
.A(n_955),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_949),
.B(n_925),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_952),
.Y(n_971)
);

INVx4_ASAP7_75t_SL g972 ( 
.A(n_951),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_940),
.Y(n_973)
);

AO22x2_ASAP7_75t_L g974 ( 
.A1(n_955),
.A2(n_924),
.B1(n_868),
.B2(n_895),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_958),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_968),
.B(n_955),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_968),
.B(n_941),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_968),
.B(n_952),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_961),
.B(n_950),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_960),
.B(n_957),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_958),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_968),
.B(n_952),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_966),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_960),
.B(n_957),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_964),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_961),
.B(n_950),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_964),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_972),
.B(n_965),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_988),
.B(n_972),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_975),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_981),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_983),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_985),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_979),
.B(n_959),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_985),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_987),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_SL g997 ( 
.A(n_989),
.B(n_978),
.Y(n_997)
);

OAI32xp33_ASAP7_75t_L g998 ( 
.A1(n_992),
.A2(n_984),
.A3(n_980),
.B1(n_988),
.B2(n_986),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_992),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_990),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_989),
.B(n_972),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_994),
.A2(n_982),
.B(n_978),
.Y(n_1002)
);

NOR2x1_ASAP7_75t_SL g1003 ( 
.A(n_1001),
.B(n_982),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_997),
.B(n_972),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_999),
.B(n_991),
.Y(n_1005)
);

INVxp67_ASAP7_75t_SL g1006 ( 
.A(n_999),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_1000),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_1002),
.B(n_979),
.Y(n_1008)
);

OAI221xp5_ASAP7_75t_L g1009 ( 
.A1(n_998),
.A2(n_962),
.B1(n_976),
.B2(n_986),
.C(n_908),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_997),
.B(n_934),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_1001),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_1001),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_1011),
.B(n_977),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1006),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1005),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1007),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1008),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1003),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1012),
.B(n_977),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1012),
.B(n_993),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1014),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_1017),
.B(n_1010),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_1018),
.A2(n_1004),
.B1(n_1009),
.B2(n_974),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1017),
.B(n_995),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_1016),
.B(n_976),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1013),
.B(n_996),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1020),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_1019),
.B(n_996),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1026),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1021),
.Y(n_1030)
);

NAND4xp75_ASAP7_75t_L g1031 ( 
.A(n_1022),
.B(n_1015),
.C(n_965),
.D(n_943),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_1023),
.A2(n_1025),
.B(n_1024),
.Y(n_1032)
);

NAND3xp33_ASAP7_75t_L g1033 ( 
.A(n_1027),
.B(n_899),
.C(n_897),
.Y(n_1033)
);

NOR2xp67_ASAP7_75t_L g1034 ( 
.A(n_1028),
.B(n_971),
.Y(n_1034)
);

NAND4xp25_ASAP7_75t_L g1035 ( 
.A(n_1025),
.B(n_856),
.C(n_861),
.D(n_913),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1034),
.B(n_969),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_1029),
.B(n_987),
.Y(n_1037)
);

NAND2x1p5_ASAP7_75t_L g1038 ( 
.A(n_1030),
.B(n_945),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1032),
.B(n_966),
.Y(n_1039)
);

OAI221xp5_ASAP7_75t_L g1040 ( 
.A1(n_1033),
.A2(n_971),
.B1(n_933),
.B2(n_891),
.C(n_953),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1031),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1035),
.B(n_945),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1032),
.B(n_934),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_SL g1044 ( 
.A1(n_1032),
.A2(n_974),
.B1(n_971),
.B2(n_967),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_1029),
.B(n_970),
.Y(n_1045)
);

INVxp67_ASAP7_75t_L g1046 ( 
.A(n_1031),
.Y(n_1046)
);

NOR3xp33_ASAP7_75t_L g1047 ( 
.A(n_1046),
.B(n_1043),
.C(n_1041),
.Y(n_1047)
);

OAI21xp33_ASAP7_75t_L g1048 ( 
.A1(n_1039),
.A2(n_974),
.B(n_954),
.Y(n_1048)
);

AOI221xp5_ASAP7_75t_L g1049 ( 
.A1(n_1036),
.A2(n_1044),
.B1(n_1042),
.B2(n_1040),
.C(n_1045),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_1038),
.B(n_952),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_L g1051 ( 
.A(n_1037),
.B(n_894),
.C(n_893),
.Y(n_1051)
);

NAND4xp25_ASAP7_75t_L g1052 ( 
.A(n_1039),
.B(n_954),
.C(n_914),
.D(n_885),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_1043),
.A2(n_974),
.B1(n_967),
.B2(n_885),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1036),
.Y(n_1054)
);

AOI211xp5_ASAP7_75t_SL g1055 ( 
.A1(n_1046),
.A2(n_857),
.B(n_929),
.C(n_901),
.Y(n_1055)
);

AOI21xp33_ASAP7_75t_SL g1056 ( 
.A1(n_1046),
.A2(n_915),
.B(n_905),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_1043),
.A2(n_863),
.B1(n_956),
.B2(n_963),
.Y(n_1057)
);

OAI22xp33_ASAP7_75t_SL g1058 ( 
.A1(n_1050),
.A2(n_963),
.B1(n_973),
.B2(n_863),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_1054),
.B(n_973),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1047),
.B(n_942),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1049),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1051),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1056),
.A2(n_881),
.B(n_879),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1057),
.B(n_944),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_L g1065 ( 
.A(n_1055),
.B(n_863),
.C(n_938),
.Y(n_1065)
);

NAND4xp75_ASAP7_75t_L g1066 ( 
.A(n_1061),
.B(n_1052),
.C(n_1048),
.D(n_1053),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1060),
.Y(n_1067)
);

NOR2x1_ASAP7_75t_L g1068 ( 
.A(n_1062),
.B(n_935),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1059),
.B(n_944),
.Y(n_1069)
);

AND2x2_ASAP7_75t_SL g1070 ( 
.A(n_1064),
.B(n_1058),
.Y(n_1070)
);

NOR2xp67_ASAP7_75t_L g1071 ( 
.A(n_1065),
.B(n_90),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1063),
.A2(n_900),
.B1(n_942),
.B2(n_935),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_1061),
.A2(n_900),
.B1(n_938),
.B2(n_889),
.Y(n_1073)
);

XOR2x2_ASAP7_75t_L g1074 ( 
.A(n_1061),
.B(n_920),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_1067),
.A2(n_900),
.B1(n_928),
.B2(n_930),
.Y(n_1075)
);

AOI322xp5_ASAP7_75t_L g1076 ( 
.A1(n_1068),
.A2(n_930),
.A3(n_929),
.B1(n_928),
.B2(n_101),
.C1(n_102),
.C2(n_103),
.Y(n_1076)
);

XNOR2xp5_ASAP7_75t_L g1077 ( 
.A(n_1074),
.B(n_96),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_1070),
.Y(n_1078)
);

NOR2x1_ASAP7_75t_L g1079 ( 
.A(n_1066),
.B(n_1071),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_1072),
.B(n_99),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1073),
.A2(n_100),
.B(n_106),
.Y(n_1081)
);

AND4x1_ASAP7_75t_L g1082 ( 
.A(n_1069),
.B(n_107),
.C(n_108),
.D(n_109),
.Y(n_1082)
);

NOR3xp33_ASAP7_75t_L g1083 ( 
.A(n_1067),
.B(n_110),
.C(n_112),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1078),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1077),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1079),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1080),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_1080),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_1082),
.B(n_113),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1081),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_1083),
.A2(n_1075),
.B1(n_1076),
.B2(n_347),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1078),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1078),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1078),
.A2(n_114),
.B1(n_117),
.B2(n_118),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1078),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1084),
.Y(n_1096)
);

AOI21xp33_ASAP7_75t_L g1097 ( 
.A1(n_1093),
.A2(n_196),
.B(n_125),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_SL g1098 ( 
.A1(n_1092),
.A2(n_123),
.B1(n_126),
.B2(n_127),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1088),
.Y(n_1099)
);

AOI222xp33_ASAP7_75t_L g1100 ( 
.A1(n_1086),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.C1(n_133),
.C2(n_134),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1088),
.B(n_135),
.Y(n_1101)
);

NAND3xp33_ASAP7_75t_L g1102 ( 
.A(n_1091),
.B(n_137),
.C(n_138),
.Y(n_1102)
);

XNOR2x1_ASAP7_75t_L g1103 ( 
.A(n_1085),
.B(n_139),
.Y(n_1103)
);

BUFx2_ASAP7_75t_SL g1104 ( 
.A(n_1099),
.Y(n_1104)
);

OAI221xp5_ASAP7_75t_L g1105 ( 
.A1(n_1096),
.A2(n_1087),
.B1(n_1089),
.B2(n_1090),
.C(n_1094),
.Y(n_1105)
);

XNOR2xp5_ASAP7_75t_L g1106 ( 
.A(n_1103),
.B(n_1095),
.Y(n_1106)
);

AOI221xp5_ASAP7_75t_L g1107 ( 
.A1(n_1102),
.A2(n_140),
.B1(n_141),
.B2(n_145),
.C(n_146),
.Y(n_1107)
);

AOI211xp5_ASAP7_75t_L g1108 ( 
.A1(n_1101),
.A2(n_147),
.B(n_149),
.C(n_150),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_1097),
.B(n_151),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1104),
.A2(n_1098),
.B1(n_1100),
.B2(n_158),
.Y(n_1110)
);

OR5x1_ASAP7_75t_L g1111 ( 
.A(n_1105),
.B(n_154),
.C(n_155),
.D(n_159),
.E(n_160),
.Y(n_1111)
);

XNOR2x1_ASAP7_75t_L g1112 ( 
.A(n_1106),
.B(n_161),
.Y(n_1112)
);

NAND3xp33_ASAP7_75t_SL g1113 ( 
.A(n_1110),
.B(n_1109),
.C(n_1108),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1113),
.A2(n_1112),
.B(n_1107),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1114),
.A2(n_1111),
.B(n_166),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1114),
.B(n_164),
.Y(n_1116)
);

OAI222xp33_ASAP7_75t_L g1117 ( 
.A1(n_1116),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.C1(n_170),
.C2(n_171),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1115),
.Y(n_1118)
);

XOR2xp5_ASAP7_75t_L g1119 ( 
.A(n_1116),
.B(n_172),
.Y(n_1119)
);

AO221x2_ASAP7_75t_L g1120 ( 
.A1(n_1118),
.A2(n_1119),
.B1(n_1117),
.B2(n_175),
.C(n_176),
.Y(n_1120)
);

OAI21xp33_ASAP7_75t_L g1121 ( 
.A1(n_1118),
.A2(n_173),
.B(n_174),
.Y(n_1121)
);

AOI221xp5_ASAP7_75t_L g1122 ( 
.A1(n_1121),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.C(n_180),
.Y(n_1122)
);

AOI211xp5_ASAP7_75t_L g1123 ( 
.A1(n_1122),
.A2(n_1120),
.B(n_182),
.C(n_185),
.Y(n_1123)
);


endmodule