module fake_jpeg_9555_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_38),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_24),
.B(n_34),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_47),
.B1(n_17),
.B2(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_54),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_19),
.B1(n_31),
.B2(n_21),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_70),
.B1(n_29),
.B2(n_18),
.Y(n_73)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_58),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_44),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_19),
.B1(n_31),
.B2(n_21),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_68),
.B1(n_29),
.B2(n_18),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_19),
.B1(n_31),
.B2(n_21),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_19),
.B1(n_31),
.B2(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NAND2xp67_ASAP7_75t_SL g110 ( 
.A(n_72),
.B(n_38),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_73),
.A2(n_79),
.B1(n_82),
.B2(n_32),
.Y(n_121)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_94),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_70),
.B1(n_52),
.B2(n_62),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_33),
.B1(n_17),
.B2(n_25),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_85),
.B1(n_93),
.B2(n_34),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_33),
.B1(n_17),
.B2(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_87),
.Y(n_117)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_25),
.B1(n_28),
.B2(n_34),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_42),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_66),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_29),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_100),
.C(n_32),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_28),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_18),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_77),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_103),
.B(n_113),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_107),
.A2(n_22),
.B1(n_30),
.B2(n_12),
.Y(n_157)
);

XNOR2x1_ASAP7_75t_SL g108 ( 
.A(n_72),
.B(n_38),
.Y(n_108)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_122),
.C(n_16),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_109),
.B(n_127),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_110),
.B(n_130),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_91),
.Y(n_113)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_43),
.C(n_38),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_82),
.C(n_74),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_119),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_81),
.B1(n_84),
.B2(n_102),
.Y(n_148)
);

XNOR2x1_ASAP7_75t_SL g122 ( 
.A(n_78),
.B(n_14),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_131),
.Y(n_143)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_79),
.A2(n_28),
.B1(n_32),
.B2(n_30),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_129),
.A2(n_23),
.B(n_128),
.Y(n_163)
);

NOR2x1_ASAP7_75t_L g130 ( 
.A(n_73),
.B(n_22),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_65),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_97),
.B(n_96),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_105),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_144),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_88),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_139),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_87),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_92),
.B1(n_86),
.B2(n_76),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_140),
.A2(n_153),
.B(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_152),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_43),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_105),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_157),
.B1(n_106),
.B2(n_125),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_80),
.Y(n_149)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_101),
.B1(n_84),
.B2(n_81),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_151),
.B1(n_117),
.B2(n_104),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_86),
.B1(n_80),
.B2(n_67),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

NAND2x1_ASAP7_75t_SL g153 ( 
.A(n_115),
.B(n_20),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_0),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_0),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_155),
.A2(n_163),
.B(n_23),
.Y(n_192)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_161),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_43),
.Y(n_158)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_160),
.B(n_0),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_16),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_171),
.B1(n_180),
.B2(n_183),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_166),
.A2(n_192),
.B(n_156),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_111),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_168),
.B(n_178),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_111),
.B1(n_125),
.B2(n_120),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_147),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_179),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_175),
.A2(n_177),
.B1(n_194),
.B2(n_145),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_114),
.Y(n_176)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_161),
.A2(n_117),
.B1(n_124),
.B2(n_71),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_162),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_120),
.B1(n_69),
.B2(n_20),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_134),
.B(n_16),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_195),
.C(n_145),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_159),
.A2(n_20),
.B1(n_75),
.B2(n_123),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_162),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_188),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_75),
.B1(n_23),
.B2(n_15),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_189),
.A2(n_144),
.B1(n_137),
.B2(n_147),
.Y(n_224)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_23),
.A3(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_191)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_138),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_193),
.B(n_196),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_132),
.A2(n_75),
.B1(n_23),
.B2(n_2),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_142),
.B(n_23),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_151),
.Y(n_196)
);

A2O1A1O1Ixp25_ASAP7_75t_L g202 ( 
.A1(n_197),
.A2(n_192),
.B(n_168),
.C(n_185),
.D(n_191),
.Y(n_202)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_203),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_197),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_169),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_204),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_205),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_218),
.C(n_222),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_210),
.B(n_221),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_185),
.A2(n_153),
.B(n_140),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_219),
.Y(n_248)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_225),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_216),
.A2(n_224),
.B1(n_174),
.B2(n_181),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_175),
.A2(n_136),
.B1(n_133),
.B2(n_148),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_217),
.A2(n_174),
.B1(n_180),
.B2(n_183),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_133),
.C(n_153),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_190),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_165),
.B(n_152),
.Y(n_220)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_176),
.B(n_155),
.Y(n_221)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_170),
.B(n_150),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_173),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_223),
.B(n_12),
.Y(n_244)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_170),
.B(n_195),
.C(n_182),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_194),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_247),
.C(n_206),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_217),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_230),
.B(n_234),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_177),
.B1(n_166),
.B2(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_231),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_200),
.A2(n_219),
.B1(n_214),
.B2(n_225),
.Y(n_232)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_233),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_208),
.B(n_155),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_208),
.B(n_154),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_237),
.B(n_239),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_167),
.B1(n_154),
.B2(n_3),
.Y(n_238)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_201),
.A2(n_13),
.B(n_12),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_207),
.Y(n_258)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_11),
.C(n_10),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_245),
.B(n_251),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_199),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_246)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_10),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_199),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_246),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_4),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_252),
.B(n_204),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

FAx1_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_216),
.CI(n_210),
.CON(n_254),
.SN(n_254)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_254),
.A2(n_250),
.B(n_243),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_227),
.Y(n_256)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_259),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_222),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_272),
.Y(n_285)
);

INVxp33_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_266),
.B(n_270),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_218),
.C(n_215),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_259),
.C(n_261),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_209),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_228),
.B(n_202),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_273),
.A2(n_240),
.B(n_241),
.Y(n_274)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_277),
.C(n_278),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_230),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_250),
.C(n_243),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_231),
.Y(n_279)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_256),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_198),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_284),
.A2(n_271),
.B(n_257),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_242),
.B(n_213),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_286),
.A2(n_289),
.B(n_239),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_258),
.B(n_237),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_290),
.C(n_268),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_264),
.A2(n_242),
.B(n_229),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_234),
.Y(n_290)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_292),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_263),
.B1(n_267),
.B2(n_254),
.Y(n_293)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

AOI22x1_ASAP7_75t_SL g295 ( 
.A1(n_284),
.A2(n_254),
.B1(n_268),
.B2(n_260),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_282),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_281),
.A2(n_266),
.B1(n_256),
.B2(n_249),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_301),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_304),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_287),
.A2(n_283),
.B1(n_288),
.B2(n_279),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_300),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_290),
.B(n_285),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_286),
.A2(n_255),
.B1(n_265),
.B2(n_247),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_275),
.B(n_205),
.C(n_5),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_305),
.C(n_6),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_278),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_6),
.C(n_7),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_295),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_307),
.Y(n_323)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

OAI21xp33_ASAP7_75t_L g326 ( 
.A1(n_308),
.A2(n_314),
.B(n_7),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_294),
.A2(n_285),
.B(n_277),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_291),
.B(n_303),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_7),
.C(n_8),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_298),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_305),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_318),
.B(n_322),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_321),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_309),
.A2(n_291),
.B(n_302),
.Y(n_320)
);

AOI211xp5_ASAP7_75t_L g327 ( 
.A1(n_320),
.A2(n_314),
.B(n_313),
.C(n_308),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_315),
.A2(n_300),
.B1(n_8),
.B2(n_9),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_325),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_7),
.Y(n_325)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_326),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_327),
.Y(n_333)
);

OAI21x1_ASAP7_75t_SL g332 ( 
.A1(n_326),
.A2(n_323),
.B(n_307),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_316),
.Y(n_335)
);

A2O1A1O1Ixp25_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_331),
.B(n_328),
.C(n_329),
.D(n_321),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_333),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_334),
.B(n_330),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_339),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_8),
.Y(n_341)
);


endmodule