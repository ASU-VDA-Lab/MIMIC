module fake_netlist_6_2231_n_804 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_804);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_804;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_698;
wire n_617;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_758;
wire n_525;
wire n_720;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_796;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_683;
wire n_420;
wire n_620;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVxp67_ASAP7_75t_L g166 ( 
.A(n_11),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_89),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_28),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_104),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_82),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_4),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_22),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_39),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_35),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_49),
.Y(n_177)
);

NOR2xp67_ASAP7_75t_L g178 ( 
.A(n_2),
.B(n_106),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_101),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_58),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_46),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_59),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_25),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_9),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_85),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_76),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_8),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_43),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_70),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_153),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_81),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_134),
.Y(n_197)
);

NOR2xp67_ASAP7_75t_L g198 ( 
.A(n_142),
.B(n_116),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_114),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_8),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_20),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_74),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_140),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_55),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_150),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_11),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_37),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_127),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_159),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_112),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_24),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_47),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_4),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_111),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_75),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_109),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_149),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_115),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_56),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_51),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_110),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_97),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_30),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_67),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_69),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_14),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_53),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_118),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_125),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_175),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_169),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_200),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_183),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_196),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_196),
.B(n_3),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_175),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

OA21x2_ASAP7_75t_L g249 ( 
.A1(n_214),
.A2(n_5),
.B(n_6),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_215),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_169),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_194),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_194),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_215),
.Y(n_255)
);

OAI21x1_ASAP7_75t_L g256 ( 
.A1(n_217),
.A2(n_7),
.B(n_9),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g258 ( 
.A(n_168),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_217),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_194),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_194),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_200),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_227),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_178),
.Y(n_265)
);

AND2x4_ASAP7_75t_L g266 ( 
.A(n_167),
.B(n_23),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_176),
.A2(n_210),
.B1(n_203),
.B2(n_216),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_L g268 ( 
.A(n_176),
.B(n_180),
.C(n_174),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_181),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_184),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_187),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_189),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_203),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_190),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_192),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_193),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_230),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_204),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_240),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_267),
.B(n_216),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_260),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_195),
.Y(n_285)
);

NAND3xp33_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_229),
.C(n_170),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_209),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_261),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_205),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_244),
.B(n_212),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_230),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_230),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_230),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_230),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_270),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_234),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_240),
.A2(n_211),
.B1(n_198),
.B2(n_224),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_231),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_234),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_231),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g303 ( 
.A1(n_242),
.A2(n_228),
.B(n_225),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_231),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_258),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_273),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_231),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_252),
.Y(n_308)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_241),
.A2(n_219),
.B(n_221),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_263),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_231),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_262),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_236),
.Y(n_313)
);

NAND2xp33_ASAP7_75t_L g314 ( 
.A(n_251),
.B(n_171),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_263),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_236),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_L g318 ( 
.A1(n_233),
.A2(n_220),
.B1(n_222),
.B2(n_218),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_252),
.B(n_172),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_257),
.A2(n_208),
.B1(n_207),
.B2(n_202),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_236),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_236),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_245),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_245),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_232),
.A2(n_199),
.B1(n_197),
.B2(n_188),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_245),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_245),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_253),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_285),
.B(n_290),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_280),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_280),
.B(n_266),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_316),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_280),
.Y(n_334)
);

O2A1O1Ixp5_ASAP7_75t_L g335 ( 
.A1(n_303),
.A2(n_309),
.B(n_281),
.C(n_276),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_266),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_304),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_237),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_325),
.B(n_266),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_307),
.B(n_247),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_303),
.A2(n_256),
.B(n_249),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_316),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_314),
.A2(n_249),
.B1(n_256),
.B2(n_272),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_314),
.A2(n_258),
.B1(n_237),
.B2(n_246),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_321),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_282),
.B(n_177),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_322),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_299),
.B(n_247),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_322),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_327),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_307),
.B(n_247),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_328),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_328),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_282),
.B(n_246),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_328),
.B(n_272),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_327),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_318),
.A2(n_179),
.B1(n_182),
.B2(n_249),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_292),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_289),
.B(n_269),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_329),
.B(n_269),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_305),
.B(n_273),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_308),
.B(n_275),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_269),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_308),
.B(n_271),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_292),
.B(n_271),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_296),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_293),
.B(n_275),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_319),
.A2(n_249),
.B1(n_235),
.B2(n_239),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_293),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_286),
.B(n_253),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_306),
.B(n_262),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_294),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_294),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_298),
.B(n_235),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_295),
.B(n_300),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_295),
.B(n_300),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_287),
.B(n_241),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_R g380 ( 
.A(n_305),
.B(n_26),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_283),
.A2(n_259),
.B1(n_264),
.B2(n_255),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_302),
.B(n_311),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_309),
.B(n_253),
.Y(n_383)
);

AOI221xp5_ASAP7_75t_L g384 ( 
.A1(n_312),
.A2(n_239),
.B1(n_259),
.B2(n_255),
.C(n_250),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_297),
.B(n_253),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_304),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_302),
.B(n_253),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_311),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_323),
.B(n_324),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_297),
.B(n_248),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_288),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_323),
.B(n_248),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_301),
.B(n_250),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_301),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_310),
.Y(n_395)
);

A2O1A1Ixp33_ASAP7_75t_L g396 ( 
.A1(n_310),
.A2(n_264),
.B(n_238),
.C(n_13),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_313),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_332),
.A2(n_313),
.B(n_317),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_330),
.B(n_315),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_349),
.A2(n_315),
.B1(n_288),
.B2(n_291),
.Y(n_400)
);

O2A1O1Ixp33_ASAP7_75t_L g401 ( 
.A1(n_361),
.A2(n_291),
.B(n_278),
.C(n_279),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_313),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_373),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_355),
.B(n_356),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_347),
.B(n_10),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_366),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_347),
.B(n_10),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_380),
.Y(n_408)
);

INVx6_ASAP7_75t_SL g409 ( 
.A(n_363),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_349),
.B(n_356),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_370),
.B(n_324),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_339),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_336),
.A2(n_317),
.B(n_326),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_379),
.B(n_277),
.Y(n_414)
);

A2O1A1Ixp33_ASAP7_75t_L g415 ( 
.A1(n_341),
.A2(n_284),
.B(n_279),
.C(n_278),
.Y(n_415)
);

INVx3_ASAP7_75t_SL g416 ( 
.A(n_339),
.Y(n_416)
);

BUFx12f_ASAP7_75t_L g417 ( 
.A(n_394),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_335),
.A2(n_344),
.B(n_383),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_395),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_340),
.A2(n_352),
.B(n_377),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_344),
.A2(n_284),
.B(n_277),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_381),
.B(n_364),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_378),
.A2(n_317),
.B(n_326),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_376),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_379),
.B(n_304),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_382),
.A2(n_389),
.B(n_383),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_372),
.A2(n_317),
.B(n_326),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_372),
.A2(n_317),
.B(n_326),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_381),
.B(n_304),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_359),
.A2(n_326),
.B(n_304),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_357),
.A2(n_90),
.B(n_163),
.Y(n_432)
);

NOR3xp33_ASAP7_75t_L g433 ( 
.A(n_338),
.B(n_396),
.C(n_384),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_364),
.B(n_12),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_368),
.B(n_12),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_333),
.B(n_27),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_342),
.A2(n_91),
.B(n_162),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_L g438 ( 
.A1(n_343),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_338),
.Y(n_439)
);

INVx11_ASAP7_75t_L g440 ( 
.A(n_380),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_346),
.B(n_29),
.Y(n_441)
);

NOR2xp67_ASAP7_75t_L g442 ( 
.A(n_345),
.B(n_164),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_367),
.A2(n_93),
.B(n_160),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_369),
.A2(n_365),
.B(n_362),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_360),
.Y(n_445)
);

O2A1O1Ixp33_ASAP7_75t_L g446 ( 
.A1(n_393),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_446)
);

BUFx4f_ASAP7_75t_L g447 ( 
.A(n_390),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_393),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_397),
.B(n_18),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_392),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_397),
.A2(n_95),
.B(n_158),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_348),
.B(n_350),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_351),
.B(n_31),
.Y(n_453)
);

INVx11_ASAP7_75t_L g454 ( 
.A(n_385),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_387),
.A2(n_94),
.B(n_157),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_331),
.A2(n_88),
.B(n_156),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_358),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_371),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_374),
.B(n_32),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_334),
.A2(n_96),
.B(n_155),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_353),
.A2(n_87),
.B(n_154),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_375),
.B(n_33),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_354),
.B(n_19),
.Y(n_463)
);

AOI21x1_ASAP7_75t_L g464 ( 
.A1(n_388),
.A2(n_98),
.B(n_34),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_337),
.B(n_99),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_337),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_385),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_424),
.Y(n_468)
);

OAI21x1_ASAP7_75t_L g469 ( 
.A1(n_427),
.A2(n_386),
.B(n_337),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_452),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_447),
.B(n_337),
.Y(n_471)
);

AOI21x1_ASAP7_75t_L g472 ( 
.A1(n_411),
.A2(n_386),
.B(n_36),
.Y(n_472)
);

AO31x2_ASAP7_75t_L g473 ( 
.A1(n_415),
.A2(n_405),
.A3(n_407),
.B(n_449),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_452),
.Y(n_474)
);

A2O1A1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_410),
.A2(n_386),
.B(n_21),
.C(n_40),
.Y(n_475)
);

O2A1O1Ixp5_ASAP7_75t_L g476 ( 
.A1(n_431),
.A2(n_386),
.B(n_41),
.C(n_42),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_447),
.B(n_404),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_399),
.B(n_38),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_406),
.B(n_44),
.Y(n_479)
);

OAI21x1_ASAP7_75t_L g480 ( 
.A1(n_420),
.A2(n_161),
.B(n_48),
.Y(n_480)
);

AO31x2_ASAP7_75t_L g481 ( 
.A1(n_448),
.A2(n_45),
.A3(n_50),
.B(n_52),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_450),
.B(n_412),
.Y(n_482)
);

CKINVDCx6p67_ASAP7_75t_R g483 ( 
.A(n_417),
.Y(n_483)
);

OAI21xp33_ASAP7_75t_L g484 ( 
.A1(n_433),
.A2(n_54),
.B(n_57),
.Y(n_484)
);

AOI221x1_ASAP7_75t_L g485 ( 
.A1(n_431),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.C(n_63),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_422),
.B(n_64),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_418),
.A2(n_65),
.B(n_66),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_425),
.B(n_68),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_444),
.A2(n_421),
.B(n_398),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_418),
.A2(n_71),
.B(n_72),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_419),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_419),
.B(n_73),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_445),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_402),
.B(n_77),
.Y(n_494)
);

AOI211x1_ASAP7_75t_L g495 ( 
.A1(n_437),
.A2(n_78),
.B(n_79),
.C(n_80),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_421),
.A2(n_83),
.B(n_84),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_413),
.A2(n_152),
.B(n_100),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_414),
.B(n_86),
.Y(n_498)
);

AO21x2_ASAP7_75t_L g499 ( 
.A1(n_437),
.A2(n_102),
.B(n_103),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_403),
.B(n_105),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_430),
.A2(n_107),
.B(n_108),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_409),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_458),
.Y(n_503)
);

NOR2x1_ASAP7_75t_SL g504 ( 
.A(n_465),
.B(n_117),
.Y(n_504)
);

AOI221xp5_ASAP7_75t_SL g505 ( 
.A1(n_448),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.C(n_123),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_428),
.A2(n_126),
.B(n_128),
.Y(n_506)
);

AOI21xp33_ASAP7_75t_L g507 ( 
.A1(n_446),
.A2(n_129),
.B(n_130),
.Y(n_507)
);

OAI21xp33_ASAP7_75t_L g508 ( 
.A1(n_439),
.A2(n_131),
.B(n_132),
.Y(n_508)
);

OAI21x1_ASAP7_75t_SL g509 ( 
.A1(n_464),
.A2(n_133),
.B(n_135),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_467),
.B(n_434),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_408),
.B(n_136),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_466),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_426),
.A2(n_137),
.B(n_138),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_400),
.A2(n_141),
.B(n_144),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_466),
.A2(n_441),
.B(n_436),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_416),
.B(n_145),
.Y(n_516)
);

AOI221xp5_ASAP7_75t_L g517 ( 
.A1(n_457),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.C(n_151),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_435),
.B(n_453),
.Y(n_518)
);

OAI21xp33_ASAP7_75t_SL g519 ( 
.A1(n_454),
.A2(n_438),
.B(n_440),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_451),
.B(n_463),
.Y(n_520)
);

AO21x2_ASAP7_75t_L g521 ( 
.A1(n_459),
.A2(n_462),
.B(n_429),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_401),
.A2(n_423),
.B(n_432),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_486),
.A2(n_443),
.B(n_455),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_482),
.B(n_442),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_469),
.A2(n_472),
.B(n_489),
.Y(n_525)
);

O2A1O1Ixp33_ASAP7_75t_SL g526 ( 
.A1(n_475),
.A2(n_457),
.B(n_456),
.C(n_460),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_510),
.B(n_409),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_476),
.A2(n_461),
.B(n_478),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_468),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_474),
.B(n_477),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_518),
.A2(n_494),
.B(n_515),
.Y(n_531)
);

OA21x2_ASAP7_75t_L g532 ( 
.A1(n_485),
.A2(n_505),
.B(n_522),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_470),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_488),
.B(n_491),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_503),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_480),
.A2(n_522),
.B(n_497),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_491),
.B(n_479),
.Y(n_537)
);

AOI221xp5_ASAP7_75t_L g538 ( 
.A1(n_507),
.A2(n_495),
.B1(n_519),
.B2(n_514),
.C(n_517),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_493),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_491),
.B(n_512),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_506),
.A2(n_509),
.B(n_492),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_502),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_496),
.A2(n_520),
.B(n_490),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_500),
.Y(n_544)
);

OR2x6_ASAP7_75t_L g545 ( 
.A(n_516),
.B(n_514),
.Y(n_545)
);

CKINVDCx11_ASAP7_75t_R g546 ( 
.A(n_483),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_512),
.Y(n_547)
);

AOI21x1_ASAP7_75t_L g548 ( 
.A1(n_498),
.A2(n_471),
.B(n_513),
.Y(n_548)
);

OA21x2_ASAP7_75t_L g549 ( 
.A1(n_505),
.A2(n_487),
.B(n_490),
.Y(n_549)
);

OAI21x1_ASAP7_75t_L g550 ( 
.A1(n_520),
.A2(n_501),
.B(n_487),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_501),
.A2(n_484),
.B(n_508),
.Y(n_551)
);

NOR2x1_ASAP7_75t_SL g552 ( 
.A(n_499),
.B(n_521),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_SL g553 ( 
.A1(n_499),
.A2(n_511),
.B1(n_504),
.B2(n_507),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_473),
.B(n_481),
.Y(n_554)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_521),
.A2(n_473),
.B(n_481),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_481),
.Y(n_556)
);

NAND2x1p5_ASAP7_75t_L g557 ( 
.A(n_473),
.B(n_491),
.Y(n_557)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_469),
.A2(n_472),
.B(n_489),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_491),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_L g560 ( 
.A1(n_486),
.A2(n_410),
.B(n_418),
.Y(n_560)
);

AOI221xp5_ASAP7_75t_L g561 ( 
.A1(n_507),
.A2(n_410),
.B1(n_318),
.B2(n_283),
.C(n_439),
.Y(n_561)
);

OAI21x1_ASAP7_75t_L g562 ( 
.A1(n_469),
.A2(n_472),
.B(n_489),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_510),
.B(n_355),
.Y(n_563)
);

OAI21x1_ASAP7_75t_L g564 ( 
.A1(n_469),
.A2(n_472),
.B(n_489),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_468),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_468),
.Y(n_566)
);

OAI21x1_ASAP7_75t_L g567 ( 
.A1(n_469),
.A2(n_472),
.B(n_489),
.Y(n_567)
);

AO21x2_ASAP7_75t_L g568 ( 
.A1(n_552),
.A2(n_554),
.B(n_536),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_547),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_547),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_557),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_540),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_557),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_525),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_529),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_563),
.B(n_534),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_533),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_525),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_546),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_540),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_558),
.Y(n_581)
);

CKINVDCx6p67_ASAP7_75t_R g582 ( 
.A(n_546),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_527),
.B(n_561),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_558),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_565),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_533),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_566),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_535),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_559),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_539),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_542),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_555),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_562),
.Y(n_593)
);

AO21x1_ASAP7_75t_L g594 ( 
.A1(n_560),
.A2(n_551),
.B(n_550),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_562),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_544),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_555),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_556),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_540),
.B(n_538),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_559),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_564),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_556),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_530),
.Y(n_603)
);

OA21x2_ASAP7_75t_L g604 ( 
.A1(n_567),
.A2(n_543),
.B(n_551),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_556),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_545),
.B(n_549),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_556),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_537),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_574),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_574),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_574),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_583),
.B(n_545),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_583),
.B(n_545),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_598),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_576),
.A2(n_524),
.B1(n_553),
.B2(n_530),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_599),
.B(n_549),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_598),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_599),
.B(n_549),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_608),
.B(n_532),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_608),
.B(n_532),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_602),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_602),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_586),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_576),
.B(n_532),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_569),
.B(n_530),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_605),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_605),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_586),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_607),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_596),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_578),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_577),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_606),
.B(n_543),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_589),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_591),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_606),
.B(n_553),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_572),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_569),
.B(n_528),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_607),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_603),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_570),
.B(n_548),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_571),
.B(n_541),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_592),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_570),
.B(n_585),
.Y(n_644)
);

NOR2x1p5_ASAP7_75t_L g645 ( 
.A(n_582),
.B(n_526),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_600),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_575),
.B(n_531),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_575),
.B(n_526),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_572),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_592),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_580),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_585),
.B(n_523),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_580),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_587),
.B(n_588),
.Y(n_654)
);

INVxp67_ASAP7_75t_SL g655 ( 
.A(n_628),
.Y(n_655)
);

NAND2x1p5_ASAP7_75t_L g656 ( 
.A(n_632),
.B(n_573),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_642),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_654),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_630),
.B(n_590),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_635),
.B(n_590),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_612),
.B(n_588),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_623),
.B(n_587),
.Y(n_662)
);

NAND3xp33_ASAP7_75t_L g663 ( 
.A(n_615),
.B(n_573),
.C(n_571),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_625),
.B(n_571),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_654),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_623),
.B(n_594),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_612),
.B(n_594),
.Y(n_667)
);

NAND4xp25_ASAP7_75t_L g668 ( 
.A(n_632),
.B(n_597),
.C(n_584),
.D(n_581),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_643),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_613),
.B(n_604),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_643),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_650),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_609),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_609),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_613),
.B(n_582),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_645),
.A2(n_640),
.B1(n_652),
.B2(n_647),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_644),
.B(n_604),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_640),
.B(n_604),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_625),
.B(n_601),
.Y(n_679)
);

INVxp67_ASAP7_75t_SL g680 ( 
.A(n_646),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_642),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_650),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_624),
.B(n_604),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_637),
.B(n_601),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_610),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_610),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_624),
.B(n_597),
.Y(n_687)
);

NAND4xp25_ASAP7_75t_L g688 ( 
.A(n_634),
.B(n_584),
.C(n_593),
.D(n_595),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_644),
.B(n_645),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_636),
.B(n_568),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_634),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_611),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_669),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_667),
.B(n_636),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_680),
.B(n_661),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_670),
.B(n_618),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_690),
.B(n_633),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_671),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_655),
.B(n_652),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_683),
.B(n_618),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_679),
.B(n_633),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_657),
.B(n_616),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_672),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_682),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_678),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_659),
.B(n_616),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_657),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_660),
.B(n_647),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_691),
.B(n_638),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_673),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_681),
.Y(n_711)
);

AND2x2_ASAP7_75t_SL g712 ( 
.A(n_676),
.B(n_648),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_662),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_681),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_666),
.B(n_631),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_673),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_664),
.B(n_638),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_683),
.B(n_620),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_685),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_679),
.B(n_620),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_664),
.B(n_619),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_674),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_693),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_705),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_693),
.Y(n_725)
);

NOR2x1_ASAP7_75t_L g726 ( 
.A(n_699),
.B(n_668),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_697),
.B(n_677),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_713),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_708),
.B(n_676),
.C(n_663),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_697),
.B(n_687),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_703),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_703),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_698),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_704),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_709),
.B(n_664),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_707),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_700),
.B(n_679),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_694),
.B(n_675),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_695),
.B(n_706),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_718),
.B(n_685),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_712),
.A2(n_675),
.B1(n_688),
.B2(n_689),
.Y(n_741)
);

INVx1_ASAP7_75t_SL g742 ( 
.A(n_724),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_739),
.B(n_694),
.Y(n_743)
);

OAI221xp5_ASAP7_75t_L g744 ( 
.A1(n_741),
.A2(n_656),
.B1(n_717),
.B2(n_714),
.C(n_711),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_724),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_741),
.A2(n_712),
.B1(n_656),
.B2(n_721),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_738),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_723),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_728),
.B(n_696),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_L g750 ( 
.A(n_726),
.B(n_579),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_728),
.B(n_696),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_733),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_748),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_742),
.Y(n_754)
);

AOI322xp5_ASAP7_75t_L g755 ( 
.A1(n_750),
.A2(n_700),
.A3(n_718),
.B1(n_734),
.B2(n_729),
.C1(n_731),
.C2(n_725),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_743),
.B(n_737),
.Y(n_756)
);

XOR2x2_ASAP7_75t_L g757 ( 
.A(n_746),
.B(n_735),
.Y(n_757)
);

XNOR2x1_ASAP7_75t_L g758 ( 
.A(n_742),
.B(n_737),
.Y(n_758)
);

NOR3xp33_ASAP7_75t_L g759 ( 
.A(n_754),
.B(n_744),
.C(n_753),
.Y(n_759)
);

AOI221x1_ASAP7_75t_L g760 ( 
.A1(n_756),
.A2(n_745),
.B1(n_736),
.B2(n_752),
.C(n_751),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_755),
.B(n_747),
.Y(n_761)
);

NAND4xp25_ASAP7_75t_L g762 ( 
.A(n_755),
.B(n_749),
.C(n_727),
.D(n_732),
.Y(n_762)
);

OAI21xp33_ASAP7_75t_SL g763 ( 
.A1(n_758),
.A2(n_730),
.B(n_740),
.Y(n_763)
);

OAI211xp5_ASAP7_75t_SL g764 ( 
.A1(n_757),
.A2(n_715),
.B(n_719),
.C(n_665),
.Y(n_764)
);

AOI211xp5_ASAP7_75t_SL g765 ( 
.A1(n_761),
.A2(n_715),
.B(n_719),
.C(n_622),
.Y(n_765)
);

OAI21xp33_ASAP7_75t_L g766 ( 
.A1(n_763),
.A2(n_701),
.B(n_702),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_759),
.B(n_701),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_760),
.B(n_701),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_762),
.Y(n_769)
);

NOR2x1_ASAP7_75t_L g770 ( 
.A(n_769),
.B(n_764),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_765),
.B(n_658),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_766),
.B(n_702),
.Y(n_772)
);

NOR2x1_ASAP7_75t_L g773 ( 
.A(n_770),
.B(n_768),
.Y(n_773)
);

NAND3x1_ASAP7_75t_L g774 ( 
.A(n_771),
.B(n_767),
.C(n_648),
.Y(n_774)
);

NOR4xp75_ASAP7_75t_L g775 ( 
.A(n_772),
.B(n_651),
.C(n_649),
.D(n_720),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_774),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_773),
.B(n_720),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_775),
.A2(n_637),
.B1(n_653),
.B2(n_684),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_773),
.B(n_722),
.Y(n_779)
);

OAI211xp5_ASAP7_75t_L g780 ( 
.A1(n_773),
.A2(n_627),
.B(n_621),
.C(n_626),
.Y(n_780)
);

OA22x2_ASAP7_75t_L g781 ( 
.A1(n_776),
.A2(n_629),
.B1(n_622),
.B2(n_621),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_777),
.A2(n_780),
.B1(n_779),
.B2(n_778),
.Y(n_782)
);

NAND4xp25_ASAP7_75t_SL g783 ( 
.A(n_777),
.B(n_639),
.C(n_629),
.D(n_627),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_SL g784 ( 
.A1(n_776),
.A2(n_651),
.B1(n_649),
.B2(n_637),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_777),
.A2(n_626),
.B1(n_639),
.B2(n_617),
.Y(n_785)
);

AND3x2_ASAP7_75t_L g786 ( 
.A(n_779),
.B(n_617),
.C(n_614),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_777),
.Y(n_787)
);

INVx1_ASAP7_75t_SL g788 ( 
.A(n_787),
.Y(n_788)
);

XOR2xp5_ASAP7_75t_L g789 ( 
.A(n_782),
.B(n_653),
.Y(n_789)
);

XNOR2xp5_ASAP7_75t_L g790 ( 
.A(n_784),
.B(n_653),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_781),
.Y(n_791)
);

AND3x1_ASAP7_75t_L g792 ( 
.A(n_783),
.B(n_614),
.C(n_722),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_788),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_791),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_789),
.A2(n_785),
.B1(n_786),
.B2(n_684),
.Y(n_795)
);

AOI21x1_ASAP7_75t_L g796 ( 
.A1(n_790),
.A2(n_716),
.B(n_710),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_794),
.B(n_792),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_793),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_795),
.B(n_716),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_796),
.A2(n_641),
.B(n_710),
.Y(n_800)
);

OA22x2_ASAP7_75t_L g801 ( 
.A1(n_798),
.A2(n_684),
.B1(n_619),
.B2(n_641),
.Y(n_801)
);

OA21x2_ASAP7_75t_L g802 ( 
.A1(n_801),
.A2(n_797),
.B(n_799),
.Y(n_802)
);

AO21x2_ASAP7_75t_L g803 ( 
.A1(n_802),
.A2(n_800),
.B(n_692),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_803),
.A2(n_686),
.B(n_674),
.Y(n_804)
);


endmodule