module fake_netlist_1_5233_n_548 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_548);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_548;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_14), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_6), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_14), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_1), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_77), .Y(n_83) );
BUFx6f_ASAP7_75t_L g84 ( .A(n_6), .Y(n_84) );
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_12), .Y(n_85) );
INVxp67_ASAP7_75t_L g86 ( .A(n_64), .Y(n_86) );
CKINVDCx16_ASAP7_75t_R g87 ( .A(n_22), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_70), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_52), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_32), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_76), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_31), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_30), .Y(n_93) );
HB1xp67_ASAP7_75t_L g94 ( .A(n_74), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_73), .Y(n_95) );
INVx3_ASAP7_75t_L g96 ( .A(n_16), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_71), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_39), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_57), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_49), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_35), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_50), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_20), .Y(n_103) );
INVxp33_ASAP7_75t_L g104 ( .A(n_67), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_38), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_51), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_54), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_29), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_41), .Y(n_109) );
NOR2xp67_ASAP7_75t_L g110 ( .A(n_63), .B(n_8), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_78), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_13), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_55), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_59), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_33), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_65), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_89), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_89), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_94), .B(n_0), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_93), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_96), .Y(n_121) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_88), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_104), .B(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_96), .Y(n_124) );
NAND2xp33_ASAP7_75t_L g125 ( .A(n_88), .B(n_28), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_96), .B(n_1), .Y(n_126) );
BUFx8_ASAP7_75t_L g127 ( .A(n_93), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_79), .B(n_2), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_97), .B(n_98), .Y(n_132) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_81), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_87), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_99), .B(n_101), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_90), .Y(n_136) );
AOI22xp5_ASAP7_75t_L g137 ( .A1(n_85), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_90), .Y(n_138) );
AND2x2_ASAP7_75t_SL g139 ( .A(n_91), .B(n_75), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_129), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_122), .B(n_100), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_128), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_126), .B(n_81), .Y(n_143) );
INVx5_ASAP7_75t_L g144 ( .A(n_117), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_127), .B(n_100), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_136), .B(n_116), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_128), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_136), .B(n_103), .Y(n_148) );
CKINVDCx8_ASAP7_75t_R g149 ( .A(n_134), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_127), .B(n_107), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_127), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_133), .B(n_82), .Y(n_152) );
INVx5_ASAP7_75t_L g153 ( .A(n_117), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_128), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_138), .B(n_107), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_120), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_120), .Y(n_157) );
BUFx8_ASAP7_75t_SL g158 ( .A(n_119), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_120), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_132), .B(n_105), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_138), .B(n_121), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_123), .B(n_106), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_123), .B(n_86), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_135), .B(n_102), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_155), .B(n_127), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_160), .B(n_126), .Y(n_166) );
OR2x2_ASAP7_75t_L g167 ( .A(n_162), .B(n_137), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_163), .B(n_139), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_143), .B(n_139), .Y(n_169) );
INVx2_ASAP7_75t_SL g170 ( .A(n_151), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_142), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_142), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_147), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_143), .A2(n_139), .B1(n_131), .B2(n_130), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_143), .B(n_130), .Y(n_176) );
INVx2_ASAP7_75t_SL g177 ( .A(n_151), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_151), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_143), .B(n_124), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_154), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_154), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_156), .Y(n_182) );
INVxp33_ASAP7_75t_L g183 ( .A(n_158), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_152), .B(n_121), .Y(n_184) );
AO22x1_ASAP7_75t_L g185 ( .A1(n_146), .A2(n_80), .B1(n_111), .B2(n_91), .Y(n_185) );
INVxp67_ASAP7_75t_L g186 ( .A(n_152), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_164), .B(n_124), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_161), .B(n_82), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_146), .B(n_112), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
AND2x6_ASAP7_75t_L g191 ( .A(n_161), .B(n_109), .Y(n_191) );
AOI211xp5_ASAP7_75t_L g192 ( .A1(n_141), .A2(n_137), .B(n_112), .C(n_125), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_157), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_159), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_159), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_153), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_165), .A2(n_145), .B(n_150), .Y(n_198) );
CKINVDCx8_ASAP7_75t_R g199 ( .A(n_191), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_178), .Y(n_200) );
OR2x2_ASAP7_75t_L g201 ( .A(n_167), .B(n_148), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_174), .A2(n_148), .B1(n_92), .B2(n_114), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_169), .A2(n_84), .B1(n_117), .B2(n_118), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_170), .A2(n_114), .B(n_92), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_178), .Y(n_205) );
INVx5_ASAP7_75t_L g206 ( .A(n_178), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_193), .Y(n_207) );
NOR2x1_ASAP7_75t_L g208 ( .A(n_167), .B(n_110), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_168), .A2(n_115), .B1(n_95), .B2(n_108), .Y(n_209) );
BUFx4f_ASAP7_75t_SL g210 ( .A(n_184), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_170), .B(n_149), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_179), .B(n_149), .Y(n_212) );
NAND2x1p5_ASAP7_75t_L g213 ( .A(n_182), .B(n_115), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_179), .B(n_111), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_182), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_186), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_177), .B(n_95), .Y(n_217) );
INVx1_ASAP7_75t_SL g218 ( .A(n_188), .Y(n_218) );
INVxp33_ASAP7_75t_SL g219 ( .A(n_166), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_179), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_190), .Y(n_221) );
BUFx12f_ASAP7_75t_L g222 ( .A(n_189), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_187), .B(n_108), .Y(n_223) );
BUFx2_ASAP7_75t_L g224 ( .A(n_191), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_171), .A2(n_109), .B(n_113), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_176), .A2(n_113), .B1(n_84), .B2(n_118), .Y(n_226) );
AOI22xp33_ASAP7_75t_SL g227 ( .A1(n_189), .A2(n_84), .B1(n_118), .B2(n_117), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_188), .B(n_3), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_190), .Y(n_229) );
OAI21x1_ASAP7_75t_L g230 ( .A1(n_171), .A2(n_140), .B(n_153), .Y(n_230) );
INVx5_ASAP7_75t_L g231 ( .A(n_200), .Y(n_231) );
OAI21x1_ASAP7_75t_L g232 ( .A1(n_230), .A2(n_181), .B(n_175), .Y(n_232) );
CKINVDCx11_ASAP7_75t_R g233 ( .A(n_222), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_215), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_215), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_218), .B(n_189), .Y(n_236) );
OAI21x1_ASAP7_75t_L g237 ( .A1(n_230), .A2(n_175), .B(n_181), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_201), .B(n_193), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_201), .B(n_196), .Y(n_239) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_225), .A2(n_173), .B(n_172), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_206), .Y(n_241) );
INVxp33_ASAP7_75t_L g242 ( .A(n_216), .Y(n_242) );
BUFx4f_ASAP7_75t_SL g243 ( .A(n_222), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_207), .Y(n_244) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_198), .A2(n_173), .B(n_172), .Y(n_245) );
NOR2xp67_ASAP7_75t_L g246 ( .A(n_206), .B(n_196), .Y(n_246) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_213), .A2(n_180), .B(n_195), .Y(n_247) );
OAI21x1_ASAP7_75t_SL g248 ( .A1(n_221), .A2(n_180), .B(n_194), .Y(n_248) );
AOI21x1_ASAP7_75t_L g249 ( .A1(n_208), .A2(n_185), .B(n_140), .Y(n_249) );
INVx6_ASAP7_75t_L g250 ( .A(n_206), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_213), .A2(n_192), .B1(n_177), .B2(n_84), .Y(n_251) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_203), .A2(n_140), .B(n_197), .Y(n_252) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_221), .A2(n_197), .B(n_191), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_207), .Y(n_254) );
INVx8_ASAP7_75t_L g255 ( .A(n_206), .Y(n_255) );
INVx1_ASAP7_75t_SL g256 ( .A(n_213), .Y(n_256) );
OAI21x1_ASAP7_75t_L g257 ( .A1(n_204), .A2(n_191), .B(n_185), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_244), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_234), .B(n_229), .Y(n_259) );
OR2x6_ASAP7_75t_L g260 ( .A(n_255), .B(n_224), .Y(n_260) );
AOI21xp33_ASAP7_75t_L g261 ( .A1(n_251), .A2(n_228), .B(n_223), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_238), .B(n_219), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_231), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_247), .A2(n_229), .B(n_217), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_242), .A2(n_219), .B1(n_212), .B2(n_191), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_238), .B(n_214), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_239), .A2(n_199), .B1(n_202), .B2(n_209), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_244), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_239), .B(n_214), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_234), .B(n_212), .Y(n_270) );
AOI221xp5_ASAP7_75t_L g271 ( .A1(n_236), .A2(n_183), .B1(n_220), .B2(n_226), .C(n_224), .Y(n_271) );
AOI221xp5_ASAP7_75t_L g272 ( .A1(n_236), .A2(n_211), .B1(n_227), .B2(n_117), .C(n_118), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_235), .B(n_206), .Y(n_273) );
OR2x6_ASAP7_75t_L g274 ( .A(n_255), .B(n_200), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_256), .B(n_199), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_244), .Y(n_276) );
OAI211xp5_ASAP7_75t_L g277 ( .A1(n_233), .A2(n_117), .B(n_118), .C(n_129), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_243), .A2(n_191), .B1(n_251), .B2(n_256), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_254), .Y(n_279) );
OAI22xp33_ASAP7_75t_L g280 ( .A1(n_235), .A2(n_210), .B1(n_178), .B2(n_205), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_258), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_258), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_258), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_268), .Y(n_284) );
INVx2_ASAP7_75t_SL g285 ( .A(n_263), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_268), .Y(n_286) );
NAND2x1p5_ASAP7_75t_L g287 ( .A(n_263), .B(n_231), .Y(n_287) );
OAI221xp5_ASAP7_75t_L g288 ( .A1(n_265), .A2(n_249), .B1(n_246), .B2(n_240), .C(n_245), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_268), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_259), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_262), .B(n_191), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_276), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_276), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_276), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_259), .B(n_246), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_259), .B(n_254), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_279), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_279), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_279), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_259), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_266), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_270), .Y(n_302) );
AOI221xp5_ASAP7_75t_L g303 ( .A1(n_302), .A2(n_270), .B1(n_261), .B2(n_267), .C(n_271), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_296), .B(n_273), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_301), .B(n_266), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_281), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_282), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_283), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_283), .B(n_267), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_286), .B(n_263), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_302), .B(n_269), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_286), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_290), .A2(n_269), .B1(n_278), .B2(n_273), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_288), .B(n_292), .C(n_297), .Y(n_315) );
OAI33xp33_ASAP7_75t_L g316 ( .A1(n_291), .A2(n_280), .A3(n_275), .B1(n_7), .B2(n_8), .B3(n_9), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_292), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_297), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_295), .B(n_273), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_281), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_300), .A2(n_273), .B1(n_272), .B2(n_260), .Y(n_321) );
OAI221xp5_ASAP7_75t_L g322 ( .A1(n_300), .A2(n_249), .B1(n_277), .B2(n_264), .C(n_241), .Y(n_322) );
OAI21xp5_ASAP7_75t_SL g323 ( .A1(n_295), .A2(n_263), .B(n_241), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_296), .B(n_254), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_284), .B(n_263), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_284), .B(n_263), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_289), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_289), .A2(n_248), .B(n_247), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_293), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_295), .B(n_4), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_285), .B(n_274), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_293), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_307), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_317), .B(n_294), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_317), .B(n_294), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_307), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_308), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_308), .B(n_298), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_306), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_305), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_305), .B(n_299), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_312), .B(n_299), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_309), .B(n_298), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_309), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_313), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_313), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_318), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_318), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_332), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_306), .B(n_285), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_306), .B(n_287), .Y(n_351) );
NAND4xp25_ASAP7_75t_L g352 ( .A(n_330), .B(n_5), .C(n_7), .D(n_9), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_327), .B(n_287), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_332), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_324), .B(n_287), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_310), .B(n_245), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_324), .B(n_240), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_327), .B(n_253), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_327), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_325), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_325), .B(n_253), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_320), .Y(n_362) );
INVx2_ASAP7_75t_SL g363 ( .A(n_311), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_311), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_326), .B(n_253), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_303), .B(n_240), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_304), .B(n_240), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_320), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_319), .B(n_5), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_311), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_304), .B(n_310), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_329), .B(n_326), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_329), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_311), .B(n_315), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_331), .B(n_231), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_315), .B(n_253), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_340), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_333), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_374), .B(n_331), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_333), .Y(n_380) );
INVx2_ASAP7_75t_SL g381 ( .A(n_375), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_336), .Y(n_382) );
INVxp67_ASAP7_75t_L g383 ( .A(n_374), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_360), .B(n_331), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_371), .B(n_323), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_341), .B(n_323), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_336), .Y(n_387) );
OAI21xp5_ASAP7_75t_L g388 ( .A1(n_352), .A2(n_328), .B(n_321), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_337), .B(n_314), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_339), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_337), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_370), .B(n_331), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_344), .B(n_10), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_344), .Y(n_394) );
OR2x6_ASAP7_75t_L g395 ( .A(n_375), .B(n_260), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_372), .B(n_10), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_370), .B(n_11), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_364), .B(n_11), .Y(n_398) );
OAI21xp5_ASAP7_75t_L g399 ( .A1(n_352), .A2(n_247), .B(n_257), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_345), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_369), .A2(n_316), .B1(n_260), .B2(n_322), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_363), .B(n_12), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_345), .B(n_13), .Y(n_403) );
INVx1_ASAP7_75t_SL g404 ( .A(n_342), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_346), .B(n_15), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_339), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_363), .B(n_274), .Y(n_407) );
XNOR2xp5_ASAP7_75t_L g408 ( .A(n_375), .B(n_15), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_338), .B(n_16), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_346), .B(n_17), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_347), .Y(n_411) );
OAI31xp33_ASAP7_75t_L g412 ( .A1(n_366), .A2(n_241), .A3(n_18), .B(n_19), .Y(n_412) );
NOR2x1_ASAP7_75t_SL g413 ( .A(n_335), .B(n_274), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_347), .B(n_17), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_348), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_348), .Y(n_416) );
NAND3xp33_ASAP7_75t_L g417 ( .A(n_376), .B(n_129), .C(n_118), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_349), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_356), .B(n_18), .Y(n_419) );
INVx3_ASAP7_75t_SL g420 ( .A(n_375), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_362), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_376), .A2(n_248), .B(n_274), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_335), .B(n_231), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_349), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_354), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_356), .B(n_19), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_354), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_338), .B(n_245), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_377), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_421), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_388), .A2(n_355), .B1(n_367), .B2(n_353), .Y(n_431) );
INVx1_ASAP7_75t_SL g432 ( .A(n_420), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_408), .A2(n_357), .B1(n_373), .B2(n_368), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_404), .B(n_343), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_385), .B(n_343), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_378), .Y(n_436) );
OAI21xp5_ASAP7_75t_L g437 ( .A1(n_419), .A2(n_257), .B(n_351), .Y(n_437) );
NOR2xp33_ASAP7_75t_R g438 ( .A(n_420), .B(n_353), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_384), .B(n_350), .Y(n_439) );
AOI21xp33_ASAP7_75t_L g440 ( .A1(n_419), .A2(n_373), .B(n_368), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_426), .A2(n_351), .B1(n_361), .B2(n_365), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_379), .B(n_350), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_426), .B(n_334), .Y(n_443) );
AOI322xp5_ASAP7_75t_L g444 ( .A1(n_383), .A2(n_365), .A3(n_361), .B1(n_358), .B2(n_334), .C1(n_359), .C2(n_362), .Y(n_444) );
OAI22xp33_ASAP7_75t_SL g445 ( .A1(n_395), .A2(n_359), .B1(n_362), .B2(n_260), .Y(n_445) );
OAI21xp33_ASAP7_75t_SL g446 ( .A1(n_423), .A2(n_358), .B(n_274), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_421), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_380), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_383), .B(n_129), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_389), .B(n_245), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_396), .B(n_129), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_386), .B(n_245), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_414), .B(n_129), .Y(n_453) );
AO22x1_ASAP7_75t_L g454 ( .A1(n_397), .A2(n_381), .B1(n_379), .B2(n_407), .Y(n_454) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_412), .A2(n_257), .B(n_241), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_382), .B(n_252), .Y(n_456) );
OAI222xp33_ASAP7_75t_L g457 ( .A1(n_395), .A2(n_260), .B1(n_231), .B2(n_255), .C1(n_205), .C2(n_250), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_401), .A2(n_232), .B(n_237), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_379), .B(n_237), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_409), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_387), .B(n_252), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_392), .B(n_237), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_391), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_414), .A2(n_255), .B(n_232), .C(n_231), .Y(n_464) );
NAND3xp33_ASAP7_75t_L g465 ( .A(n_423), .B(n_231), .C(n_153), .Y(n_465) );
AOI211xp5_ASAP7_75t_L g466 ( .A1(n_398), .A2(n_232), .B(n_255), .C(n_178), .Y(n_466) );
OAI221xp5_ASAP7_75t_L g467 ( .A1(n_399), .A2(n_250), .B1(n_252), .B2(n_153), .C(n_144), .Y(n_467) );
OAI21xp33_ASAP7_75t_L g468 ( .A1(n_402), .A2(n_200), .B(n_23), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_394), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_400), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_407), .A2(n_250), .B1(n_252), .B2(n_200), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_411), .B(n_153), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_395), .Y(n_473) );
INVxp67_ASAP7_75t_L g474 ( .A(n_413), .Y(n_474) );
AO22x2_ASAP7_75t_L g475 ( .A1(n_429), .A2(n_418), .B1(n_427), .B2(n_425), .Y(n_475) );
INVxp67_ASAP7_75t_L g476 ( .A(n_451), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_436), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_448), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_463), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g480 ( .A1(n_431), .A2(n_405), .B1(n_403), .B2(n_410), .C(n_393), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_431), .B(n_415), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_446), .B(n_417), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_433), .A2(n_407), .B1(n_416), .B2(n_424), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_469), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_444), .B(n_406), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_435), .B(n_406), .Y(n_486) );
XNOR2xp5_ASAP7_75t_L g487 ( .A(n_432), .B(n_422), .Y(n_487) );
AOI322xp5_ASAP7_75t_L g488 ( .A1(n_460), .A2(n_428), .A3(n_390), .B1(n_422), .B2(n_153), .C1(n_144), .C2(n_200), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_441), .B(n_390), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_473), .A2(n_250), .B1(n_144), .B2(n_25), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_442), .B(n_144), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_445), .B(n_144), .Y(n_492) );
INVxp33_ASAP7_75t_L g493 ( .A(n_438), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_439), .B(n_144), .Y(n_494) );
INVx2_ASAP7_75t_SL g495 ( .A(n_454), .Y(n_495) );
NOR3xp33_ASAP7_75t_L g496 ( .A(n_451), .B(n_250), .C(n_24), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_434), .B(n_21), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_474), .A2(n_26), .B(n_27), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_449), .Y(n_499) );
OAI311xp33_ASAP7_75t_L g500 ( .A1(n_458), .A2(n_72), .A3(n_36), .B1(n_37), .C1(n_40), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_452), .B(n_69), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_474), .B(n_34), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_443), .Y(n_503) );
XOR2xp5_ASAP7_75t_L g504 ( .A(n_462), .B(n_42), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_SL g505 ( .A1(n_493), .A2(n_457), .B(n_464), .C(n_440), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_475), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_493), .A2(n_453), .B1(n_437), .B2(n_470), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_499), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_495), .Y(n_509) );
NAND3xp33_ASAP7_75t_L g510 ( .A(n_492), .B(n_455), .C(n_465), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_499), .B(n_450), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_475), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_475), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_476), .A2(n_468), .B1(n_459), .B2(n_466), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_481), .B(n_430), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_480), .A2(n_482), .B1(n_495), .B2(n_503), .Y(n_516) );
AOI221xp5_ASAP7_75t_L g517 ( .A1(n_485), .A2(n_467), .B1(n_472), .B2(n_457), .C(n_447), .Y(n_517) );
BUFx3_ASAP7_75t_L g518 ( .A(n_494), .Y(n_518) );
OAI21xp33_ASAP7_75t_L g519 ( .A1(n_487), .A2(n_467), .B(n_471), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_477), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_483), .A2(n_482), .B1(n_489), .B2(n_491), .Y(n_521) );
INVxp33_ASAP7_75t_L g522 ( .A(n_492), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g523 ( .A1(n_505), .A2(n_478), .B1(n_479), .B2(n_484), .C(n_486), .Y(n_523) );
AOI221x1_ASAP7_75t_L g524 ( .A1(n_506), .A2(n_496), .B1(n_498), .B2(n_497), .C(n_501), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_509), .B(n_488), .Y(n_525) );
AOI321xp33_ASAP7_75t_L g526 ( .A1(n_516), .A2(n_502), .A3(n_490), .B1(n_504), .B2(n_461), .C(n_456), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_508), .Y(n_527) );
INVx2_ASAP7_75t_SL g528 ( .A(n_518), .Y(n_528) );
CKINVDCx6p67_ASAP7_75t_R g529 ( .A(n_522), .Y(n_529) );
OAI211xp5_ASAP7_75t_L g530 ( .A1(n_516), .A2(n_502), .B(n_500), .C(n_45), .Y(n_530) );
OAI22xp33_ASAP7_75t_L g531 ( .A1(n_522), .A2(n_43), .B1(n_44), .B2(n_46), .Y(n_531) );
AOI21xp33_ASAP7_75t_L g532 ( .A1(n_513), .A2(n_47), .B(n_48), .Y(n_532) );
NOR3xp33_ASAP7_75t_SL g533 ( .A(n_530), .B(n_510), .C(n_519), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_527), .Y(n_534) );
AOI321xp33_ASAP7_75t_L g535 ( .A1(n_523), .A2(n_521), .A3(n_517), .B1(n_507), .B2(n_512), .C(n_514), .Y(n_535) );
NAND4xp25_ASAP7_75t_SL g536 ( .A(n_523), .B(n_505), .C(n_515), .D(n_511), .Y(n_536) );
NAND2x1_ASAP7_75t_SL g537 ( .A(n_525), .B(n_520), .Y(n_537) );
NOR4xp25_ASAP7_75t_L g538 ( .A(n_536), .B(n_529), .C(n_528), .D(n_526), .Y(n_538) );
INVxp67_ASAP7_75t_SL g539 ( .A(n_534), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_533), .Y(n_540) );
NAND3xp33_ASAP7_75t_L g541 ( .A(n_540), .B(n_535), .C(n_524), .Y(n_541) );
OAI22x1_ASAP7_75t_L g542 ( .A1(n_540), .A2(n_537), .B1(n_532), .B2(n_531), .Y(n_542) );
OAI22xp5_ASAP7_75t_SL g543 ( .A1(n_541), .A2(n_538), .B1(n_539), .B2(n_532), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_542), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_544), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_545), .A2(n_543), .B(n_56), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_546), .A2(n_53), .B1(n_58), .B2(n_60), .Y(n_547) );
AO221x1_ASAP7_75t_L g548 ( .A1(n_547), .A2(n_61), .B1(n_62), .B2(n_66), .C(n_68), .Y(n_548) );
endmodule