module fake_jpeg_22018_n_345 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_44),
.Y(n_71)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_41),
.B(n_42),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_0),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_31),
.B1(n_18),
.B2(n_29),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_53),
.A2(n_61),
.B1(n_70),
.B2(n_77),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_57),
.Y(n_83)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_62),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_31),
.B1(n_18),
.B2(n_33),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_31),
.B1(n_29),
.B2(n_19),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_74),
.Y(n_100)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_72),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_29),
.B1(n_17),
.B2(n_25),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_46),
.B1(n_43),
.B2(n_37),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_37),
.A2(n_25),
.B1(n_23),
.B2(n_17),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_80),
.Y(n_99)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_84),
.B(n_86),
.Y(n_134)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_41),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_87),
.B(n_88),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_63),
.Y(n_88)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_93),
.Y(n_145)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_0),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_94),
.B(n_8),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_42),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_97),
.Y(n_136)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_107),
.Y(n_143)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

BUFx4f_ASAP7_75t_SL g111 ( 
.A(n_63),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_47),
.Y(n_113)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_117),
.B1(n_118),
.B2(n_24),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_16),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_79),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_55),
.A2(n_23),
.B1(n_34),
.B2(n_35),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_27),
.Y(n_146)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_68),
.B1(n_56),
.B2(n_52),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_124),
.A2(n_128),
.B1(n_142),
.B2(n_148),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_50),
.B1(n_48),
.B2(n_38),
.Y(n_128)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_50),
.C(n_48),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_139),
.C(n_121),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_101),
.A2(n_65),
.B1(n_35),
.B2(n_34),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_147),
.B1(n_112),
.B2(n_96),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_26),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_94),
.A2(n_27),
.B1(n_24),
.B2(n_20),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_86),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_116),
.A2(n_33),
.B1(n_32),
.B2(n_27),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_114),
.A2(n_27),
.B1(n_24),
.B2(n_20),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_149),
.B(n_88),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_111),
.B1(n_108),
.B2(n_92),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_154),
.A2(n_162),
.B1(n_165),
.B2(n_176),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_143),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_156),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_157),
.A2(n_160),
.B(n_152),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_99),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_166),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_128),
.A2(n_120),
.B1(n_90),
.B2(n_83),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_146),
.B1(n_140),
.B2(n_136),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_111),
.B(n_85),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_161),
.B(n_168),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_177),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_125),
.B(n_110),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_98),
.Y(n_167)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_167),
.Y(n_214)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_133),
.A2(n_97),
.B(n_93),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_169),
.A2(n_179),
.B(n_186),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_115),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_170),
.Y(n_218)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_173),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_127),
.B(n_10),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_177),
.Y(n_189)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_130),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_175),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_0),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_149),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_178),
.A2(n_183),
.B1(n_129),
.B2(n_123),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_133),
.A2(n_26),
.B(n_20),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_0),
.Y(n_182)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_122),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_132),
.B(n_1),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_187),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_138),
.A2(n_92),
.B1(n_24),
.B2(n_20),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_185),
.A2(n_7),
.B1(n_12),
.B2(n_10),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_132),
.A2(n_149),
.B(n_126),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_126),
.B(n_26),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_195),
.B1(n_200),
.B2(n_201),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_140),
.C(n_144),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_206),
.C(n_210),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_211),
.B(n_213),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_155),
.A2(n_146),
.B1(n_136),
.B2(n_144),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_169),
.A2(n_152),
.B(n_151),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_197),
.A2(n_179),
.B(n_187),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_155),
.A2(n_146),
.B1(n_151),
.B2(n_129),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_123),
.B1(n_89),
.B2(n_16),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_202),
.A2(n_205),
.B1(n_178),
.B2(n_165),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_89),
.B1(n_16),
.B2(n_26),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_26),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_216),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_153),
.B(n_26),
.C(n_2),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_160),
.A2(n_1),
.B(n_2),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_6),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_217),
.C(n_172),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_157),
.A2(n_1),
.B(n_2),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_153),
.B(n_3),
.Y(n_215)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_154),
.B(n_7),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_168),
.B(n_3),
.C(n_4),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_219),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_190),
.B(n_164),
.Y(n_221)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_199),
.A2(n_162),
.B1(n_171),
.B2(n_180),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_224),
.A2(n_239),
.B1(n_246),
.B2(n_247),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_156),
.Y(n_227)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_228),
.A2(n_235),
.B(n_236),
.Y(n_268)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_193),
.B(n_170),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_230),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_174),
.Y(n_231)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_231),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_203),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_232),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_183),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_166),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_196),
.A2(n_186),
.B(n_167),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_202),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_185),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_241),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_182),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_248),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_189),
.B(n_173),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_245),
.B(n_208),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_201),
.A2(n_161),
.B1(n_184),
.B2(n_175),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_219),
.B1(n_209),
.B2(n_208),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_189),
.B(n_3),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_192),
.B(n_6),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g249 ( 
.A1(n_243),
.A2(n_209),
.B(n_194),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_249),
.A2(n_264),
.B1(n_266),
.B2(n_270),
.Y(n_282)
);

NAND4xp25_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_204),
.C(n_214),
.D(n_197),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_251),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_224),
.A2(n_195),
.B1(n_191),
.B2(n_196),
.Y(n_252)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_238),
.A2(n_198),
.B1(n_216),
.B2(n_212),
.Y(n_259)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_259),
.Y(n_283)
);

BUFx4f_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_228),
.A2(n_236),
.B(n_225),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_SL g281 ( 
.A1(n_263),
.A2(n_242),
.B(n_5),
.C(n_4),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_222),
.B1(n_246),
.B2(n_223),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_210),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_257),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_223),
.A2(n_211),
.B1(n_217),
.B2(n_213),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_229),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_244),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_268),
.A2(n_225),
.B(n_235),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_272),
.A2(n_279),
.B(n_251),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_237),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_280),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_237),
.C(n_240),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_288),
.C(n_263),
.Y(n_294)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_241),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_277),
.B(n_284),
.Y(n_302)
);

FAx1_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_245),
.CI(n_226),
.CON(n_279),
.SN(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_248),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_281),
.B(n_271),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_9),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_262),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_286),
.Y(n_301)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_267),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_282),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_9),
.C(n_10),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_289),
.B(n_268),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_289),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_292),
.A2(n_281),
.B(n_265),
.Y(n_318)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_290),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_293),
.A2(n_303),
.B(n_253),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_275),
.C(n_253),
.Y(n_311)
);

NOR3xp33_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_250),
.C(n_254),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_278),
.Y(n_307)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_299),
.Y(n_309)
);

BUFx5_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_252),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_272),
.B(n_261),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_258),
.Y(n_306)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_311),
.C(n_315),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_317),
.B(n_318),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_298),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_273),
.B1(n_255),
.B2(n_281),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_313),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_314),
.B(n_293),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_256),
.C(n_255),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_259),
.Y(n_317)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_321),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_292),
.B(n_301),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_326),
.C(n_308),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_291),
.C(n_304),
.Y(n_326)
);

AO22x1_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_312),
.B1(n_316),
.B2(n_318),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_296),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_331),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_333),
.C(n_327),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_319),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_334),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_325),
.A2(n_309),
.B(n_305),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_305),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_335),
.A2(n_332),
.B(n_330),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_320),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_336),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_338),
.Y(n_341)
);

O2A1O1Ixp33_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_339),
.B(n_337),
.C(n_320),
.Y(n_342)
);

AO21x1_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_281),
.B(n_15),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_15),
.B(n_5),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_5),
.Y(n_345)
);


endmodule