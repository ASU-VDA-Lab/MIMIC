module fake_jpeg_14183_n_203 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_7),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_5),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_7),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_40),
.B(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_25),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_41),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_5),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_54),
.Y(n_65)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_15),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_18),
.B(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_8),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_21),
.B(n_8),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_26),
.B(n_2),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_57),
.Y(n_73)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_1),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_25),
.B(n_1),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_27),
.C(n_32),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_59),
.A2(n_32),
.B1(n_38),
.B2(n_57),
.Y(n_91)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_26),
.B(n_4),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_31),
.B(n_28),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_67),
.B(n_39),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_13),
.B1(n_34),
.B2(n_30),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_13),
.B1(n_34),
.B2(n_30),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_78),
.B1(n_91),
.B2(n_93),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_83),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_23),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_88),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_37),
.A2(n_23),
.B1(n_20),
.B2(n_19),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_72),
.A2(n_82),
.B1(n_90),
.B2(n_71),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_20),
.B(n_19),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_67),
.C(n_83),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_41),
.A2(n_27),
.B1(n_35),
.B2(n_32),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_9),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_84),
.B(n_94),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_50),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_36),
.A2(n_32),
.B1(n_11),
.B2(n_12),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_39),
.B(n_47),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_51),
.B1(n_54),
.B2(n_39),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_85),
.B1(n_76),
.B2(n_62),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_96),
.B(n_99),
.Y(n_144)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_86),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_64),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_101),
.B(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_65),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_63),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_110),
.B(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_119),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_115),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_75),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_118),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_77),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_75),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_93),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_121),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_92),
.Y(n_121)
);

NOR2xp67_ASAP7_75t_SL g122 ( 
.A(n_91),
.B(n_72),
.Y(n_122)
);

NAND2x1_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_62),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_71),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_142),
.C(n_106),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_139),
.B1(n_120),
.B2(n_103),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_85),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_132),
.B(n_133),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_74),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_116),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_140),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_98),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_74),
.B1(n_122),
.B2(n_114),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_74),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_113),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_154),
.C(n_158),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_113),
.B1(n_112),
.B2(n_102),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_148),
.A2(n_159),
.B1(n_130),
.B2(n_129),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_139),
.A2(n_112),
.B1(n_98),
.B2(n_109),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_157),
.Y(n_165)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_151),
.B(n_153),
.Y(n_167)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_134),
.A2(n_143),
.B1(n_138),
.B2(n_125),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_99),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_138),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_159)
);

AOI32xp33_ASAP7_75t_L g161 ( 
.A1(n_125),
.A2(n_132),
.A3(n_137),
.B1(n_133),
.B2(n_144),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_SL g174 ( 
.A(n_161),
.B(n_144),
.C(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_162),
.B(n_163),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_123),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_135),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_SL g181 ( 
.A(n_164),
.B(n_170),
.C(n_174),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_175),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_137),
.C(n_124),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_144),
.B(n_136),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_167),
.B(n_171),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_145),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_145),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_131),
.Y(n_185)
);

BUFx12_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_179),
.B1(n_184),
.B2(n_169),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_165),
.A2(n_156),
.B1(n_149),
.B2(n_154),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_172),
.A2(n_151),
.B(n_158),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_180),
.A2(n_173),
.B1(n_168),
.B2(n_166),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_163),
.C(n_162),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_183),
.C(n_185),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_165),
.A2(n_150),
.B(n_152),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_167),
.B1(n_174),
.B2(n_171),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_190),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_189),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_177),
.A2(n_173),
.B1(n_126),
.B2(n_131),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_184),
.A2(n_126),
.B1(n_180),
.B2(n_183),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_179),
.B(n_181),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_188),
.B(n_182),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_178),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_SL g197 ( 
.A1(n_193),
.A2(n_189),
.B(n_190),
.C(n_185),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_193),
.A2(n_188),
.B(n_186),
.C(n_191),
.Y(n_196)
);

A2O1A1O1Ixp25_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_197),
.B(n_194),
.C(n_195),
.D(n_178),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_198),
.B(n_195),
.Y(n_199)
);

OAI21x1_ASAP7_75t_SL g201 ( 
.A1(n_199),
.A2(n_200),
.B(n_194),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_178),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_126),
.Y(n_203)
);


endmodule