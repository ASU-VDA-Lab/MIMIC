module fake_jpeg_19829_n_173 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx2_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_5),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_15),
.Y(n_50)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_41),
.Y(n_66)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_0),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx2_ASAP7_75t_SL g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_48),
.B(n_50),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_19),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_64),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_18),
.B1(n_30),
.B2(n_24),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_18),
.B1(n_17),
.B2(n_31),
.Y(n_70)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_25),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_28),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_69),
.B1(n_57),
.B2(n_65),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_71),
.B(n_83),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_74),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_30),
.B1(n_18),
.B2(n_21),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_35),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_88),
.C(n_40),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_21),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_86),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_27),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_49),
.B(n_45),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_54),
.B(n_25),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_59),
.Y(n_100)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_69),
.B1(n_59),
.B2(n_47),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_102),
.B1(n_106),
.B2(n_91),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_28),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_86),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_23),
.Y(n_104)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_69),
.B1(n_65),
.B2(n_57),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_98),
.A2(n_83),
.B1(n_70),
.B2(n_85),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_31),
.B(n_107),
.Y(n_126)
);

AO22x2_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_106),
.B1(n_103),
.B2(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_114),
.B(n_116),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_76),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_119),
.C(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_72),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_23),
.C(n_107),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_122),
.Y(n_130)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_92),
.B(n_88),
.CI(n_53),
.CON(n_122),
.SN(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_108),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_132),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_110),
.A2(n_73),
.B1(n_88),
.B2(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_113),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_129),
.B(n_138),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_136),
.Y(n_139)
);

AOI221xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_75),
.B1(n_27),
.B2(n_95),
.C(n_22),
.Y(n_134)
);

OAI322xp33_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_111),
.A3(n_27),
.B1(n_22),
.B2(n_119),
.C1(n_115),
.C2(n_42),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_122),
.A2(n_96),
.B1(n_108),
.B2(n_73),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_142),
.A2(n_145),
.B(n_146),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_112),
.C(n_118),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_143),
.B(n_144),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_112),
.C(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_121),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_SL g150 ( 
.A(n_148),
.B(n_130),
.C(n_126),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_152),
.Y(n_156)
);

OAI321xp33_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_112),
.A3(n_143),
.B1(n_141),
.B2(n_133),
.C(n_127),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_141),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_SL g152 ( 
.A(n_139),
.B(n_136),
.C(n_129),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_144),
.A2(n_135),
.B1(n_79),
.B2(n_87),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_154),
.B1(n_1),
.B2(n_2),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_61),
.B1(n_2),
.B2(n_3),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_158),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_42),
.C(n_84),
.Y(n_158)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_4),
.C(n_7),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_4),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_1),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_150),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_165),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_156),
.B1(n_161),
.B2(n_158),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_167),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_12),
.Y(n_167)
);

AOI31xp67_ASAP7_75t_SL g170 ( 
.A1(n_168),
.A2(n_162),
.A3(n_12),
.B(n_13),
.Y(n_170)
);

AOI21x1_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_14),
.B(n_3),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_169),
.B(n_14),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g173 ( 
.A(n_172),
.Y(n_173)
);


endmodule