module fake_jpeg_3637_n_248 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_12),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_46),
.B(n_50),
.Y(n_121)
);

HAxp5_ASAP7_75t_SL g47 ( 
.A(n_19),
.B(n_21),
.CON(n_47),
.SN(n_47)
);

HAxp5_ASAP7_75t_SL g101 ( 
.A(n_47),
.B(n_48),
.CON(n_101),
.SN(n_101)
);

HAxp5_ASAP7_75t_SL g48 ( 
.A(n_21),
.B(n_0),
.CON(n_48),
.SN(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_3),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_4),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_61),
.B(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_16),
.B(n_4),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_6),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_65),
.B(n_73),
.Y(n_102)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_30),
.B(n_11),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_16),
.B(n_6),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_38),
.B(n_7),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_7),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_22),
.B(n_8),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_76),
.B(n_22),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

BUFx16f_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_27),
.Y(n_95)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_27),
.B1(n_36),
.B2(n_34),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_82),
.A2(n_119),
.B1(n_8),
.B2(n_10),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_103),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_25),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_96),
.B(n_105),
.Y(n_150)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_25),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_68),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_33),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_42),
.B(n_33),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_106),
.B(n_107),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_44),
.B(n_26),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_43),
.B(n_26),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_115),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_59),
.B(n_29),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_45),
.A2(n_29),
.B1(n_34),
.B2(n_36),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_51),
.B(n_37),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_90),
.Y(n_149)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_37),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_136),
.Y(n_159)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

BUFx24_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_125),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_126),
.B(n_137),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_82),
.A2(n_57),
.B1(n_54),
.B2(n_80),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_129),
.A2(n_135),
.B1(n_138),
.B2(n_152),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_93),
.A2(n_66),
.B1(n_72),
.B2(n_77),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_130),
.A2(n_132),
.B(n_142),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g131 ( 
.A(n_89),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_149),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_101),
.A2(n_77),
.B1(n_58),
.B2(n_74),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_8),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_SL g163 ( 
.A(n_134),
.B(n_143),
.C(n_99),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_10),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_87),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_10),
.B1(n_85),
.B2(n_97),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_94),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_140),
.B(n_144),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_100),
.A2(n_108),
.B(n_91),
.Y(n_142)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_81),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_116),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_85),
.A2(n_92),
.B1(n_97),
.B2(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_152),
.Y(n_161)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_148),
.Y(n_175)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_88),
.B(n_104),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_153),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_117),
.A2(n_118),
.B1(n_88),
.B2(n_84),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_94),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_156),
.B(n_111),
.Y(n_165)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_166),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_127),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_125),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_104),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_98),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_98),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_99),
.C(n_126),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_179),
.C(n_128),
.Y(n_192)
);

NAND2x1_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_99),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_130),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_122),
.B(n_156),
.C(n_142),
.Y(n_179)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_138),
.B1(n_145),
.B2(n_140),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_196),
.B1(n_200),
.B2(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_187),
.B(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

HAxp5_ASAP7_75t_SL g203 ( 
.A(n_190),
.B(n_172),
.CON(n_203),
.SN(n_203)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_195),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_193),
.C(n_180),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_148),
.C(n_146),
.Y(n_193)
);

NOR4xp25_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_143),
.C(n_150),
.D(n_134),
.Y(n_194)
);

NOR4xp25_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_174),
.C(n_160),
.D(n_176),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_155),
.B1(n_139),
.B2(n_154),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_197),
.B(n_198),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_183),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_133),
.B1(n_157),
.B2(n_141),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

OAI321xp33_ASAP7_75t_L g204 ( 
.A1(n_201),
.A2(n_159),
.A3(n_169),
.B1(n_166),
.B2(n_163),
.C(n_171),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_206),
.B(n_188),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_210),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_SL g211 ( 
.A1(n_201),
.A2(n_176),
.B(n_174),
.C(n_177),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_190),
.B(n_186),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_214),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_158),
.C(n_165),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_170),
.B1(n_178),
.B2(n_164),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_202),
.Y(n_224)
);

AO221x1_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_200),
.B1(n_196),
.B2(n_177),
.C(n_191),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_212),
.Y(n_232)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_224),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_219),
.A2(n_211),
.B1(n_203),
.B2(n_209),
.Y(n_226)
);

AOI321xp33_ASAP7_75t_L g228 ( 
.A1(n_223),
.A2(n_188),
.A3(n_211),
.B1(n_214),
.B2(n_208),
.C(n_205),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_211),
.A2(n_186),
.B(n_193),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_185),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_232),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_213),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_227),
.B(n_230),
.Y(n_235)
);

NOR3xp33_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_231),
.C(n_225),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_212),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_229),
.A2(n_221),
.B1(n_220),
.B2(n_222),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_178),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_234),
.A2(n_237),
.B(n_230),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_226),
.A2(n_219),
.B1(n_184),
.B2(n_162),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_227),
.Y(n_238)
);

INVxp33_ASAP7_75t_SL g244 ( 
.A(n_238),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_241),
.C(n_177),
.Y(n_243)
);

AOI322xp5_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_236),
.A3(n_162),
.B1(n_158),
.B2(n_175),
.C1(n_237),
.C2(n_124),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_175),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_243),
.B(n_241),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_246),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g246 ( 
.A(n_244),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_177),
.Y(n_248)
);


endmodule