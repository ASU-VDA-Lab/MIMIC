module fake_netlist_1_2015_n_885 (n_103, n_52, n_50, n_7, n_3, n_34, n_25, n_9, n_96, n_72, n_77, n_90, n_99, n_43, n_73, n_62, n_97, n_33, n_4, n_59, n_76, n_6, n_74, n_8, n_61, n_44, n_66, n_88, n_46, n_37, n_18, n_65, n_87, n_5, n_81, n_85, n_102, n_47, n_1, n_16, n_78, n_95, n_40, n_68, n_36, n_11, n_15, n_71, n_70, n_94, n_2, n_17, n_58, n_20, n_84, n_12, n_56, n_80, n_67, n_22, n_19, n_26, n_39, n_101, n_98, n_38, n_104, n_100, n_24, n_35, n_91, n_32, n_93, n_48, n_63, n_54, n_41, n_55, n_29, n_60, n_10, n_30, n_13, n_92, n_75, n_82, n_53, n_64, n_69, n_83, n_23, n_0, n_57, n_51, n_45, n_42, n_21, n_86, n_27, n_89, n_28, n_79, n_49, n_14, n_31, n_885, n_884);
input n_103;
input n_52;
input n_50;
input n_7;
input n_3;
input n_34;
input n_25;
input n_9;
input n_96;
input n_72;
input n_77;
input n_90;
input n_99;
input n_43;
input n_73;
input n_62;
input n_97;
input n_33;
input n_4;
input n_59;
input n_76;
input n_6;
input n_74;
input n_8;
input n_61;
input n_44;
input n_66;
input n_88;
input n_46;
input n_37;
input n_18;
input n_65;
input n_87;
input n_5;
input n_81;
input n_85;
input n_102;
input n_47;
input n_1;
input n_16;
input n_78;
input n_95;
input n_40;
input n_68;
input n_36;
input n_11;
input n_15;
input n_71;
input n_70;
input n_94;
input n_2;
input n_17;
input n_58;
input n_20;
input n_84;
input n_12;
input n_56;
input n_80;
input n_67;
input n_22;
input n_19;
input n_26;
input n_39;
input n_101;
input n_98;
input n_38;
input n_104;
input n_100;
input n_24;
input n_35;
input n_91;
input n_32;
input n_93;
input n_48;
input n_63;
input n_54;
input n_41;
input n_55;
input n_29;
input n_60;
input n_10;
input n_30;
input n_13;
input n_92;
input n_75;
input n_82;
input n_53;
input n_64;
input n_69;
input n_83;
input n_23;
input n_0;
input n_57;
input n_51;
input n_45;
input n_42;
input n_21;
input n_86;
input n_27;
input n_89;
input n_28;
input n_79;
input n_49;
input n_14;
input n_31;
output n_885;
output n_884;
wire n_107;
wire n_646;
wire n_759;
wire n_658;
wire n_673;
wire n_156;
wire n_154;
wire n_239;
wire n_7;
wire n_309;
wire n_356;
wire n_327;
wire n_25;
wire n_204;
wire n_592;
wire n_769;
wire n_169;
wire n_370;
wire n_384;
wire n_439;
wire n_545;
wire n_180;
wire n_604;
wire n_99;
wire n_43;
wire n_73;
wire n_440;
wire n_199;
wire n_279;
wire n_786;
wire n_831;
wire n_357;
wire n_74;
wire n_729;
wire n_308;
wire n_518;
wire n_44;
wire n_394;
wire n_189;
wire n_681;
wire n_226;
wire n_352;
wire n_447;
wire n_66;
wire n_379;
wire n_535;
wire n_689;
wire n_595;
wire n_875;
wire n_626;
wire n_316;
wire n_285;
wire n_564;
wire n_586;
wire n_471;
wire n_47;
wire n_766;
wire n_475;
wire n_744;
wire n_850;
wire n_281;
wire n_645;
wire n_497;
wire n_399;
wire n_11;
wire n_295;
wire n_371;
wire n_579;
wire n_516;
wire n_608;
wire n_368;
wire n_805;
wire n_373;
wire n_139;
wire n_342;
wire n_151;
wire n_71;
wire n_288;
wire n_557;
wire n_176;
wire n_753;
wire n_859;
wire n_436;
wire n_438;
wire n_869;
wire n_359;
wire n_195;
wire n_300;
wire n_487;
wire n_461;
wire n_723;
wire n_223;
wire n_833;
wire n_405;
wire n_830;
wire n_562;
wire n_19;
wire n_409;
wire n_482;
wire n_838;
wire n_534;
wire n_569;
wire n_707;
wire n_526;
wire n_261;
wire n_483;
wire n_423;
wire n_220;
wire n_353;
wire n_410;
wire n_104;
wire n_709;
wire n_303;
wire n_502;
wire n_821;
wire n_468;
wire n_159;
wire n_566;
wire n_91;
wire n_301;
wire n_340;
wire n_148;
wire n_149;
wire n_567;
wire n_378;
wire n_752;
wire n_246;
wire n_676;
wire n_823;
wire n_191;
wire n_143;
wire n_780;
wire n_864;
wire n_629;
wire n_446;
wire n_63;
wire n_402;
wire n_54;
wire n_876;
wire n_387;
wire n_125;
wire n_145;
wire n_166;
wire n_558;
wire n_596;
wire n_492;
wire n_181;
wire n_123;
wire n_219;
wire n_343;
wire n_494;
wire n_555;
wire n_553;
wire n_135;
wire n_481;
wire n_621;
wire n_817;
wire n_776;
wire n_315;
wire n_397;
wire n_53;
wire n_880;
wire n_213;
wire n_196;
wire n_293;
wire n_797;
wire n_836;
wire n_127;
wire n_312;
wire n_742;
wire n_424;
wire n_23;
wire n_110;
wire n_182;
wire n_269;
wire n_663;
wire n_529;
wire n_656;
wire n_751;
wire n_186;
wire n_137;
wire n_507;
wire n_334;
wire n_164;
wire n_433;
wire n_806;
wire n_120;
wire n_392;
wire n_650;
wire n_660;
wire n_155;
wire n_162;
wire n_114;
wire n_772;
wire n_50;
wire n_789;
wire n_816;
wire n_3;
wire n_331;
wire n_651;
wire n_574;
wire n_882;
wire n_636;
wire n_330;
wire n_614;
wire n_231;
wire n_884;
wire n_9;
wire n_737;
wire n_428;
wire n_178;
wire n_478;
wire n_814;
wire n_652;
wire n_678;
wire n_708;
wire n_229;
wire n_97;
wire n_133;
wire n_324;
wire n_442;
wire n_422;
wire n_192;
wire n_699;
wire n_857;
wire n_329;
wire n_6;
wire n_8;
wire n_578;
wire n_187;
wire n_548;
wire n_188;
wire n_443;
wire n_304;
wire n_18;
wire n_682;
wire n_801;
wire n_441;
wire n_868;
wire n_628;
wire n_425;
wire n_314;
wire n_824;
wire n_601;
wire n_307;
wire n_517;
wire n_215;
wire n_736;
wire n_172;
wire n_109;
wire n_332;
wire n_198;
wire n_386;
wire n_653;
wire n_351;
wire n_1;
wire n_16;
wire n_670;
wire n_95;
wire n_40;
wire n_210;
wire n_426;
wire n_755;
wire n_716;
wire n_228;
wire n_863;
wire n_671;
wire n_278;
wire n_115;
wire n_270;
wire n_476;
wire n_765;
wire n_829;
wire n_599;
wire n_715;
wire n_849;
wire n_179;
wire n_289;
wire n_404;
wire n_366;
wire n_721;
wire n_362;
wire n_617;
wire n_688;
wire n_837;
wire n_485;
wire n_396;
wire n_549;
wire n_354;
wire n_720;
wire n_152;
wire n_851;
wire n_70;
wire n_588;
wire n_458;
wire n_375;
wire n_855;
wire n_17;
wire n_322;
wire n_317;
wire n_221;
wire n_328;
wire n_506;
wire n_711;
wire n_491;
wire n_800;
wire n_388;
wire n_773;
wire n_266;
wire n_763;
wire n_80;
wire n_632;
wire n_793;
wire n_679;
wire n_522;
wire n_546;
wire n_615;
wire n_684;
wire n_701;
wire n_326;
wire n_532;
wire n_756;
wire n_635;
wire n_544;
wire n_879;
wire n_576;
wire n_275;
wire n_691;
wire n_622;
wire n_661;
wire n_493;
wire n_274;
wire n_150;
wire n_235;
wire n_690;
wire n_38;
wire n_533;
wire n_272;
wire n_686;
wire n_299;
wire n_100;
wire n_561;
wire n_581;
wire n_280;
wire n_141;
wire n_509;
wire n_160;
wire n_499;
wire n_377;
wire n_263;
wire n_757;
wire n_844;
wire n_695;
wire n_193;
wire n_232;
wire n_344;
wire n_878;
wire n_783;
wire n_812;
wire n_147;
wire n_185;
wire n_367;
wire n_795;
wire n_267;
wire n_687;
wire n_171;
wire n_638;
wire n_873;
wire n_450;
wire n_585;
wire n_140;
wire n_644;
wire n_111;
wire n_779;
wire n_212;
wire n_746;
wire n_30;
wire n_634;
wire n_13;
wire n_254;
wire n_559;
wire n_704;
wire n_435;
wire n_728;
wire n_583;
wire n_841;
wire n_64;
wire n_69;
wire n_248;
wire n_866;
wire n_407;
wire n_527;
wire n_83;
wire n_200;
wire n_603;
wire n_262;
wire n_119;
wire n_667;
wire n_503;
wire n_856;
wire n_339;
wire n_347;
wire n_124;
wire n_696;
wire n_748;
wire n_79;
wire n_129;
wire n_611;
wire n_521;
wire n_157;
wire n_774;
wire n_103;
wire n_808;
wire n_421;
wire n_52;
wire n_253;
wire n_434;
wire n_677;
wire n_624;
wire n_273;
wire n_325;
wire n_571;
wire n_524;
wire n_692;
wire n_530;
wire n_743;
wire n_163;
wire n_348;
wire n_96;
wire n_685;
wire n_669;
wire n_77;
wire n_72;
wire n_90;
wire n_594;
wire n_762;
wire n_214;
wire n_740;
wire n_787;
wire n_770;
wire n_167;
wire n_861;
wire n_809;
wire n_364;
wire n_33;
wire n_464;
wire n_76;
wire n_470;
wire n_590;
wire n_61;
wire n_463;
wire n_216;
wire n_153;
wire n_355;
wire n_609;
wire n_121;
wire n_286;
wire n_408;
wire n_247;
wire n_431;
wire n_161;
wire n_224;
wire n_484;
wire n_165;
wire n_860;
wire n_413;
wire n_65;
wire n_537;
wire n_710;
wire n_525;
wire n_560;
wire n_5;
wire n_496;
wire n_393;
wire n_843;
wire n_211;
wire n_85;
wire n_320;
wire n_264;
wire n_102;
wire n_283;
wire n_733;
wire n_846;
wire n_290;
wire n_217;
wire n_201;
wire n_791;
wire n_792;
wire n_277;
wire n_259;
wire n_612;
wire n_244;
wire n_666;
wire n_771;
wire n_827;
wire n_276;
wire n_297;
wire n_225;
wire n_631;
wire n_350;
wire n_747;
wire n_208;
wire n_616;
wire n_815;
wire n_523;
wire n_854;
wire n_528;
wire n_419;
wire n_252;
wire n_519;
wire n_168;
wire n_839;
wire n_271;
wire n_693;
wire n_785;
wire n_739;
wire n_94;
wire n_194;
wire n_858;
wire n_758;
wire n_825;
wire n_282;
wire n_58;
wire n_775;
wire n_113;
wire n_242;
wire n_498;
wire n_501;
wire n_321;
wire n_284;
wire n_302;
wire n_538;
wire n_703;
wire n_811;
wire n_116;
wire n_734;
wire n_292;
wire n_547;
wire n_593;
wire n_118;
wire n_587;
wire n_233;
wire n_597;
wire n_554;
wire n_698;
wire n_705;
wire n_257;
wire n_741;
wire n_828;
wire n_722;
wire n_203;
wire n_26;
wire n_477;
wire n_460;
wire n_243;
wire n_318;
wire n_346;
wire n_98;
wire n_345;
wire n_230;
wire n_452;
wire n_714;
wire n_146;
wire n_337;
wire n_32;
wire n_726;
wire n_641;
wire n_637;
wire n_531;
wire n_872;
wire n_93;
wire n_539;
wire n_847;
wire n_406;
wire n_372;
wire n_842;
wire n_820;
wire n_713;
wire n_467;
wire n_702;
wire n_41;
wire n_760;
wire n_826;
wire n_623;
wire n_417;
wire n_451;
wire n_665;
wire n_647;
wire n_445;
wire n_500;
wire n_732;
wire n_845;
wire n_575;
wire n_10;
wire n_390;
wire n_600;
wire n_818;
wire n_75;
wire n_82;
wire n_183;
wire n_731;
wire n_550;
wire n_132;
wire n_643;
wire n_761;
wire n_778;
wire n_582;
wire n_784;
wire n_170;
wire n_205;
wire n_158;
wire n_126;
wire n_473;
wire n_249;
wire n_389;
wire n_834;
wire n_510;
wire n_360;
wire n_363;
wire n_749;
wire n_427;
wire n_724;
wire n_106;
wire n_296;
wire n_605;
wire n_42;
wire n_21;
wire n_835;
wire n_437;
wire n_871;
wire n_620;
wire n_89;
wire n_480;
wire n_130;
wire n_341;
wire n_310;
wire n_700;
wire n_640;
wire n_14;
wire n_236;
wire n_639;
wire n_727;
wire n_136;
wire n_260;
wire n_580;
wire n_610;
wire n_222;
wire n_657;
wire n_822;
wire n_381;
wire n_142;
wire n_34;
wire n_853;
wire n_754;
wire n_385;
wire n_798;
wire n_227;
wire n_395;
wire n_454;
wire n_453;
wire n_250;
wire n_551;
wire n_268;
wire n_190;
wire n_606;
wire n_62;
wire n_712;
wire n_777;
wire n_4;
wire n_59;
wire n_323;
wire n_565;
wire n_781;
wire n_852;
wire n_376;
wire n_694;
wire n_240;
wire n_459;
wire n_768;
wire n_88;
wire n_568;
wire n_46;
wire n_174;
wire n_717;
wire n_807;
wire n_108;
wire n_335;
wire n_37;
wire n_122;
wire n_374;
wire n_613;
wire n_380;
wire n_515;
wire n_802;
wire n_865;
wire n_672;
wire n_867;
wire n_87;
wire n_466;
wire n_349;
wire n_207;
wire n_197;
wire n_81;
wire n_541;
wire n_572;
wire n_298;
wire n_112;
wire n_630;
wire n_735;
wire n_649;
wire n_602;
wire n_78;
wire n_552;
wire n_68;
wire n_444;
wire n_105;
wire n_251;
wire n_598;
wire n_810;
wire n_36;
wire n_416;
wire n_870;
wire n_432;
wire n_465;
wire n_414;
wire n_680;
wire n_730;
wire n_469;
wire n_369;
wire n_361;
wire n_767;
wire n_237;
wire n_881;
wire n_654;
wire n_15;
wire n_520;
wire n_633;
wire n_429;
wire n_803;
wire n_256;
wire n_398;
wire n_668;
wire n_117;
wire n_238;
wire n_365;
wire n_577;
wire n_796;
wire n_804;
wire n_294;
wire n_2;
wire n_338;
wire n_662;
wire n_591;
wire n_391;
wire n_241;
wire n_209;
wire n_874;
wire n_20;
wire n_84;
wire n_782;
wire n_449;
wire n_832;
wire n_56;
wire n_12;
wire n_412;
wire n_455;
wire n_67;
wire n_504;
wire n_618;
wire n_790;
wire n_456;
wire n_22;
wire n_683;
wire n_479;
wire n_584;
wire n_311;
wire n_401;
wire n_877;
wire n_383;
wire n_813;
wire n_202;
wire n_319;
wire n_542;
wire n_725;
wire n_819;
wire n_862;
wire n_39;
wire n_101;
wire n_291;
wire n_489;
wire n_245;
wire n_664;
wire n_508;
wire n_764;
wire n_719;
wire n_486;
wire n_788;
wire n_24;
wire n_35;
wire n_655;
wire n_490;
wire n_472;
wire n_540;
wire n_840;
wire n_400;
wire n_794;
wire n_457;
wire n_659;
wire n_134;
wire n_48;
wire n_255;
wire n_563;
wire n_513;
wire n_55;
wire n_718;
wire n_543;
wire n_336;
wire n_29;
wire n_218;
wire n_173;
wire n_556;
wire n_488;
wire n_648;
wire n_382;
wire n_799;
wire n_138;
wire n_60;
wire n_462;
wire n_573;
wire n_536;
wire n_474;
wire n_745;
wire n_305;
wire n_495;
wire n_430;
wire n_418;
wire n_505;
wire n_92;
wire n_313;
wire n_333;
wire n_358;
wire n_627;
wire n_750;
wire n_706;
wire n_589;
wire n_175;
wire n_128;
wire n_306;
wire n_415;
wire n_697;
wire n_0;
wire n_512;
wire n_258;
wire n_675;
wire n_619;
wire n_642;
wire n_234;
wire n_607;
wire n_848;
wire n_184;
wire n_265;
wire n_57;
wire n_674;
wire n_51;
wire n_570;
wire n_411;
wire n_514;
wire n_287;
wire n_144;
wire n_403;
wire n_625;
wire n_45;
wire n_131;
wire n_420;
wire n_86;
wire n_27;
wire n_738;
wire n_177;
wire n_28;
wire n_511;
wire n_448;
wire n_49;
wire n_206;
wire n_31;
INVx1_ASAP7_75t_L g105 ( .A(n_2), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_54), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_21), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_53), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_43), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_62), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_65), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_87), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_33), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_96), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_35), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_77), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_36), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_71), .Y(n_119) );
CKINVDCx14_ASAP7_75t_R g120 ( .A(n_79), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_63), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_93), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_32), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_55), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_1), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_95), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_44), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_74), .Y(n_128) );
BUFx3_ASAP7_75t_L g129 ( .A(n_88), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_50), .Y(n_130) );
CKINVDCx14_ASAP7_75t_R g131 ( .A(n_68), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_9), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_80), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_15), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_6), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_17), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_41), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_104), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_92), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_28), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_94), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_22), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_56), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_125), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_138), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_138), .B(n_0), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_138), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_138), .B(n_0), .Y(n_148) );
BUFx8_ASAP7_75t_L g149 ( .A(n_140), .Y(n_149) );
INVx5_ASAP7_75t_L g150 ( .A(n_119), .Y(n_150) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_105), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_114), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_119), .Y(n_153) );
NAND3xp33_ASAP7_75t_L g154 ( .A(n_105), .B(n_47), .C(n_102), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_134), .B(n_1), .Y(n_155) );
OAI22xp5_ASAP7_75t_SL g156 ( .A1(n_134), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_114), .B(n_3), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_140), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_119), .Y(n_159) );
INVx6_ASAP7_75t_L g160 ( .A(n_124), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_132), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_124), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_132), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_140), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_120), .B(n_4), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_108), .Y(n_167) );
NOR2xp33_ASAP7_75t_R g168 ( .A(n_149), .B(n_131), .Y(n_168) );
INVx2_ASAP7_75t_SL g169 ( .A(n_149), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_149), .B(n_106), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_151), .B(n_135), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_147), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_147), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_166), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
INVxp33_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
INVx2_ASAP7_75t_SL g177 ( .A(n_148), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_161), .B(n_124), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_152), .B(n_129), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_148), .B(n_107), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_147), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_145), .B(n_110), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_155), .A2(n_122), .B1(n_128), .B2(n_141), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_153), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_153), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_148), .B(n_112), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_145), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_153), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_158), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_158), .Y(n_191) );
CKINVDCx6p67_ASAP7_75t_R g192 ( .A(n_166), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_155), .B(n_116), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_155), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_157), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_165), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_153), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_165), .Y(n_198) );
INVx8_ASAP7_75t_L g199 ( .A(n_157), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_167), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_167), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_157), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_146), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_153), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_150), .B(n_123), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_162), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_163), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_160), .B(n_126), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_162), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_162), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_164), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_150), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_150), .B(n_136), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_162), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_159), .A2(n_136), .B1(n_109), .B2(n_111), .Y(n_215) );
NOR2xp33_ASAP7_75t_R g216 ( .A(n_192), .B(n_137), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_193), .B(n_160), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_174), .B(n_160), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_183), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_174), .B(n_160), .Y(n_220) );
INVxp67_ASAP7_75t_L g221 ( .A(n_184), .Y(n_221) );
NAND2xp33_ASAP7_75t_L g222 ( .A(n_169), .B(n_130), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_199), .B(n_133), .Y(n_223) );
OAI22xp33_ASAP7_75t_L g224 ( .A1(n_176), .A2(n_127), .B1(n_118), .B2(n_109), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_169), .B(n_154), .Y(n_225) );
AND2x2_ASAP7_75t_SL g226 ( .A(n_202), .B(n_111), .Y(n_226) );
NOR2xp33_ASAP7_75t_R g227 ( .A(n_192), .B(n_139), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_199), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_199), .B(n_142), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_168), .B(n_143), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_180), .B(n_113), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_194), .B(n_113), .Y(n_232) );
OAI221xp5_ASAP7_75t_L g233 ( .A1(n_195), .A2(n_156), .B1(n_115), .B2(n_127), .C(n_118), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_199), .A2(n_121), .B1(n_115), .B2(n_108), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_183), .Y(n_235) );
NAND3xp33_ASAP7_75t_L g236 ( .A(n_187), .B(n_150), .C(n_159), .Y(n_236) );
INVx2_ASAP7_75t_SL g237 ( .A(n_171), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_203), .B(n_121), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_199), .B(n_150), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_183), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_203), .B(n_117), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_178), .B(n_159), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_177), .B(n_117), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_202), .B(n_129), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_171), .B(n_159), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_172), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_207), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_190), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_177), .A2(n_162), .B(n_129), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_170), .B(n_18), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_182), .B(n_5), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_188), .B(n_19), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_188), .A2(n_5), .B(n_6), .C(n_7), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_207), .B(n_7), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_208), .B(n_52), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_172), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_211), .B(n_8), .Y(n_257) );
OAI221xp5_ASAP7_75t_L g258 ( .A1(n_211), .A2(n_8), .B1(n_9), .B2(n_10), .C(n_11), .Y(n_258) );
CKINVDCx11_ASAP7_75t_R g259 ( .A(n_200), .Y(n_259) );
INVxp67_ASAP7_75t_L g260 ( .A(n_200), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_201), .B(n_10), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_201), .B(n_11), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_205), .B(n_59), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_190), .B(n_12), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_179), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_191), .B(n_13), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_213), .B(n_15), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_191), .B(n_16), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_173), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_173), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_196), .B(n_16), .Y(n_271) );
AO21x1_ASAP7_75t_L g272 ( .A1(n_252), .A2(n_175), .B(n_214), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_247), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_226), .B(n_196), .Y(n_274) );
INVxp67_ASAP7_75t_L g275 ( .A(n_237), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_226), .B(n_198), .Y(n_276) );
OR2x6_ASAP7_75t_L g277 ( .A(n_228), .B(n_213), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_248), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g279 ( .A1(n_238), .A2(n_175), .B(n_215), .Y(n_279) );
O2A1O1Ixp33_ASAP7_75t_L g280 ( .A1(n_221), .A2(n_198), .B(n_181), .C(n_206), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_259), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_228), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_260), .A2(n_181), .B1(n_212), .B2(n_206), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_248), .B(n_212), .Y(n_284) );
AND2x6_ASAP7_75t_SL g285 ( .A(n_231), .B(n_17), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_243), .A2(n_214), .B(n_186), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_232), .B(n_212), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_231), .B(n_212), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_243), .A2(n_214), .B(n_186), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_239), .A2(n_185), .B(n_186), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_238), .B(n_206), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_224), .B(n_206), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_241), .A2(n_189), .B(n_185), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_264), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_227), .B(n_204), .Y(n_295) );
NAND3xp33_ASAP7_75t_L g296 ( .A(n_222), .B(n_210), .C(n_209), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_267), .B(n_210), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_245), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g299 ( .A1(n_233), .A2(n_209), .B(n_197), .C(n_189), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_230), .B(n_197), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_241), .A2(n_189), .B(n_185), .Y(n_301) );
OA22x2_ASAP7_75t_L g302 ( .A1(n_216), .A2(n_20), .B1(n_23), .B2(n_24), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_244), .A2(n_204), .B(n_26), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_216), .B(n_204), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_254), .Y(n_305) );
AO32x1_ASAP7_75t_L g306 ( .A1(n_253), .A2(n_204), .A3(n_27), .B1(n_29), .B2(n_30), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_244), .A2(n_204), .B(n_31), .Y(n_307) );
O2A1O1Ixp33_ASAP7_75t_L g308 ( .A1(n_258), .A2(n_204), .B(n_34), .C(n_37), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_242), .A2(n_25), .B(n_38), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_249), .A2(n_39), .B(n_40), .Y(n_310) );
NOR2x1_ASAP7_75t_L g311 ( .A(n_254), .B(n_42), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_267), .A2(n_45), .B1(n_46), .B2(n_48), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_227), .B(n_223), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_266), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g315 ( .A1(n_257), .A2(n_49), .B1(n_51), .B2(n_57), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_294), .B(n_234), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_305), .A2(n_229), .B1(n_218), .B2(n_220), .Y(n_317) );
AO31x2_ASAP7_75t_L g318 ( .A1(n_272), .A2(n_261), .A3(n_262), .B(n_268), .Y(n_318) );
AOI21x1_ASAP7_75t_L g319 ( .A1(n_303), .A2(n_255), .B(n_252), .Y(n_319) );
OAI21xp5_ASAP7_75t_L g320 ( .A1(n_280), .A2(n_251), .B(n_250), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_273), .B(n_217), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_275), .A2(n_217), .B1(n_265), .B2(n_271), .C(n_236), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_277), .B(n_225), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_274), .B(n_250), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_276), .A2(n_298), .B1(n_277), .B2(n_292), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_277), .B(n_225), .Y(n_326) );
AOI21x1_ASAP7_75t_L g327 ( .A1(n_307), .A2(n_219), .B(n_235), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_282), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_297), .A2(n_263), .B1(n_240), .B2(n_270), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_282), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_282), .B(n_263), .Y(n_331) );
AOI221x1_ASAP7_75t_L g332 ( .A1(n_309), .A2(n_269), .B1(n_256), .B2(n_246), .C(n_64), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_291), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_299), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_290), .A2(n_58), .B(n_60), .Y(n_335) );
AOI21xp33_ASAP7_75t_L g336 ( .A1(n_304), .A2(n_61), .B(n_66), .Y(n_336) );
OAI21x1_ASAP7_75t_L g337 ( .A1(n_311), .A2(n_67), .B(n_69), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_288), .A2(n_70), .B(n_72), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_278), .Y(n_339) );
OAI21x1_ASAP7_75t_L g340 ( .A1(n_310), .A2(n_73), .B(n_75), .Y(n_340) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_293), .A2(n_76), .B(n_78), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_313), .B(n_81), .Y(n_342) );
INVx4_ASAP7_75t_L g343 ( .A(n_302), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_328), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_327), .Y(n_345) );
OAI21x1_ASAP7_75t_L g346 ( .A1(n_332), .A2(n_319), .B(n_341), .Y(n_346) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_341), .A2(n_301), .B(n_286), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_333), .Y(n_348) );
NAND2x1p5_ASAP7_75t_L g349 ( .A(n_343), .B(n_314), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_328), .Y(n_350) );
OA21x2_ASAP7_75t_L g351 ( .A1(n_320), .A2(n_315), .B(n_312), .Y(n_351) );
AO31x2_ASAP7_75t_L g352 ( .A1(n_334), .A2(n_289), .A3(n_283), .B(n_300), .Y(n_352) );
OAI21x1_ASAP7_75t_L g353 ( .A1(n_340), .A2(n_295), .B(n_315), .Y(n_353) );
NAND2x1p5_ASAP7_75t_L g354 ( .A(n_343), .B(n_314), .Y(n_354) );
OAI21x1_ASAP7_75t_L g355 ( .A1(n_340), .A2(n_308), .B(n_279), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_316), .B(n_285), .Y(n_356) );
BUFx6f_ASAP7_75t_SL g357 ( .A(n_343), .Y(n_357) );
INVx6_ASAP7_75t_L g358 ( .A(n_328), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_325), .B(n_281), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_323), .B(n_287), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_328), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_323), .B(n_314), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_324), .A2(n_306), .B(n_296), .Y(n_363) );
INVxp67_ASAP7_75t_SL g364 ( .A(n_330), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_321), .Y(n_365) );
OA21x2_ASAP7_75t_L g366 ( .A1(n_337), .A2(n_306), .B(n_284), .Y(n_366) );
OA21x2_ASAP7_75t_L g367 ( .A1(n_337), .A2(n_306), .B(n_83), .Y(n_367) );
NOR2x1_ASAP7_75t_R g368 ( .A(n_342), .B(n_323), .Y(n_368) );
OAI21x1_ASAP7_75t_L g369 ( .A1(n_335), .A2(n_82), .B(n_84), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_326), .B(n_85), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_326), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_339), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_348), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_348), .B(n_318), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_365), .B(n_318), .Y(n_375) );
OAI21x1_ASAP7_75t_L g376 ( .A1(n_346), .A2(n_338), .B(n_331), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_344), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_345), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_372), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_372), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_345), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_365), .B(n_318), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
NAND2x1_ASAP7_75t_L g384 ( .A(n_350), .B(n_342), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_349), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_345), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_349), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_344), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_344), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_361), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_346), .Y(n_391) );
BUFx10_ASAP7_75t_L g392 ( .A(n_357), .Y(n_392) );
AO31x2_ASAP7_75t_L g393 ( .A1(n_363), .A2(n_317), .A3(n_329), .B(n_318), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_361), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_367), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_367), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_370), .B(n_342), .Y(n_397) );
AO21x2_ASAP7_75t_L g398 ( .A1(n_355), .A2(n_336), .B(n_322), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_354), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_367), .Y(n_400) );
INVxp67_ASAP7_75t_L g401 ( .A(n_368), .Y(n_401) );
OAI21x1_ASAP7_75t_L g402 ( .A1(n_353), .A2(n_339), .B(n_89), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_370), .B(n_339), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_361), .Y(n_404) );
BUFx3_ASAP7_75t_L g405 ( .A(n_358), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_354), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_367), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_366), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_354), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_366), .Y(n_410) );
AO21x2_ASAP7_75t_L g411 ( .A1(n_355), .A2(n_86), .B(n_90), .Y(n_411) );
INVx3_ASAP7_75t_L g412 ( .A(n_357), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_350), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_359), .B(n_91), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_357), .Y(n_415) );
AO21x2_ASAP7_75t_L g416 ( .A1(n_353), .A2(n_97), .B(n_98), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_358), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_368), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_350), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_373), .B(n_356), .Y(n_420) );
INVxp67_ASAP7_75t_L g421 ( .A(n_414), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_375), .B(n_362), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_375), .B(n_362), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_374), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_374), .B(n_359), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_375), .B(n_362), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_378), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_374), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_378), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_388), .Y(n_430) );
NOR2xp33_ASAP7_75t_R g431 ( .A(n_392), .B(n_357), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_378), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_382), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_414), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_414), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_382), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_382), .B(n_362), .Y(n_437) );
AND2x2_ASAP7_75t_SL g438 ( .A(n_418), .B(n_351), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_381), .Y(n_439) );
INVx4_ASAP7_75t_SL g440 ( .A(n_418), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_381), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_381), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_386), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_386), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_373), .B(n_352), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_379), .B(n_352), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_379), .B(n_352), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_386), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_380), .B(n_352), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_380), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_408), .Y(n_451) );
BUFx3_ASAP7_75t_L g452 ( .A(n_392), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_388), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_408), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_408), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_410), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_410), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_389), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_410), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_395), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_395), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_395), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_396), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_396), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_397), .B(n_364), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_396), .Y(n_466) );
INVxp67_ASAP7_75t_L g467 ( .A(n_389), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_400), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_400), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_394), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_400), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_407), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_394), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_390), .B(n_350), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_390), .B(n_352), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_401), .B(n_371), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_407), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_407), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_419), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_390), .B(n_352), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_413), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_391), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_392), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_391), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_419), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_397), .B(n_351), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_391), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_402), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_397), .B(n_351), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_413), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_403), .B(n_351), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_403), .B(n_360), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_377), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_393), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_403), .B(n_366), .Y(n_495) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_383), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_393), .B(n_366), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_452), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_450), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_486), .B(n_393), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_486), .B(n_393), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_489), .B(n_393), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_422), .B(n_406), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_450), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_455), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_420), .B(n_401), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_425), .B(n_385), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_483), .B(n_412), .Y(n_508) );
INVxp67_ASAP7_75t_L g509 ( .A(n_496), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_424), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_424), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_425), .B(n_385), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_455), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_428), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_433), .B(n_399), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_428), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_455), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_479), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_489), .B(n_393), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_433), .B(n_399), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_436), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_436), .B(n_393), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_465), .B(n_406), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_481), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_422), .B(n_390), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_483), .B(n_415), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_423), .B(n_390), .Y(n_527) );
INVx4_ASAP7_75t_L g528 ( .A(n_452), .Y(n_528) );
AND2x4_ASAP7_75t_L g529 ( .A(n_475), .B(n_415), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_457), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_485), .Y(n_531) );
AND2x4_ASAP7_75t_L g532 ( .A(n_475), .B(n_415), .Y(n_532) );
BUFx2_ASAP7_75t_L g533 ( .A(n_431), .Y(n_533) );
INVxp67_ASAP7_75t_L g534 ( .A(n_453), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_423), .B(n_377), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_475), .B(n_415), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_481), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_426), .B(n_387), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_457), .Y(n_539) );
INVx3_ASAP7_75t_L g540 ( .A(n_457), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_490), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_452), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_490), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_458), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_473), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_465), .Y(n_546) );
OAI221xp5_ASAP7_75t_L g547 ( .A1(n_476), .A2(n_384), .B1(n_409), .B2(n_387), .C(n_383), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_426), .B(n_409), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_430), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_475), .B(n_415), .Y(n_550) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_430), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_492), .B(n_404), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_474), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_459), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_437), .B(n_404), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_492), .B(n_404), .Y(n_556) );
NAND2x1p5_ASAP7_75t_L g557 ( .A(n_474), .B(n_412), .Y(n_557) );
NAND2x1p5_ASAP7_75t_L g558 ( .A(n_474), .B(n_412), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_434), .B(n_412), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_451), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_437), .B(n_417), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_445), .B(n_412), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_435), .B(n_417), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_451), .Y(n_564) );
INVx5_ASAP7_75t_L g565 ( .A(n_474), .Y(n_565) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_467), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_470), .B(n_417), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_445), .B(n_405), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_491), .B(n_377), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_491), .B(n_377), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_459), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_454), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_495), .B(n_377), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_421), .B(n_405), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_454), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_456), .B(n_377), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_456), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_446), .B(n_405), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_439), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_459), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_440), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_446), .B(n_377), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_495), .B(n_416), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_439), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_440), .B(n_392), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_462), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_438), .A2(n_384), .B1(n_441), .B2(n_442), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_441), .B(n_398), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_442), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_462), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_443), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_447), .B(n_392), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_443), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_447), .B(n_416), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_462), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_449), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_449), .B(n_416), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_464), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_427), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_497), .B(n_398), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_564), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_596), .B(n_497), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_500), .B(n_480), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_518), .B(n_448), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_546), .B(n_494), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_506), .B(n_438), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_555), .B(n_480), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_564), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_544), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_568), .B(n_480), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_545), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_524), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_561), .B(n_480), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_534), .B(n_438), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_525), .B(n_493), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_500), .B(n_494), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_521), .B(n_461), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_525), .B(n_493), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_527), .B(n_444), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_580), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_537), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_527), .B(n_444), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_501), .B(n_460), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_541), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_518), .B(n_444), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_510), .B(n_472), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_580), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_566), .B(n_477), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_543), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_501), .B(n_460), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_511), .B(n_463), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_540), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_533), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_531), .B(n_427), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_514), .B(n_463), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_516), .B(n_469), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_540), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_531), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_499), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_504), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_535), .B(n_448), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_535), .B(n_448), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_528), .B(n_440), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_572), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_502), .B(n_471), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_592), .B(n_432), .Y(n_646) );
AND2x4_ASAP7_75t_L g647 ( .A(n_529), .B(n_440), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_572), .Y(n_648) );
BUFx2_ASAP7_75t_L g649 ( .A(n_528), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_503), .B(n_432), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_507), .B(n_432), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_538), .B(n_429), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_502), .B(n_469), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_540), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_505), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_560), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_519), .B(n_472), .Y(n_657) );
INVx2_ASAP7_75t_SL g658 ( .A(n_528), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_519), .B(n_471), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_505), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_512), .B(n_427), .Y(n_661) );
INVx1_ASAP7_75t_SL g662 ( .A(n_498), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_513), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_575), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_552), .B(n_429), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_522), .B(n_461), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_513), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_522), .B(n_515), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_529), .B(n_440), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_517), .Y(n_670) );
NAND2xp33_ASAP7_75t_L g671 ( .A(n_585), .B(n_429), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_520), .B(n_477), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_509), .B(n_478), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_577), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_579), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_584), .Y(n_676) );
OR2x2_ASAP7_75t_L g677 ( .A(n_556), .B(n_478), .Y(n_677) );
INVx1_ASAP7_75t_SL g678 ( .A(n_542), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_517), .Y(n_679) );
OR2x2_ASAP7_75t_L g680 ( .A(n_578), .B(n_468), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_548), .B(n_468), .Y(n_681) );
INVx1_ASAP7_75t_SL g682 ( .A(n_523), .Y(n_682) );
INVxp67_ASAP7_75t_L g683 ( .A(n_549), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_573), .B(n_466), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_589), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_573), .B(n_466), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_591), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_530), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_530), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_562), .B(n_464), .Y(n_690) );
AND2x4_ASAP7_75t_SL g691 ( .A(n_529), .B(n_487), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_593), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_549), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_569), .B(n_487), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_567), .B(n_487), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_569), .B(n_484), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_551), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_563), .B(n_484), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_551), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_570), .B(n_484), .Y(n_700) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_598), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_559), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_599), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_508), .Y(n_704) );
INVx2_ASAP7_75t_SL g705 ( .A(n_633), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_638), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_612), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_603), .B(n_532), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_603), .B(n_532), .Y(n_709) );
INVxp67_ASAP7_75t_L g710 ( .A(n_649), .Y(n_710) );
OR2x2_ASAP7_75t_L g711 ( .A(n_623), .B(n_582), .Y(n_711) );
NOR2xp67_ASAP7_75t_L g712 ( .A(n_658), .B(n_585), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_621), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_607), .B(n_550), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_623), .B(n_550), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_616), .B(n_600), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_624), .Y(n_717) );
INVx3_ASAP7_75t_L g718 ( .A(n_647), .Y(n_718) );
INVxp67_ASAP7_75t_L g719 ( .A(n_662), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_629), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_616), .B(n_597), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_630), .B(n_597), .Y(n_722) );
OAI21xp33_ASAP7_75t_SL g723 ( .A1(n_643), .A2(n_526), .B(n_508), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_701), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_609), .B(n_547), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_639), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_630), .B(n_550), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_645), .B(n_594), .Y(n_728) );
OR2x2_ASAP7_75t_L g729 ( .A(n_645), .B(n_570), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_611), .B(n_574), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_640), .Y(n_731) );
OR2x2_ASAP7_75t_L g732 ( .A(n_653), .B(n_553), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_701), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_653), .B(n_583), .Y(n_734) );
NAND2x2_ASAP7_75t_L g735 ( .A(n_658), .B(n_581), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_677), .Y(n_736) );
OR2x2_ASAP7_75t_L g737 ( .A(n_657), .B(n_576), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_682), .B(n_526), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_656), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_657), .B(n_583), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_659), .B(n_610), .Y(n_741) );
NAND3xp33_ASAP7_75t_SL g742 ( .A(n_643), .B(n_557), .C(n_558), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_664), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_659), .B(n_588), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_613), .B(n_532), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_646), .B(n_536), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_644), .B(n_586), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_606), .A2(n_536), .B1(n_587), .B2(n_565), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_674), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_675), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_648), .B(n_571), .Y(n_751) );
INVxp67_ASAP7_75t_SL g752 ( .A(n_601), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_678), .B(n_536), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_676), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_685), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_702), .B(n_565), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_687), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_692), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_693), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_697), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_601), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_681), .B(n_565), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_668), .B(n_565), .Y(n_763) );
NAND4xp75_ASAP7_75t_L g764 ( .A(n_614), .B(n_598), .C(n_595), .D(n_590), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_619), .B(n_557), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_699), .B(n_595), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_622), .B(n_558), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_673), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_666), .B(n_590), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_615), .B(n_586), .Y(n_770) );
OR2x2_ASAP7_75t_L g771 ( .A(n_602), .B(n_571), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_618), .B(n_554), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_665), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_690), .B(n_554), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_628), .Y(n_775) );
INVxp67_ASAP7_75t_SL g776 ( .A(n_608), .Y(n_776) );
OAI33xp33_ASAP7_75t_L g777 ( .A1(n_605), .A2(n_539), .A3(n_488), .B1(n_482), .B2(n_416), .B3(n_411), .Y(n_777) );
NOR2xp67_ASAP7_75t_SL g778 ( .A(n_704), .B(n_358), .Y(n_778) );
INVx1_ASAP7_75t_SL g779 ( .A(n_691), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_628), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_707), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_768), .B(n_683), .Y(n_782) );
OR2x6_ASAP7_75t_L g783 ( .A(n_712), .B(n_669), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_713), .Y(n_784) );
OAI22xp33_ASAP7_75t_L g785 ( .A1(n_735), .A2(n_669), .B1(n_647), .B2(n_606), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_717), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_720), .Y(n_787) );
INVx2_ASAP7_75t_SL g788 ( .A(n_705), .Y(n_788) );
NAND2x1p5_ASAP7_75t_L g789 ( .A(n_779), .B(n_647), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_775), .B(n_683), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_719), .B(n_614), .Y(n_791) );
NAND3xp33_ASAP7_75t_L g792 ( .A(n_723), .B(n_608), .C(n_671), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_726), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_731), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_718), .A2(n_669), .B1(n_691), .B2(n_680), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_780), .B(n_650), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_739), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_742), .A2(n_671), .B1(n_652), .B2(n_627), .Y(n_798) );
OAI221xp5_ASAP7_75t_L g799 ( .A1(n_725), .A2(n_695), .B1(n_698), .B2(n_672), .C(n_604), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_773), .B(n_641), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_724), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_743), .Y(n_802) );
OR2x2_ASAP7_75t_L g803 ( .A(n_744), .B(n_634), .Y(n_803) );
OAI21xp5_ASAP7_75t_L g804 ( .A1(n_710), .A2(n_625), .B(n_620), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_749), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_730), .A2(n_620), .B1(n_627), .B2(n_696), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_750), .Y(n_807) );
NAND3xp33_ASAP7_75t_SL g808 ( .A(n_779), .B(n_661), .C(n_651), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_753), .B(n_684), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_754), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g811 ( .A1(n_752), .A2(n_617), .B(n_636), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_716), .B(n_642), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_716), .B(n_686), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_755), .Y(n_814) );
OR2x2_ASAP7_75t_L g815 ( .A(n_744), .B(n_694), .Y(n_815) );
OAI21xp5_ASAP7_75t_SL g816 ( .A1(n_748), .A2(n_700), .B(n_696), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_757), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_758), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_736), .B(n_700), .Y(n_819) );
O2A1O1Ixp5_ASAP7_75t_R g820 ( .A1(n_721), .A2(n_631), .B(n_635), .C(n_626), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_718), .A2(n_694), .B1(n_703), .B2(n_689), .Y(n_821) );
NAND2xp67_ASAP7_75t_SL g822 ( .A(n_762), .B(n_411), .Y(n_822) );
OAI21xp5_ASAP7_75t_L g823 ( .A1(n_776), .A2(n_632), .B(n_637), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_759), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_801), .Y(n_825) );
O2A1O1Ixp5_ASAP7_75t_L g826 ( .A1(n_820), .A2(n_738), .B(n_706), .C(n_760), .Y(n_826) );
A2O1A1Ixp33_ASAP7_75t_L g827 ( .A1(n_792), .A2(n_763), .B(n_756), .C(n_765), .Y(n_827) );
OAI32xp33_ASAP7_75t_L g828 ( .A1(n_789), .A2(n_729), .A3(n_711), .B1(n_732), .B2(n_737), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_799), .B(n_709), .Y(n_829) );
AOI21xp5_ASAP7_75t_L g830 ( .A1(n_785), .A2(n_769), .B(n_766), .Y(n_830) );
AOI221x1_ASAP7_75t_L g831 ( .A1(n_811), .A2(n_761), .B1(n_747), .B2(n_751), .C(n_766), .Y(n_831) );
OAI22xp33_ASAP7_75t_L g832 ( .A1(n_783), .A2(n_721), .B1(n_722), .B2(n_734), .Y(n_832) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_808), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_803), .Y(n_834) );
AOI322xp5_ASAP7_75t_L g835 ( .A1(n_791), .A2(n_722), .A3(n_734), .B1(n_740), .B2(n_728), .C1(n_741), .C2(n_727), .Y(n_835) );
BUFx2_ASAP7_75t_SL g836 ( .A(n_788), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_782), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_783), .A2(n_740), .B1(n_764), .B2(n_728), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_790), .Y(n_839) );
OAI211xp5_ASAP7_75t_SL g840 ( .A1(n_816), .A2(n_769), .B(n_747), .C(n_751), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_781), .B(n_733), .Y(n_841) );
O2A1O1Ixp5_ASAP7_75t_L g842 ( .A1(n_795), .A2(n_777), .B(n_778), .C(n_708), .Y(n_842) );
INVx1_ASAP7_75t_SL g843 ( .A(n_796), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_784), .Y(n_844) );
AOI222xp33_ASAP7_75t_L g845 ( .A1(n_821), .A2(n_715), .B1(n_772), .B2(n_770), .C1(n_767), .C2(n_746), .Y(n_845) );
AOI211x1_ASAP7_75t_L g846 ( .A1(n_804), .A2(n_745), .B(n_714), .C(n_771), .Y(n_846) );
OAI211xp5_ASAP7_75t_L g847 ( .A1(n_798), .A2(n_774), .B(n_632), .C(n_637), .Y(n_847) );
NOR3xp33_ASAP7_75t_L g848 ( .A(n_798), .B(n_654), .C(n_688), .Y(n_848) );
AND4x1_ASAP7_75t_L g849 ( .A(n_842), .B(n_806), .C(n_823), .D(n_787), .Y(n_849) );
AOI21xp5_ASAP7_75t_L g850 ( .A1(n_827), .A2(n_824), .B(n_807), .Y(n_850) );
OAI221xp5_ASAP7_75t_L g851 ( .A1(n_827), .A2(n_806), .B1(n_786), .B2(n_818), .C(n_817), .Y(n_851) );
AOI221xp5_ASAP7_75t_L g852 ( .A1(n_833), .A2(n_797), .B1(n_793), .B2(n_802), .C(n_814), .Y(n_852) );
XNOR2xp5_ASAP7_75t_L g853 ( .A(n_836), .B(n_805), .Y(n_853) );
AND5x1_ASAP7_75t_L g854 ( .A(n_835), .B(n_822), .C(n_819), .D(n_800), .E(n_815), .Y(n_854) );
NAND4xp25_ASAP7_75t_L g855 ( .A(n_846), .B(n_810), .C(n_794), .D(n_813), .Y(n_855) );
AOI221xp5_ASAP7_75t_L g856 ( .A1(n_833), .A2(n_812), .B1(n_809), .B2(n_654), .C(n_688), .Y(n_856) );
NOR4xp25_ASAP7_75t_L g857 ( .A(n_840), .B(n_689), .C(n_679), .D(n_670), .Y(n_857) );
AOI221xp5_ASAP7_75t_L g858 ( .A1(n_832), .A2(n_679), .B1(n_670), .B2(n_667), .C(n_663), .Y(n_858) );
NOR3xp33_ASAP7_75t_L g859 ( .A(n_838), .B(n_369), .C(n_402), .Y(n_859) );
OAI32xp33_ASAP7_75t_L g860 ( .A1(n_848), .A2(n_667), .A3(n_663), .B1(n_660), .B2(n_655), .Y(n_860) );
OAI322xp33_ASAP7_75t_L g861 ( .A1(n_832), .A2(n_660), .A3(n_655), .B1(n_539), .B2(n_488), .C1(n_482), .C2(n_411), .Y(n_861) );
NAND3xp33_ASAP7_75t_L g862 ( .A(n_849), .B(n_831), .C(n_826), .Y(n_862) );
AOI211xp5_ASAP7_75t_L g863 ( .A1(n_859), .A2(n_828), .B(n_847), .C(n_829), .Y(n_863) );
OAI211xp5_ASAP7_75t_L g864 ( .A1(n_852), .A2(n_845), .B(n_829), .C(n_830), .Y(n_864) );
AND4x1_ASAP7_75t_L g865 ( .A(n_856), .B(n_837), .C(n_839), .D(n_844), .Y(n_865) );
AOI211xp5_ASAP7_75t_L g866 ( .A1(n_851), .A2(n_843), .B(n_834), .C(n_841), .Y(n_866) );
NOR2xp33_ASAP7_75t_L g867 ( .A(n_853), .B(n_825), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_855), .Y(n_868) );
NOR3x1_ASAP7_75t_L g869 ( .A(n_868), .B(n_854), .C(n_857), .Y(n_869) );
AOI211x1_ASAP7_75t_L g870 ( .A1(n_862), .A2(n_850), .B(n_860), .C(n_861), .Y(n_870) );
AOI21xp5_ASAP7_75t_L g871 ( .A1(n_867), .A2(n_864), .B(n_863), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_866), .B(n_858), .Y(n_872) );
HB1xp67_ASAP7_75t_L g873 ( .A(n_869), .Y(n_873) );
AOI221xp5_ASAP7_75t_L g874 ( .A1(n_871), .A2(n_865), .B1(n_488), .B2(n_411), .C(n_482), .Y(n_874) );
O2A1O1Ixp33_ASAP7_75t_L g875 ( .A1(n_872), .A2(n_398), .B(n_369), .C(n_358), .Y(n_875) );
NOR2x1_ASAP7_75t_L g876 ( .A(n_873), .B(n_870), .Y(n_876) );
NAND3xp33_ASAP7_75t_L g877 ( .A(n_874), .B(n_99), .C(n_100), .Y(n_877) );
INVx3_ASAP7_75t_L g878 ( .A(n_876), .Y(n_878) );
INVx1_ASAP7_75t_SL g879 ( .A(n_877), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_879), .A2(n_878), .B1(n_875), .B2(n_398), .Y(n_880) );
OAI21xp5_ASAP7_75t_SL g881 ( .A1(n_880), .A2(n_878), .B(n_103), .Y(n_881) );
AOI21xp5_ASAP7_75t_L g882 ( .A1(n_881), .A2(n_347), .B(n_402), .Y(n_882) );
OA21x2_ASAP7_75t_L g883 ( .A1(n_882), .A2(n_347), .B(n_376), .Y(n_883) );
UNKNOWN g884 ( );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_884), .A2(n_101), .B1(n_376), .B2(n_873), .Y(n_885) );
endmodule