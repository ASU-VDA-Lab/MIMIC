module real_jpeg_12026_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_263, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_263;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_139;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_0),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_0),
.A2(n_9),
.B(n_34),
.C(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_0),
.A2(n_38),
.B1(n_51),
.B2(n_52),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_0),
.B(n_39),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_0),
.B(n_49),
.C(n_52),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_0),
.B(n_65),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_0),
.B(n_31),
.C(n_35),
.Y(n_207)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_3),
.Y(n_98)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_61),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_61),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_61),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_57),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_8),
.A2(n_51),
.B1(n_52),
.B2(n_57),
.Y(n_102)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

AO22x1_ASAP7_75t_L g65 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_63),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_23)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_11),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_11),
.A2(n_28),
.B1(n_46),
.B2(n_47),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_11),
.A2(n_28),
.B1(n_51),
.B2(n_52),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_111),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_110),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_77),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_16),
.B(n_77),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_71),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_68),
.B2(n_70),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_40),
.B2(n_41),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_20),
.B(n_124),
.C(n_125),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_20),
.A2(n_21),
.B1(n_84),
.B2(n_85),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_20),
.A2(n_21),
.B1(n_124),
.B2(n_139),
.Y(n_249)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_21),
.B(n_84),
.C(n_218),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_29),
.B1(n_37),
.B2(n_39),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OA21x2_ASAP7_75t_L g68 ( 
.A1(n_23),
.A2(n_33),
.B(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_25),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_25),
.B(n_207),
.Y(n_206)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_29),
.B(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_29),
.B(n_39),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_35),
.A2(n_63),
.B(n_64),
.C(n_65),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_63),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_SL g145 ( 
.A1(n_38),
.A2(n_47),
.B(n_63),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_38),
.B(n_101),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_38),
.B(n_55),
.Y(n_188)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_42),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_68),
.C(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_42),
.A2(n_67),
.B1(n_72),
.B2(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_55),
.B(n_56),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_43),
.A2(n_55),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_44),
.A2(n_50),
.B1(n_90),
.B2(n_92),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_44),
.B(n_105),
.Y(n_104)
);

AO22x1_ASAP7_75t_SL g129 ( 
.A1(n_44),
.A2(n_50),
.B1(n_105),
.B2(n_130),
.Y(n_129)
);

NOR2x1_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_46),
.B(n_170),
.Y(n_169)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AO22x1_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_51),
.B(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_55),
.A2(n_91),
.B(n_104),
.Y(n_103)
);

OA21x2_ASAP7_75t_L g140 ( 
.A1(n_55),
.A2(n_104),
.B(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_70),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_68),
.A2(n_70),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_68),
.A2(n_70),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_70),
.B(n_124),
.C(n_212),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_70),
.B(n_228),
.C(n_233),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_72),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B(n_75),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_73),
.A2(n_75),
.B(n_87),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_73),
.A2(n_86),
.B(n_88),
.Y(n_233)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.C(n_93),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_78),
.A2(n_82),
.B1(n_83),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_84),
.B(n_89),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_89),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_84),
.A2(n_85),
.B1(n_151),
.B2(n_159),
.Y(n_150)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_85),
.B(n_152),
.C(n_155),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_106),
.B(n_107),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_95),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_103),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_96),
.A2(n_106),
.B1(n_107),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_96),
.A2(n_103),
.B1(n_106),
.B2(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_102),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_99),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_100),
.A2(n_101),
.B1(n_147),
.B2(n_156),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_101),
.A2(n_156),
.B(n_157),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_101),
.A2(n_128),
.B(n_157),
.Y(n_221)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_103),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_105),
.Y(n_213)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_131),
.B(n_260),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_113),
.B(n_116),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_123),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_117),
.A2(n_121),
.B1(n_122),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_117),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_123),
.B(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_124),
.A2(n_139),
.B1(n_140),
.B2(n_182),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_124),
.A2(n_139),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_125),
.A2(n_126),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_127),
.A2(n_129),
.B1(n_164),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_127),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_129),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_129),
.A2(n_164),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_129),
.B(n_174),
.C(n_176),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_129),
.B(n_149),
.C(n_163),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_254),
.B(n_259),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_243),
.B(n_253),
.Y(n_133)
);

OAI321xp33_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_215),
.A3(n_238),
.B1(n_241),
.B2(n_242),
.C(n_263),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_199),
.B(n_214),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_165),
.B(n_198),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_148),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_138),
.B(n_148),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.C(n_142),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_140),
.B(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_140),
.A2(n_169),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_140),
.A2(n_182),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_142),
.A2(n_143),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_146),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_160),
.B2(n_161),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_154),
.B(n_180),
.Y(n_190)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_192),
.B(n_197),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_178),
.B(n_191),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_168),
.B(n_171),
.Y(n_191)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_171)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_173),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_176),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_176),
.B(n_188),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_205),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_183),
.B(n_190),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_221),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_187),
.B(n_189),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_193),
.B(n_194),
.Y(n_197)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_200),
.B(n_201),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_208),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_204),
.C(n_208),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_224),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_224),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.C(n_223),
.Y(n_216)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_217),
.B(n_220),
.CI(n_223),
.CON(n_240),
.SN(n_240)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_237),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_234),
.B2(n_235),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_235),
.C(n_237),
.Y(n_252)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_239),
.B(n_240),
.Y(n_241)
);

BUFx24_ASAP7_75t_SL g262 ( 
.A(n_240),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_252),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_252),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_247),
.C(n_250),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_256),
.Y(n_259)
);


endmodule