module fake_jpeg_30592_n_415 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_415);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_415;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_45),
.Y(n_116)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_59),
.Y(n_93)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_17),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_53),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_15),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_13),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_67),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_58),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_18),
.B(n_13),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_21),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_71),
.Y(n_110)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_0),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_84),
.Y(n_115)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_41),
.B1(n_19),
.B2(n_30),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g96 ( 
.A(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_22),
.B(n_0),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_83),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_22),
.B(n_1),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_35),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_24),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_86),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_52),
.A2(n_20),
.B1(n_40),
.B2(n_35),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_88),
.A2(n_107),
.B1(n_54),
.B2(n_37),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_109),
.B1(n_19),
.B2(n_41),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_57),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_100),
.B(n_122),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_55),
.A2(n_20),
.B1(n_76),
.B2(n_63),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_44),
.B(n_24),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_108),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_78),
.A2(n_32),
.B1(n_29),
.B2(n_40),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_58),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_49),
.B(n_26),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_123),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_44),
.B(n_26),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_135),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_62),
.A2(n_32),
.B1(n_27),
.B2(n_28),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_126),
.A2(n_130),
.B1(n_41),
.B2(n_19),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_65),
.A2(n_32),
.B1(n_27),
.B2(n_28),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_56),
.B(n_30),
.Y(n_133)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_66),
.B(n_28),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_137),
.A2(n_144),
.B1(n_167),
.B2(n_88),
.Y(n_181)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_92),
.A2(n_85),
.B1(n_83),
.B2(n_81),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_87),
.A2(n_30),
.B1(n_20),
.B2(n_75),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_146),
.Y(n_183)
);

AO22x1_ASAP7_75t_SL g148 ( 
.A1(n_109),
.A2(n_80),
.B1(n_79),
.B2(n_77),
.Y(n_148)
);

AO22x1_ASAP7_75t_SL g175 ( 
.A1(n_148),
.A2(n_162),
.B1(n_89),
.B2(n_131),
.Y(n_175)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_89),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_96),
.A2(n_69),
.B1(n_64),
.B2(n_61),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_96),
.A2(n_32),
.B1(n_40),
.B2(n_35),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_73),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_163),
.Y(n_185)
);

INVx3_ASAP7_75t_SL g161 ( 
.A(n_95),
.Y(n_161)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_43),
.B1(n_37),
.B2(n_56),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_91),
.B(n_40),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_165),
.Y(n_182)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_102),
.B(n_2),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_115),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_102),
.A2(n_37),
.B1(n_4),
.B2(n_5),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

CKINVDCx11_ASAP7_75t_R g171 ( 
.A(n_168),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_175),
.A2(n_127),
.B1(n_169),
.B2(n_159),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_136),
.B(n_114),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_176),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_180),
.A2(n_138),
.B1(n_161),
.B2(n_127),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_181),
.B(n_187),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_147),
.A2(n_142),
.B1(n_139),
.B2(n_131),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_136),
.B(n_112),
.C(n_117),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_189),
.B(n_167),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_110),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_191),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_156),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

AOI22x1_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_162),
.B1(n_137),
.B2(n_148),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_193),
.A2(n_197),
.B1(n_199),
.B2(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_196),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_170),
.A2(n_165),
.B1(n_138),
.B2(n_107),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_195),
.A2(n_170),
.B1(n_172),
.B2(n_174),
.Y(n_219)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_148),
.B1(n_156),
.B2(n_149),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_149),
.B1(n_145),
.B2(n_162),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_143),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_206),
.Y(n_212)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_203),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_171),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_204),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_L g208 ( 
.A1(n_175),
.A2(n_146),
.B1(n_162),
.B2(n_106),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_185),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_211),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_210),
.A2(n_181),
.B1(n_144),
.B2(n_176),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_143),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_202),
.B(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_214),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_211),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_209),
.B(n_185),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_232),
.C(n_193),
.Y(n_250)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_169),
.B(n_166),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_218),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_219),
.A2(n_192),
.B1(n_199),
.B2(n_231),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_183),
.Y(n_220)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

FAx1_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_183),
.CI(n_175),
.CON(n_222),
.SN(n_222)
);

NAND2xp33_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_193),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_205),
.B(n_176),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_223),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_204),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_226),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_229),
.A2(n_200),
.B1(n_193),
.B2(n_195),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_189),
.Y(n_230)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_230),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_203),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_231),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_147),
.C(n_182),
.Y(n_232)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_206),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_250),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_210),
.B1(n_197),
.B2(n_207),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_239),
.A2(n_252),
.B1(n_228),
.B2(n_178),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_240),
.A2(n_221),
.B1(n_213),
.B2(n_201),
.Y(n_265)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_244),
.Y(n_258)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_248),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_247),
.A2(n_222),
.B(n_216),
.Y(n_254)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_249),
.A2(n_229),
.B1(n_219),
.B2(n_222),
.Y(n_262)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_251),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_224),
.A2(n_201),
.B1(n_182),
.B2(n_172),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_230),
.C(n_232),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_259),
.Y(n_293)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_224),
.B1(n_229),
.B2(n_214),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_270),
.B1(n_242),
.B2(n_251),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_249),
.B(n_235),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_256),
.A2(n_261),
.B(n_266),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_212),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_212),
.C(n_217),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_260),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_235),
.A2(n_222),
.B(n_216),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_262),
.A2(n_238),
.B1(n_239),
.B2(n_234),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_243),
.A2(n_226),
.B1(n_221),
.B2(n_222),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_264),
.A2(n_265),
.B1(n_272),
.B2(n_271),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_236),
.A2(n_228),
.B(n_184),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_217),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_238),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_244),
.A2(n_228),
.B(n_184),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_268),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_264),
.A2(n_242),
.B(n_248),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_273),
.A2(n_282),
.B(n_291),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_274),
.A2(n_277),
.B1(n_279),
.B2(n_261),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_278),
.B(n_153),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_270),
.A2(n_234),
.B1(n_237),
.B2(n_236),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_280),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_237),
.Y(n_281)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_256),
.A2(n_252),
.B(n_246),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_286),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_265),
.A2(n_245),
.B1(n_228),
.B2(n_196),
.Y(n_287)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

O2A1O1Ixp33_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_171),
.B(n_194),
.C(n_179),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_292),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_258),
.B(n_141),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_289),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_87),
.B1(n_93),
.B2(n_141),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_272),
.A2(n_178),
.B(n_203),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_161),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_281),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_296),
.B(n_299),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_260),
.B1(n_271),
.B2(n_255),
.Y(n_298)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_298),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_311),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_274),
.A2(n_253),
.B1(n_254),
.B2(n_259),
.Y(n_303)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_303),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_279),
.A2(n_267),
.B1(n_263),
.B2(n_174),
.Y(n_304)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_304),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_293),
.B(n_263),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_308),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_174),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_277),
.A2(n_275),
.B1(n_294),
.B2(n_276),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_309),
.A2(n_276),
.B1(n_287),
.B2(n_284),
.Y(n_321)
);

OA22x2_ASAP7_75t_L g310 ( 
.A1(n_275),
.A2(n_179),
.B1(n_186),
.B2(n_177),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_310),
.A2(n_121),
.B1(n_119),
.B2(n_90),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_186),
.C(n_164),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_284),
.C(n_291),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_168),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_316),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_273),
.B(n_157),
.Y(n_316)
);

NAND2xp33_ASAP7_75t_SL g322 ( 
.A(n_317),
.B(n_280),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_321),
.A2(n_334),
.B1(n_297),
.B2(n_312),
.Y(n_342)
);

XNOR2x1_ASAP7_75t_L g354 ( 
.A(n_322),
.B(n_327),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_315),
.A2(n_286),
.B(n_283),
.Y(n_323)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_309),
.A2(n_288),
.B(n_140),
.Y(n_328)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_328),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_315),
.A2(n_94),
.B(n_98),
.Y(n_329)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_329),
.Y(n_351)
);

NOR2xp67_ASAP7_75t_SL g330 ( 
.A(n_313),
.B(n_150),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_330),
.B(n_331),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_125),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_158),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_332),
.A2(n_337),
.B1(n_132),
.B2(n_106),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_306),
.A2(n_90),
.B1(n_121),
.B2(n_119),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_155),
.C(n_98),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_338),
.C(n_340),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_95),
.C(n_105),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_301),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_339),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_300),
.B(n_103),
.C(n_105),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_342),
.A2(n_337),
.B1(n_111),
.B2(n_116),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_300),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_347),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_306),
.C(n_312),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_346),
.B(n_349),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_311),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_325),
.A2(n_295),
.B1(n_318),
.B2(n_317),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_335),
.Y(n_352)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_352),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_310),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_355),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_310),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_356),
.A2(n_334),
.B1(n_336),
.B2(n_338),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_324),
.A2(n_310),
.B1(n_111),
.B2(n_125),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_358),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_326),
.C(n_333),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_326),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_360),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_358),
.B(n_340),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_362),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_354),
.B(n_322),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_345),
.A2(n_354),
.B(n_351),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_365),
.A2(n_355),
.B(n_350),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_348),
.Y(n_368)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_368),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_369),
.B(n_371),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_343),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_346),
.A2(n_103),
.B1(n_120),
.B2(n_128),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_128),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_341),
.C(n_353),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_373),
.B(n_383),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_370),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_377),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_347),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_376),
.B(n_37),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_366),
.B(n_341),
.Y(n_377)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_378),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_364),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_382),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_362),
.B(n_120),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_381),
.B(n_367),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_385),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_374),
.A2(n_367),
.B1(n_366),
.B2(n_369),
.Y(n_386)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_386),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_387),
.B(n_5),
.C(n_6),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_384),
.B(n_3),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_389),
.A2(n_391),
.B(n_392),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_379),
.B(n_3),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_375),
.A2(n_37),
.B(n_4),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_393),
.A2(n_386),
.B1(n_390),
.B2(n_380),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_396),
.B(n_401),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_394),
.A2(n_376),
.B(n_4),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_399),
.A2(n_6),
.B(n_7),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_388),
.A2(n_3),
.B(n_4),
.Y(n_400)
);

AOI21x1_ASAP7_75t_L g404 ( 
.A1(n_400),
.A2(n_6),
.B(n_7),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_395),
.B(n_387),
.C(n_7),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_402),
.B(n_403),
.Y(n_408)
);

AO221x1_ASAP7_75t_L g407 ( 
.A1(n_404),
.A2(n_398),
.B1(n_397),
.B2(n_10),
.C(n_11),
.Y(n_407)
);

OAI21x1_ASAP7_75t_SL g405 ( 
.A1(n_396),
.A2(n_8),
.B(n_9),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_405),
.A2(n_8),
.B(n_9),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_407),
.A2(n_408),
.B(n_406),
.Y(n_410)
);

NAND3xp33_ASAP7_75t_L g411 ( 
.A(n_409),
.B(n_8),
.C(n_9),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_410),
.B(n_411),
.C(n_8),
.Y(n_412)
);

BUFx24_ASAP7_75t_SL g413 ( 
.A(n_412),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_413),
.A2(n_10),
.B(n_11),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_414),
.A2(n_10),
.B(n_407),
.Y(n_415)
);


endmodule