module fake_jpeg_3163_n_649 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_649);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_649;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_15),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_8),
.B(n_14),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_58),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_60),
.Y(n_166)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_61),
.Y(n_149)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_62),
.Y(n_179)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_63),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_65),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_34),
.A2(n_9),
.B(n_1),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_66),
.B(n_97),
.Y(n_154)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_68),
.Y(n_176)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_69),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_70),
.Y(n_171)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_73),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_74),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_75),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_76),
.Y(n_210)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_78),
.Y(n_196)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_79),
.Y(n_178)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_80),
.Y(n_222)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_81),
.Y(n_180)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_82),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_86),
.Y(n_202)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_87),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_89),
.Y(n_187)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_90),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_91),
.Y(n_207)
);

BUFx8_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_92),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_93),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_94),
.Y(n_217)
);

CKINVDCx9p33_ASAP7_75t_R g95 ( 
.A(n_43),
.Y(n_95)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_34),
.B(n_9),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_35),
.B(n_11),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_98),
.B(n_119),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_99),
.Y(n_133)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_100),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_101),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_103),
.Y(n_219)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_105),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_35),
.B(n_8),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_27),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_109),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_110),
.Y(n_211)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_112),
.Y(n_223)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_113),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_21),
.Y(n_114)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_114),
.Y(n_225)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_24),
.Y(n_115)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_24),
.Y(n_116)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_116),
.Y(n_228)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_28),
.Y(n_117)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_28),
.Y(n_118)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_31),
.B(n_19),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_25),
.Y(n_120)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_21),
.Y(n_123)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_25),
.Y(n_124)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_40),
.Y(n_125)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_125),
.Y(n_200)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_40),
.Y(n_126)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_126),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_40),
.Y(n_127)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_127),
.Y(n_213)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_37),
.Y(n_128)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_129),
.Y(n_226)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_36),
.Y(n_130)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_97),
.B(n_37),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_139),
.B(n_155),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_44),
.B1(n_55),
.B2(n_48),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_143),
.A2(n_147),
.B1(n_0),
.B2(n_1),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_92),
.A2(n_42),
.B1(n_27),
.B2(n_38),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_146),
.A2(n_184),
.B1(n_188),
.B2(n_93),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_42),
.B1(n_27),
.B2(n_38),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_129),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_153),
.B(n_201),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_125),
.B(n_55),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_156),
.B(n_164),
.Y(n_261)
);

INVx6_ASAP7_75t_SL g157 ( 
.A(n_101),
.Y(n_157)
);

INVx13_ASAP7_75t_L g278 ( 
.A(n_157),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_123),
.A2(n_57),
.B1(n_33),
.B2(n_39),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_161),
.B(n_99),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_65),
.B(n_33),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_126),
.A2(n_54),
.B1(n_26),
.B2(n_57),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_173),
.A2(n_197),
.B1(n_206),
.B2(n_94),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_73),
.B(n_45),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_181),
.B(n_183),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_127),
.B(n_44),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_182),
.B(n_218),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_80),
.B(n_48),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_77),
.A2(n_42),
.B1(n_31),
.B2(n_51),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_82),
.B(n_45),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_185),
.B(n_193),
.Y(n_274)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_100),
.Y(n_186)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_89),
.A2(n_42),
.B1(n_51),
.B2(n_39),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_113),
.B(n_26),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_59),
.A2(n_54),
.B1(n_43),
.B2(n_56),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_60),
.Y(n_199)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_199),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_121),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_70),
.Y(n_205)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_108),
.A2(n_43),
.B1(n_56),
.B2(n_2),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_75),
.B(n_12),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_208),
.B(n_216),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_76),
.B(n_12),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_83),
.B(n_106),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_84),
.B(n_43),
.C(n_56),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_220),
.B(n_0),
.C(n_4),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_164),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_230),
.B(n_231),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_181),
.Y(n_231)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_145),
.Y(n_233)
);

INVx3_ASAP7_75t_SL g342 ( 
.A(n_233),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_234),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_236),
.A2(n_311),
.B1(n_217),
.B2(n_215),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_165),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_237),
.B(n_260),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_145),
.Y(n_239)
);

INVx5_ASAP7_75t_L g357 ( 
.A(n_239),
.Y(n_357)
);

O2A1O1Ixp33_ASAP7_75t_SL g240 ( 
.A1(n_154),
.A2(n_43),
.B(n_91),
.C(n_88),
.Y(n_240)
);

O2A1O1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_240),
.A2(n_296),
.B(n_234),
.C(n_269),
.Y(n_344)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_242),
.Y(n_320)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_243),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_244),
.Y(n_316)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_166),
.Y(n_246)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_246),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_177),
.Y(n_247)
);

BUFx2_ASAP7_75t_SL g366 ( 
.A(n_247),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_248),
.A2(n_211),
.B1(n_198),
.B2(n_195),
.Y(n_321)
);

BUFx8_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_249),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_165),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_250),
.Y(n_372)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_131),
.Y(n_251)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_251),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_166),
.Y(n_252)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_252),
.Y(n_354)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_254),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_185),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_255),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_171),
.Y(n_256)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_256),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_156),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_257),
.B(n_267),
.Y(n_314)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_135),
.Y(n_258)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_258),
.Y(n_327)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_140),
.Y(n_259)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_259),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_193),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_132),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_263)
);

OAI22x1_ASAP7_75t_L g368 ( 
.A1(n_263),
.A2(n_269),
.B1(n_277),
.B2(n_6),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_174),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_264),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_154),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_265),
.A2(n_300),
.B(n_190),
.Y(n_352)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_168),
.Y(n_266)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_266),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_179),
.B(n_13),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_159),
.B(n_19),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_268),
.B(n_287),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_146),
.A2(n_142),
.B1(n_174),
.B2(n_138),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_158),
.Y(n_270)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_270),
.Y(n_334)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_167),
.Y(n_271)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_271),
.Y(n_348)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_149),
.Y(n_272)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_272),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_226),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_273),
.B(n_281),
.Y(n_335)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_169),
.Y(n_275)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_275),
.Y(n_351)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_171),
.Y(n_276)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_276),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_192),
.A2(n_12),
.B1(n_4),
.B2(n_5),
.Y(n_277)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_151),
.Y(n_279)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_279),
.Y(n_365)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_228),
.Y(n_280)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_280),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_209),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_172),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_282),
.B(n_283),
.Y(n_359)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_187),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_163),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_285),
.B(n_286),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_196),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_202),
.B(n_14),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_214),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_288),
.B(n_289),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_175),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_178),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_290),
.B(n_292),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_204),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_291),
.Y(n_347)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_180),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_200),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_293),
.B(n_294),
.Y(n_338)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_189),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_194),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_301),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_296),
.B(n_147),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_160),
.B(n_15),
.Y(n_297)
);

INVx3_ASAP7_75t_SL g298 ( 
.A(n_191),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_224),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_208),
.A2(n_15),
.B1(n_5),
.B2(n_6),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_204),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_219),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_303),
.Y(n_332)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_175),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_176),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_304),
.B(n_305),
.Y(n_356)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_212),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_133),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_306),
.B(n_307),
.Y(n_360)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_226),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_182),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_308),
.A2(n_262),
.B1(n_232),
.B2(n_274),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_210),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_309),
.A2(n_312),
.B1(n_313),
.B2(n_150),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_141),
.B(n_5),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_310),
.B(n_190),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_133),
.A2(n_222),
.B1(n_213),
.B2(n_210),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_222),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_134),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_257),
.B(n_261),
.C(n_255),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_315),
.B(n_345),
.C(n_299),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_321),
.A2(n_329),
.B1(n_337),
.B2(n_264),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_322),
.B(n_265),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_244),
.A2(n_184),
.B(n_188),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_325),
.A2(n_370),
.B(n_263),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_326),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_330),
.B(n_361),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_236),
.A2(n_217),
.B1(n_215),
.B2(n_207),
.Y(n_337)
);

O2A1O1Ixp33_ASAP7_75t_L g402 ( 
.A1(n_344),
.A2(n_278),
.B(n_298),
.C(n_301),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_284),
.B(n_190),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_248),
.A2(n_170),
.B1(n_152),
.B2(n_207),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_346),
.A2(n_358),
.B1(n_362),
.B2(n_252),
.Y(n_405)
);

AOI21xp33_ASAP7_75t_L g395 ( 
.A1(n_352),
.A2(n_311),
.B(n_313),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_240),
.A2(n_134),
.B1(n_137),
.B2(n_136),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_229),
.A2(n_137),
.B1(n_136),
.B2(n_148),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_238),
.A2(n_144),
.B1(n_162),
.B2(n_0),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_363),
.A2(n_250),
.B1(n_270),
.B2(n_304),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_367),
.B(n_254),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_368),
.A2(n_277),
.B1(n_303),
.B2(n_289),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_249),
.A2(n_7),
.B(n_16),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_335),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_374),
.B(n_384),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_375),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_376),
.B(n_381),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_322),
.B(n_300),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_377),
.B(n_398),
.Y(n_423)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_318),
.Y(n_378)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_378),
.Y(n_425)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_364),
.Y(n_379)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_379),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_323),
.B(n_253),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_380),
.B(n_392),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_345),
.B(n_235),
.C(n_241),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_382),
.B(n_388),
.C(n_415),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_316),
.A2(n_283),
.B1(n_282),
.B2(n_275),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_383),
.A2(n_385),
.B1(n_393),
.B2(n_397),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_340),
.B(n_249),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_318),
.Y(n_386)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_386),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_338),
.Y(n_387)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_387),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_315),
.B(n_286),
.C(n_293),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_328),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_389),
.B(n_407),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_342),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_390),
.Y(n_448)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_391),
.Y(n_440)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_360),
.Y(n_394)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_394),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_395),
.A2(n_396),
.B(n_411),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_353),
.B(n_288),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_330),
.B(n_276),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_358),
.A2(n_233),
.B1(n_309),
.B2(n_256),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_400),
.A2(n_403),
.B1(n_410),
.B2(n_371),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_314),
.B(n_246),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_401),
.B(n_404),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_402),
.A2(n_416),
.B(n_418),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_316),
.A2(n_325),
.B1(n_344),
.B2(n_346),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_314),
.B(n_239),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_405),
.A2(n_357),
.B1(n_369),
.B2(n_365),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_323),
.B(n_291),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_406),
.B(n_408),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_355),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_332),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_373),
.B(n_7),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_409),
.B(n_413),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_321),
.A2(n_278),
.B1(n_16),
.B2(n_18),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_368),
.A2(n_7),
.B1(n_16),
.B2(n_18),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_353),
.B(n_19),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_412),
.A2(n_419),
.B(n_420),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_373),
.B(n_317),
.Y(n_413)
);

MAJx2_ASAP7_75t_L g414 ( 
.A(n_352),
.B(n_327),
.C(n_348),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_414),
.B(n_421),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_327),
.B(n_362),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_349),
.A2(n_338),
.B(n_356),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_332),
.B(n_356),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_417),
.B(n_391),
.Y(n_456)
);

FAx1_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_361),
.CI(n_359),
.CON(n_418),
.SN(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_359),
.A2(n_334),
.B(n_351),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_359),
.A2(n_342),
.B1(n_347),
.B2(n_351),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_396),
.A2(n_347),
.B1(n_342),
.B2(n_334),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_424),
.A2(n_450),
.B(n_458),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_419),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_427),
.B(n_456),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_403),
.A2(n_364),
.B1(n_348),
.B2(n_324),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_429),
.A2(n_438),
.B1(n_441),
.B2(n_442),
.Y(n_490)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_379),
.Y(n_436)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_436),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_415),
.A2(n_324),
.B1(n_354),
.B2(n_339),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_408),
.A2(n_354),
.B1(n_339),
.B2(n_369),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_443),
.A2(n_405),
.B1(n_396),
.B2(n_387),
.Y(n_469)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_378),
.Y(n_447)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_447),
.Y(n_463)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_386),
.Y(n_449)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_449),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_375),
.A2(n_336),
.B(n_331),
.Y(n_450)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_417),
.Y(n_453)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_453),
.Y(n_482)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_406),
.Y(n_455)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_455),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_418),
.A2(n_331),
.B(n_333),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_394),
.A2(n_357),
.B1(n_350),
.B2(n_365),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_459),
.A2(n_385),
.B1(n_400),
.B2(n_389),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_381),
.B(n_350),
.C(n_333),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_461),
.C(n_437),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_382),
.B(n_319),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_420),
.Y(n_462)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_462),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_464),
.B(n_483),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_453),
.A2(n_398),
.B1(n_418),
.B2(n_393),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_465),
.A2(n_488),
.B1(n_455),
.B2(n_428),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_413),
.Y(n_466)
);

NAND3xp33_ASAP7_75t_L g524 ( 
.A(n_466),
.B(n_472),
.C(n_486),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_432),
.A2(n_418),
.B(n_402),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_467),
.A2(n_487),
.B(n_499),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_469),
.A2(n_473),
.B1(n_478),
.B2(n_494),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_451),
.A2(n_407),
.B1(n_416),
.B2(n_414),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g525 ( 
.A(n_471),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_434),
.B(n_422),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_443),
.A2(n_401),
.B1(n_421),
.B2(n_377),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_404),
.Y(n_474)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_474),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_431),
.B(n_388),
.Y(n_475)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_475),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_437),
.B(n_414),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_476),
.B(n_477),
.C(n_480),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_462),
.A2(n_376),
.B1(n_392),
.B2(n_412),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_446),
.B(n_380),
.C(n_412),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_457),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_481),
.B(n_492),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_458),
.Y(n_483)
);

AND2x6_ASAP7_75t_L g484 ( 
.A(n_432),
.B(n_402),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_484),
.B(n_489),
.Y(n_508)
);

OAI22x1_ASAP7_75t_L g485 ( 
.A1(n_435),
.A2(n_411),
.B1(n_410),
.B2(n_390),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_485),
.A2(n_444),
.B(n_429),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_434),
.B(n_409),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_435),
.A2(n_384),
.B(n_399),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_440),
.A2(n_390),
.B1(n_319),
.B2(n_343),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_438),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_431),
.B(n_320),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_436),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_459),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_446),
.B(n_423),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_477),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_426),
.A2(n_320),
.B1(n_343),
.B2(n_341),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_439),
.B(n_366),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_497),
.B(n_460),
.C(n_433),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_450),
.A2(n_341),
.B(n_372),
.Y(n_499)
);

A2O1A1O1Ixp25_ASAP7_75t_L g500 ( 
.A1(n_423),
.A2(n_439),
.B(n_433),
.C(n_445),
.D(n_440),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_500),
.A2(n_441),
.B(n_452),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_491),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_502),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_476),
.B(n_461),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_503),
.B(n_514),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_479),
.A2(n_426),
.B(n_444),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g550 ( 
.A1(n_505),
.A2(n_513),
.B(n_519),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_482),
.B(n_445),
.Y(n_509)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_509),
.Y(n_539)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_510),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_511),
.B(n_498),
.C(n_478),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_482),
.A2(n_447),
.B1(n_449),
.B2(n_425),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_516),
.A2(n_518),
.B1(n_526),
.B2(n_529),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_496),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_517),
.B(n_496),
.Y(n_560)
);

CKINVDCx14_ASAP7_75t_R g518 ( 
.A(n_487),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_467),
.A2(n_427),
.B(n_430),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_468),
.B(n_430),
.Y(n_520)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_520),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_468),
.B(n_425),
.Y(n_522)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_522),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_499),
.Y(n_523)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_523),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_488),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_527),
.A2(n_463),
.B1(n_470),
.B2(n_500),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_479),
.Y(n_528)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_528),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_495),
.B(n_428),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_495),
.B(n_452),
.Y(n_530)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_530),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_493),
.B(n_424),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_531),
.B(n_532),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_497),
.B(n_475),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_533),
.A2(n_494),
.B1(n_489),
.B2(n_498),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_480),
.B(n_448),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_534),
.B(n_465),
.Y(n_542)
);

CKINVDCx16_ASAP7_75t_R g535 ( 
.A(n_469),
.Y(n_535)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_535),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_511),
.B(n_532),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_537),
.B(n_541),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_534),
.B(n_473),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_SL g582 ( 
.A(n_542),
.B(n_515),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_543),
.B(n_556),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_521),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g571 ( 
.A(n_544),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_503),
.B(n_483),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_547),
.B(n_531),
.Y(n_585)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_509),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_552),
.B(n_553),
.Y(n_580)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_520),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_522),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_554),
.A2(n_557),
.B1(n_561),
.B2(n_562),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_514),
.B(n_474),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_559),
.A2(n_533),
.B1(n_504),
.B2(n_513),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_560),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_515),
.A2(n_490),
.B1(n_464),
.B2(n_485),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_524),
.A2(n_463),
.B1(n_470),
.B2(n_484),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_564),
.A2(n_574),
.B1(n_551),
.B2(n_554),
.Y(n_595)
);

CKINVDCx14_ASAP7_75t_R g566 ( 
.A(n_538),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_566),
.B(n_567),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_537),
.B(n_506),
.C(n_512),
.Y(n_567)
);

BUFx24_ASAP7_75t_SL g569 ( 
.A(n_556),
.Y(n_569)
);

BUFx24_ASAP7_75t_SL g604 ( 
.A(n_569),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_543),
.B(n_506),
.C(n_512),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_570),
.B(n_586),
.C(n_540),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_561),
.A2(n_527),
.B1(n_525),
.B2(n_535),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_573),
.A2(n_575),
.B1(n_576),
.B2(n_581),
.Y(n_597)
);

CKINVDCx14_ASAP7_75t_R g574 ( 
.A(n_550),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_563),
.A2(n_548),
.B1(n_546),
.B2(n_553),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_546),
.A2(n_504),
.B1(n_508),
.B2(n_502),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_550),
.A2(n_508),
.B(n_528),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_577),
.B(n_584),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_555),
.B(n_523),
.Y(n_578)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_578),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_539),
.A2(n_501),
.B1(n_526),
.B2(n_529),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_SL g599 ( 
.A(n_582),
.B(n_585),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_548),
.A2(n_501),
.B1(n_519),
.B2(n_505),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_583),
.A2(n_549),
.B1(n_510),
.B2(n_530),
.Y(n_602)
);

CKINVDCx16_ASAP7_75t_R g584 ( 
.A(n_559),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_536),
.B(n_507),
.C(n_516),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_568),
.B(n_542),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_588),
.B(n_589),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_568),
.B(n_540),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_572),
.Y(n_590)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_590),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_591),
.B(n_592),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_571),
.B(n_541),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_570),
.B(n_536),
.C(n_558),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_593),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_567),
.B(n_547),
.C(n_551),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_594),
.B(n_598),
.C(n_600),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_SL g616 ( 
.A1(n_595),
.A2(n_575),
.B1(n_578),
.B2(n_517),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_579),
.B(n_552),
.C(n_549),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_579),
.B(n_560),
.C(n_507),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_586),
.B(n_545),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_601),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_602),
.A2(n_564),
.B1(n_580),
.B2(n_565),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_585),
.B(n_560),
.Y(n_605)
);

MAJx2_ASAP7_75t_L g614 ( 
.A(n_605),
.B(n_578),
.C(n_573),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_596),
.A2(n_577),
.B(n_580),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_SL g628 ( 
.A(n_606),
.B(n_372),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_593),
.B(n_582),
.C(n_565),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_609),
.B(n_618),
.C(n_611),
.Y(n_631)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_613),
.Y(n_625)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_614),
.B(n_599),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_587),
.A2(n_576),
.B(n_583),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_615),
.B(n_616),
.Y(n_621)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_603),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_617),
.B(n_619),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_591),
.B(n_517),
.C(n_448),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_597),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_SL g622 ( 
.A1(n_615),
.A2(n_590),
.B1(n_598),
.B2(n_594),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_622),
.B(n_624),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_616),
.A2(n_605),
.B1(n_588),
.B2(n_589),
.Y(n_623)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_623),
.Y(n_634)
);

INVx11_ASAP7_75t_L g624 ( 
.A(n_618),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_613),
.A2(n_599),
.B(n_604),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_626),
.A2(n_628),
.B(n_609),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_627),
.B(n_630),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_607),
.A2(n_620),
.B1(n_608),
.B2(n_612),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_631),
.B(n_610),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_632),
.B(n_622),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_SL g636 ( 
.A1(n_626),
.A2(n_612),
.B(n_608),
.Y(n_636)
);

AOI21xp33_ASAP7_75t_L g642 ( 
.A1(n_636),
.A2(n_638),
.B(n_625),
.Y(n_642)
);

OAI21x1_ASAP7_75t_L g639 ( 
.A1(n_637),
.A2(n_621),
.B(n_628),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_625),
.B(n_614),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_639),
.B(n_640),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_633),
.B(n_629),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_SL g643 ( 
.A1(n_641),
.A2(n_642),
.B(n_635),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_643),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_645),
.B(n_644),
.C(n_634),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g647 ( 
.A1(n_646),
.A2(n_638),
.B(n_621),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_647),
.B(n_631),
.C(n_627),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_648),
.A2(n_624),
.B(n_611),
.Y(n_649)
);


endmodule