module fake_jpeg_19871_n_355 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_355);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_55),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_19),
.B1(n_34),
.B2(n_28),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_61),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_33),
.B1(n_18),
.B2(n_20),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_59),
.A2(n_71),
.B1(n_86),
.B2(n_25),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_20),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_19),
.B1(n_34),
.B2(n_28),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_62),
.A2(n_82),
.B1(n_54),
.B2(n_17),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_65),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_35),
.B1(n_24),
.B2(n_29),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_43),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_37),
.B(n_25),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_69),
.B(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_73),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_28),
.B1(n_34),
.B2(n_27),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_16),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_23),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_27),
.B1(n_32),
.B2(n_23),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_35),
.B1(n_29),
.B2(n_31),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_43),
.B(n_17),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_30),
.Y(n_127)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_94),
.A2(n_121),
.B1(n_68),
.B2(n_1),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_32),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_97),
.B(n_103),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_64),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_100),
.B(n_108),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_66),
.B(n_32),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_103),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_67),
.B(n_17),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_16),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_105),
.B(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_25),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_107),
.A2(n_115),
.B1(n_7),
.B2(n_14),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_65),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_56),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_111),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_40),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_122),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_82),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_23),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_125),
.Y(n_149)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_83),
.B(n_38),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_129),
.C(n_52),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_72),
.A2(n_29),
.B1(n_35),
.B2(n_31),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_62),
.A2(n_40),
.B1(n_38),
.B2(n_31),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_46),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_84),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_128),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_68),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_52),
.C(n_50),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_124),
.A2(n_78),
.B1(n_81),
.B2(n_80),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_132),
.A2(n_160),
.B1(n_118),
.B2(n_128),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_133),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_139),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_81),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_79),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_142),
.B(n_118),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_93),
.B(n_87),
.C(n_50),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_148),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_30),
.Y(n_148)
);

AO22x2_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_68),
.B1(n_1),
.B2(n_2),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_150),
.B(n_0),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_112),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_151),
.B(n_157),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_30),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_158),
.Y(n_185)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_91),
.B(n_7),
.Y(n_157)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_126),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_108),
.B1(n_124),
.B2(n_110),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_163),
.A2(n_164),
.B1(n_173),
.B2(n_177),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_144),
.A2(n_104),
.B1(n_97),
.B2(n_94),
.Y(n_164)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_167),
.B(n_168),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_96),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_159),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_170),
.B(n_174),
.Y(n_224)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_121),
.B1(n_94),
.B2(n_129),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_95),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_134),
.A2(n_100),
.B1(n_109),
.B2(n_113),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_134),
.A2(n_145),
.B1(n_154),
.B2(n_150),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_142),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_183),
.B1(n_186),
.B2(n_190),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_95),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_181),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_125),
.B1(n_123),
.B2(n_101),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_139),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_188),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_133),
.A2(n_101),
.B1(n_117),
.B2(n_92),
.Y(n_186)
);

AND2x4_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_126),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_140),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_143),
.B(n_116),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_131),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_132),
.A2(n_6),
.B1(n_14),
.B2(n_12),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_197),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_155),
.A2(n_12),
.B1(n_10),
.B2(n_9),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_116),
.B1(n_1),
.B2(n_2),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_150),
.B(n_156),
.Y(n_216)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_131),
.Y(n_196)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_137),
.A2(n_116),
.B1(n_3),
.B2(n_4),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_223),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_169),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_200),
.B(n_203),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_146),
.C(n_143),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_229),
.C(n_230),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_196),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_171),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_205),
.B(n_213),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_162),
.B(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_206),
.B(n_210),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_148),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_212),
.A2(n_220),
.B(n_0),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_172),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_150),
.B(n_135),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_215),
.A2(n_216),
.B(n_187),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_135),
.Y(n_218)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_141),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_141),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_187),
.Y(n_227)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

INVx13_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_152),
.C(n_136),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_136),
.Y(n_230)
);

AOI32xp33_ASAP7_75t_SL g269 ( 
.A1(n_232),
.A2(n_233),
.A3(n_209),
.B1(n_222),
.B2(n_217),
.Y(n_269)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_187),
.B(n_195),
.Y(n_233)
);

A2O1A1O1Ixp25_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_180),
.B(n_185),
.C(n_165),
.D(n_164),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_225),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_227),
.A2(n_179),
.B1(n_173),
.B2(n_183),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_240),
.B1(n_249),
.B2(n_255),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_227),
.A2(n_184),
.B1(n_163),
.B2(n_192),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_204),
.A2(n_185),
.B1(n_165),
.B2(n_194),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_241),
.A2(n_242),
.B1(n_244),
.B2(n_211),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_212),
.A2(n_185),
.B1(n_165),
.B2(n_167),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_212),
.A2(n_161),
.B1(n_189),
.B2(n_6),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_254),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_226),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_217),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_222),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_202),
.A2(n_3),
.B(n_5),
.C(n_9),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_226),
.A2(n_231),
.B1(n_206),
.B2(n_214),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_207),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_256),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_10),
.B1(n_3),
.B2(n_5),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_257),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_214),
.A2(n_10),
.B1(n_220),
.B2(n_211),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_207),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_259),
.Y(n_275)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_237),
.Y(n_291)
);

OAI22x1_ASAP7_75t_L g263 ( 
.A1(n_233),
.A2(n_220),
.B1(n_224),
.B2(n_208),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_263),
.A2(n_240),
.B(n_241),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_223),
.C(n_199),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_270),
.C(n_276),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_253),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_267),
.B(n_272),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_263),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_230),
.C(n_201),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_252),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_243),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_278),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_235),
.B(n_210),
.C(n_209),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_281),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_245),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_244),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_249),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_235),
.B(n_198),
.C(n_221),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_281),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_198),
.C(n_221),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_284),
.A2(n_288),
.B(n_296),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_280),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_282),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_293),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_291),
.A2(n_299),
.B1(n_301),
.B2(n_260),
.Y(n_309)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_272),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_264),
.Y(n_294)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_269),
.A2(n_246),
.B(n_232),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_250),
.Y(n_298)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_298),
.Y(n_314)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_265),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_300),
.Y(n_304)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_265),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_268),
.C(n_277),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_303),
.A2(n_288),
.B(n_273),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_270),
.C(n_266),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_307),
.C(n_312),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_315),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_287),
.C(n_276),
.Y(n_307)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_309),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_262),
.C(n_255),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_290),
.Y(n_313)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_285),
.B(n_250),
.C(n_233),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_317),
.A2(n_324),
.B(n_258),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_302),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_323),
.Y(n_330)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_288),
.B(n_273),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_325),
.B(n_326),
.Y(n_334)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_310),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_311),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_289),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_268),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_328),
.A2(n_296),
.B1(n_284),
.B2(n_316),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_329),
.B(n_337),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_307),
.C(n_305),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_331),
.B(n_332),
.C(n_336),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_306),
.C(n_312),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_333),
.A2(n_321),
.B(n_328),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_318),
.A2(n_304),
.B1(n_301),
.B2(n_300),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_335),
.A2(n_291),
.B1(n_271),
.B2(n_275),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_315),
.C(n_314),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_331),
.B(n_297),
.Y(n_338)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_338),
.Y(n_345)
);

OA21x2_ASAP7_75t_L g348 ( 
.A1(n_341),
.A2(n_342),
.B(n_344),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_330),
.A2(n_319),
.B(n_322),
.Y(n_342)
);

OAI21x1_ASAP7_75t_L g343 ( 
.A1(n_336),
.A2(n_248),
.B(n_275),
.Y(n_343)
);

AO21x1_ASAP7_75t_L g347 ( 
.A1(n_343),
.A2(n_236),
.B(n_271),
.Y(n_347)
);

AOI21xp33_ASAP7_75t_L g346 ( 
.A1(n_340),
.A2(n_292),
.B(n_334),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_346),
.A2(n_254),
.B(n_247),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_347),
.A2(n_340),
.B(n_335),
.Y(n_349)
);

AOI21x1_ASAP7_75t_L g351 ( 
.A1(n_349),
.A2(n_350),
.B(n_348),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_345),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_339),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_239),
.C(n_339),
.Y(n_354)
);

BUFx24_ASAP7_75t_SL g355 ( 
.A(n_354),
.Y(n_355)
);


endmodule