module fake_jpeg_3921_n_289 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_289);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_1),
.B(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_13),
.B1(n_26),
.B2(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_15),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_50),
.B1(n_26),
.B2(n_27),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_37),
.B1(n_32),
.B2(n_23),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_23),
.B1(n_13),
.B2(n_27),
.Y(n_54)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_23),
.B1(n_27),
.B2(n_13),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_57),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_58),
.B1(n_61),
.B2(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_42),
.B1(n_26),
.B2(n_15),
.Y(n_73)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_30),
.B1(n_36),
.B2(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_59),
.B(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_40),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_65),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_34),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_62),
.B(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_31),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_36),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_33),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_18),
.C(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_31),
.C(n_28),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_78),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_68),
.B1(n_46),
.B2(n_55),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_86),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_65),
.A2(n_44),
.B1(n_39),
.B2(n_48),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_83),
.B1(n_53),
.B2(n_52),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_39),
.B1(n_42),
.B2(n_46),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_59),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_42),
.B1(n_46),
.B2(n_49),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_52),
.B1(n_57),
.B2(n_60),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_31),
.C(n_28),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_89),
.Y(n_91)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_65),
.B1(n_66),
.B2(n_58),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_92),
.B1(n_99),
.B2(n_104),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_66),
.B1(n_54),
.B2(n_67),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_100),
.B1(n_29),
.B2(n_14),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_18),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_55),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_101),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_36),
.B(n_33),
.C(n_21),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_53),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_20),
.B(n_16),
.Y(n_130)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_29),
.B1(n_31),
.B2(n_28),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_105),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g106 ( 
.A1(n_71),
.A2(n_29),
.B(n_31),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_106),
.A2(n_75),
.B(n_71),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_79),
.B(n_25),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_28),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_104),
.A2(n_70),
.B1(n_82),
.B2(n_83),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_125),
.B1(n_111),
.B2(n_123),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_70),
.C(n_88),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_120),
.C(n_113),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_71),
.B1(n_81),
.B2(n_88),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_124),
.B1(n_99),
.B2(n_28),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_71),
.B(n_79),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_109),
.B(n_94),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_129),
.B(n_130),
.Y(n_142)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_78),
.C(n_85),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_85),
.B1(n_87),
.B2(n_60),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_21),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_141),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_132),
.A2(n_139),
.B1(n_143),
.B2(n_124),
.Y(n_170)
);

AOI22x1_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_99),
.B1(n_102),
.B2(n_90),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_154),
.B(n_152),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_134),
.A2(n_136),
.B(n_150),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_125),
.Y(n_165)
);

OA21x2_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_111),
.B(n_129),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_99),
.B1(n_103),
.B2(n_96),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_115),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_99),
.B1(n_95),
.B2(n_105),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_99),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_147),
.C(n_151),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_128),
.B(n_16),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_25),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_121),
.B(n_127),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_113),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_19),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_11),
.B(n_12),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_84),
.C(n_80),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_20),
.B(n_16),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_152),
.A2(n_130),
.B(n_129),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_110),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_154),
.C(n_120),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_14),
.C(n_25),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_137),
.B(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_160),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_131),
.B(n_118),
.Y(n_162)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_164),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_146),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_165),
.A2(n_170),
.B1(n_178),
.B2(n_138),
.Y(n_181)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_19),
.C(n_25),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_172),
.B(n_142),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_173),
.A2(n_174),
.B1(n_179),
.B2(n_142),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_133),
.A2(n_128),
.B1(n_25),
.B2(n_14),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_176),
.Y(n_188)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_135),
.A2(n_21),
.B1(n_22),
.B2(n_84),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_153),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_182),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_181),
.A2(n_188),
.B1(n_159),
.B2(n_165),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_147),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_196),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_198),
.B1(n_200),
.B2(n_178),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_144),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_191),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_136),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_136),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_196),
.C(n_197),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_84),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_156),
.A2(n_167),
.B1(n_163),
.B2(n_160),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_169),
.A2(n_80),
.B1(n_22),
.B2(n_25),
.Y(n_200)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_172),
.C(n_175),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_203),
.C(n_206),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_166),
.C(n_171),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_204),
.A2(n_213),
.B1(n_216),
.B2(n_19),
.Y(n_226)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_171),
.C(n_174),
.Y(n_206)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_157),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_214),
.C(n_19),
.Y(n_230)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_184),
.B(n_193),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_212),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_155),
.B1(n_164),
.B2(n_158),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_162),
.C(n_176),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_177),
.Y(n_215)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_172),
.B1(n_179),
.B2(n_173),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_9),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_217),
.A2(n_218),
.B(n_14),
.Y(n_233)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_183),
.B(n_190),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_223),
.B1(n_232),
.B2(n_235),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_197),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_6),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_22),
.B1(n_16),
.B2(n_20),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_14),
.C(n_19),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_204),
.A2(n_22),
.B1(n_25),
.B2(n_14),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_231),
.B(n_7),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_202),
.A2(n_201),
.B(n_210),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_236),
.B(n_219),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_7),
.Y(n_235)
);

INVxp67_ASAP7_75t_SL g236 ( 
.A(n_208),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_219),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_239),
.B(n_241),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_2),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_221),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_242),
.A2(n_245),
.B(n_0),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_225),
.B(n_208),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_243),
.A2(n_248),
.B(n_249),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_19),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_247),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_19),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_14),
.C(n_1),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_14),
.C(n_1),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_2),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_232),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_251),
.B(n_259),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_244),
.A2(n_224),
.B1(n_225),
.B2(n_228),
.Y(n_254)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_248),
.A2(n_224),
.B1(n_228),
.B2(n_229),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_258),
.C(n_4),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_250),
.B(n_235),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_260),
.B(n_4),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_249),
.A2(n_223),
.B1(n_2),
.B2(n_3),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_6),
.B1(n_2),
.B2(n_3),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_261),
.B(n_5),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_4),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_3),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_263),
.A2(n_265),
.B(n_267),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_8),
.B(n_9),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_269),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_5),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_271),
.B(n_8),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_252),
.B(n_6),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_6),
.B(n_7),
.Y(n_271)
);

AO21x1_ASAP7_75t_L g275 ( 
.A1(n_272),
.A2(n_258),
.B(n_257),
.Y(n_275)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_275),
.Y(n_281)
);

OAI21x1_ASAP7_75t_L g276 ( 
.A1(n_270),
.A2(n_257),
.B(n_261),
.Y(n_276)
);

NAND4xp25_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_277),
.C(n_8),
.D(n_11),
.Y(n_280)
);

OAI21x1_ASAP7_75t_L g277 ( 
.A1(n_270),
.A2(n_7),
.B(n_8),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_278),
.B(n_279),
.Y(n_283)
);

OAI21x1_ASAP7_75t_SL g284 ( 
.A1(n_280),
.A2(n_11),
.B(n_12),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_11),
.C(n_12),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_274),
.C(n_12),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_285),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_286),
.B(n_281),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_283),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_282),
.Y(n_289)
);


endmodule