module fake_jpeg_3189_n_237 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_237);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_235;
wire n_103;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_50),
.Y(n_57)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_14),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

BUFx24_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_20),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_20),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_83),
.Y(n_87)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_81),
.Y(n_90)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_49),
.B1(n_48),
.B2(n_47),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_92),
.B(n_57),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_82),
.A2(n_55),
.B1(n_72),
.B2(n_53),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_79),
.B1(n_68),
.B2(n_58),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_56),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_66),
.C(n_75),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_72),
.B(n_71),
.C(n_64),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_99),
.B(n_79),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_65),
.B1(n_76),
.B2(n_53),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_85),
.B1(n_63),
.B2(n_55),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_101),
.B1(n_112),
.B2(n_67),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_85),
.B1(n_70),
.B2(n_65),
.Y(n_101)
);

NAND2x1_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_81),
.Y(n_102)
);

XNOR2x1_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_118),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_104),
.B(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_74),
.B1(n_77),
.B2(n_62),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_73),
.B1(n_62),
.B2(n_77),
.Y(n_121)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_111),
.B(n_0),
.Y(n_133)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_57),
.B(n_64),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_99),
.A2(n_76),
.B1(n_66),
.B2(n_70),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_54),
.Y(n_132)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_118),
.B(n_60),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_120),
.B(n_5),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_131),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_88),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_2),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_91),
.B1(n_88),
.B2(n_73),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_124),
.A2(n_127),
.B1(n_6),
.B2(n_7),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_75),
.B1(n_74),
.B2(n_93),
.Y(n_127)
);

OAI32xp33_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_58),
.A3(n_54),
.B1(n_68),
.B2(n_93),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_4),
.C(n_5),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_135),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_67),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_46),
.B1(n_45),
.B2(n_42),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_138),
.A2(n_40),
.B1(n_39),
.B2(n_38),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_1),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_31),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_124),
.A2(n_2),
.B(n_3),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_162),
.B(n_8),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_154),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_130),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_152),
.Y(n_170)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_126),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

OR2x2_ASAP7_75t_SL g153 ( 
.A(n_136),
.B(n_3),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_15),
.B(n_16),
.Y(n_182)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_37),
.B1(n_36),
.B2(n_32),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_160),
.B1(n_121),
.B2(n_127),
.Y(n_168)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_161),
.Y(n_171)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_140),
.A2(n_6),
.B(n_7),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_164),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_8),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_136),
.C(n_137),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_176),
.C(n_183),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_168),
.A2(n_178),
.B1(n_181),
.B2(n_150),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_175),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_146),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_149),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_119),
.C(n_125),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_158),
.A2(n_125),
.B(n_10),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_180),
.C(n_182),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_160),
.B(n_154),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_156),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_26),
.C(n_25),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_15),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_145),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_200),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_145),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_187),
.B(n_190),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_150),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_191),
.B(n_192),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_177),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_195),
.B1(n_182),
.B2(n_165),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_180),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_21),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_197),
.C(n_172),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_166),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_179),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_165),
.Y(n_211)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_22),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_171),
.B(n_184),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_184),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_202),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_205),
.Y(n_213)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_185),
.C(n_183),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_23),
.Y(n_218)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_211),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_212),
.A2(n_188),
.B1(n_190),
.B2(n_22),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_214),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_202),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_217),
.B(n_221),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_206),
.Y(n_222)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_224),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_208),
.B(n_203),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_206),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_226),
.B(n_213),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_227),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_223),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_229),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_231),
.A2(n_216),
.B1(n_220),
.B2(n_228),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_219),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_225),
.C(n_226),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_234),
.A2(n_218),
.B(n_204),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_235),
.B(n_210),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_23),
.Y(n_237)
);


endmodule