module fake_aes_6531_n_688 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_688);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_688;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_462;
wire n_232;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_195;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g73 ( .A(n_17), .Y(n_73) );
CKINVDCx5p33_ASAP7_75t_R g74 ( .A(n_40), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_70), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_3), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_48), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_16), .Y(n_78) );
HB1xp67_ASAP7_75t_L g79 ( .A(n_66), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_71), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_32), .Y(n_81) );
INVxp33_ASAP7_75t_SL g82 ( .A(n_27), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_5), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_17), .Y(n_84) );
INVxp67_ASAP7_75t_L g85 ( .A(n_37), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_35), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_38), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_28), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_33), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_21), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_1), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_16), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_24), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_67), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_30), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_53), .Y(n_96) );
INVxp33_ASAP7_75t_L g97 ( .A(n_60), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_36), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_55), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_21), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_57), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_7), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_47), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_6), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_34), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_52), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_7), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_26), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_50), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_29), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_0), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_3), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_2), .Y(n_114) );
CKINVDCx14_ASAP7_75t_R g115 ( .A(n_14), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_69), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_43), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_19), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_45), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_2), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_39), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_77), .Y(n_122) );
NOR3xp33_ASAP7_75t_L g123 ( .A(n_111), .B(n_1), .C(n_4), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g124 ( .A(n_97), .B(n_4), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_77), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_115), .Y(n_126) );
CKINVDCx11_ASAP7_75t_R g127 ( .A(n_94), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_80), .Y(n_128) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_80), .A2(n_5), .B(n_6), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_81), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_98), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_98), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_87), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_76), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_79), .B(n_8), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_76), .B(n_8), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_87), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_88), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_88), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_74), .Y(n_143) );
XOR2xp5_ASAP7_75t_L g144 ( .A(n_73), .B(n_9), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_89), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_92), .B(n_9), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_89), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_78), .B(n_10), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_92), .B(n_10), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_93), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_93), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_95), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_78), .B(n_11), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_95), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_85), .B(n_11), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_116), .Y(n_156) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_83), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_116), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_117), .Y(n_159) );
OAI21x1_ASAP7_75t_L g160 ( .A1(n_117), .A2(n_42), .B(n_68), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_119), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_119), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_75), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_96), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_99), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_83), .B(n_12), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_165), .B(n_122), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_134), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_143), .B(n_82), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_143), .B(n_121), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_134), .Y(n_171) );
AND2x6_ASAP7_75t_L g172 ( .A(n_146), .B(n_103), .Y(n_172) );
INVx5_ASAP7_75t_L g173 ( .A(n_151), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
NAND2x1p5_ASAP7_75t_L g175 ( .A(n_129), .B(n_105), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_146), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_146), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_122), .B(n_125), .Y(n_179) );
INVx1_ASAP7_75t_SL g180 ( .A(n_126), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_134), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_149), .Y(n_182) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_144), .Y(n_183) );
BUFx8_ASAP7_75t_SL g184 ( .A(n_126), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_149), .B(n_120), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_149), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_149), .B(n_120), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_151), .Y(n_188) );
NAND2x1p5_ASAP7_75t_L g189 ( .A(n_129), .B(n_108), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_149), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_165), .B(n_106), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_137), .A2(n_90), .B1(n_114), .B2(n_91), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_151), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_137), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_163), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_125), .B(n_109), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_151), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_127), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_128), .B(n_74), .Y(n_199) );
INVx4_ASAP7_75t_L g200 ( .A(n_130), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_128), .B(n_106), .Y(n_201) );
OAI22xp5_ASAP7_75t_SL g202 ( .A1(n_144), .A2(n_118), .B1(n_100), .B2(n_84), .Y(n_202) );
AND2x6_ASAP7_75t_L g203 ( .A(n_139), .B(n_110), .Y(n_203) );
INVx2_ASAP7_75t_SL g204 ( .A(n_157), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_151), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_151), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_134), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_127), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_134), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_134), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_151), .Y(n_211) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_160), .A2(n_114), .B(n_90), .Y(n_212) );
BUFx3_ASAP7_75t_L g213 ( .A(n_163), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_131), .B(n_101), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_134), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_151), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_154), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_131), .B(n_101), .Y(n_218) );
INVx4_ASAP7_75t_L g219 ( .A(n_130), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_134), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_157), .B(n_139), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_154), .Y(n_222) );
OR2x2_ASAP7_75t_L g223 ( .A(n_138), .B(n_91), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_154), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_132), .B(n_113), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_132), .B(n_107), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_154), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_138), .A2(n_84), .B1(n_104), .B2(n_102), .Y(n_228) );
OR2x2_ASAP7_75t_L g229 ( .A(n_136), .B(n_150), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_154), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_154), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_154), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_154), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_158), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_229), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_200), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_194), .B(n_139), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_194), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_229), .Y(n_239) );
BUFx3_ASAP7_75t_L g240 ( .A(n_172), .Y(n_240) );
BUFx12f_ASAP7_75t_L g241 ( .A(n_198), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_221), .A2(n_147), .B(n_141), .C(n_140), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_174), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_174), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_204), .B(n_152), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_204), .B(n_166), .Y(n_246) );
OR2x6_ASAP7_75t_L g247 ( .A(n_202), .B(n_166), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_221), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_185), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_199), .B(n_152), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_201), .B(n_136), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_179), .A2(n_150), .B(n_140), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_185), .B(n_187), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_174), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_223), .B(n_155), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_185), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_185), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_178), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_218), .B(n_162), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_200), .Y(n_260) );
AND3x1_ASAP7_75t_SL g261 ( .A(n_202), .B(n_144), .C(n_112), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_200), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_187), .B(n_166), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_187), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_200), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_219), .Y(n_266) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_178), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_223), .B(n_155), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_203), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_214), .B(n_162), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_219), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_182), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_172), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_178), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_219), .Y(n_275) );
INVx1_ASAP7_75t_SL g276 ( .A(n_180), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_191), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_187), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_182), .B(n_123), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_219), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_170), .B(n_153), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_182), .B(n_123), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_167), .B(n_142), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_175), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_182), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_175), .Y(n_286) );
AOI22x1_ASAP7_75t_L g287 ( .A1(n_175), .A2(n_164), .B1(n_147), .B2(n_141), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_172), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_169), .B(n_148), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_186), .B(n_145), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_186), .B(n_148), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_203), .A2(n_124), .B1(n_153), .B2(n_130), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_203), .B(n_145), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_L g294 ( .A1(n_176), .A2(n_141), .B(n_147), .C(n_133), .Y(n_294) );
OR2x6_ASAP7_75t_L g295 ( .A(n_192), .B(n_124), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_186), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_186), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_172), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_172), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_203), .B(n_145), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_189), .B(n_145), .Y(n_301) );
NOR2xp67_ASAP7_75t_L g302 ( .A(n_208), .B(n_130), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_183), .B(n_142), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_203), .B(n_160), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_176), .Y(n_305) );
OR2x6_ASAP7_75t_L g306 ( .A(n_176), .B(n_160), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_243), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_253), .Y(n_308) );
INVx3_ASAP7_75t_L g309 ( .A(n_243), .Y(n_309) );
BUFx12f_ASAP7_75t_L g310 ( .A(n_241), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_243), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_236), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_236), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_305), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_260), .Y(n_315) );
INVx4_ASAP7_75t_L g316 ( .A(n_253), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_243), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_260), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_262), .Y(n_319) );
AOI21xp33_ASAP7_75t_L g320 ( .A1(n_238), .A2(n_228), .B(n_190), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_240), .Y(n_321) );
A2O1A1Ixp33_ASAP7_75t_L g322 ( .A1(n_281), .A2(n_190), .B(n_177), .C(n_196), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_240), .Y(n_323) );
NOR2xp67_ASAP7_75t_L g324 ( .A(n_272), .B(n_177), .Y(n_324) );
CKINVDCx6p67_ASAP7_75t_R g325 ( .A(n_241), .Y(n_325) );
INVx5_ASAP7_75t_L g326 ( .A(n_244), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_262), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_263), .B(n_203), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_301), .A2(n_177), .B(n_190), .Y(n_329) );
AOI222xp33_ASAP7_75t_L g330 ( .A1(n_248), .A2(n_208), .B1(n_225), .B2(n_226), .C1(n_203), .C2(n_172), .Y(n_330) );
AND2x6_ASAP7_75t_L g331 ( .A(n_273), .B(n_172), .Y(n_331) );
INVx8_ASAP7_75t_L g332 ( .A(n_253), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_273), .Y(n_333) );
INVx2_ASAP7_75t_SL g334 ( .A(n_238), .Y(n_334) );
AOI22xp33_ASAP7_75t_SL g335 ( .A1(n_247), .A2(n_189), .B1(n_129), .B2(n_130), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_265), .Y(n_336) );
INVx4_ASAP7_75t_L g337 ( .A(n_288), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_263), .B(n_135), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_301), .A2(n_212), .B(n_189), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_279), .B(n_164), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_290), .A2(n_212), .B(n_188), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_265), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_288), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_244), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_266), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_266), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_271), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_276), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_244), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_303), .Y(n_350) );
CKINVDCx6p67_ASAP7_75t_R g351 ( .A(n_247), .Y(n_351) );
NOR2xp67_ASAP7_75t_L g352 ( .A(n_272), .B(n_296), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_271), .Y(n_353) );
INVx3_ASAP7_75t_L g354 ( .A(n_244), .Y(n_354) );
CKINVDCx11_ASAP7_75t_R g355 ( .A(n_247), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_290), .A2(n_212), .B(n_188), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_275), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_298), .Y(n_358) );
CKINVDCx11_ASAP7_75t_R g359 ( .A(n_295), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_248), .B(n_184), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_277), .B(n_135), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_298), .Y(n_362) );
OR2x6_ASAP7_75t_L g363 ( .A(n_299), .B(n_129), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_359), .A2(n_282), .B1(n_279), .B2(n_295), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_350), .A2(n_268), .B1(n_255), .B2(n_289), .C(n_281), .Y(n_365) );
NOR2xp67_ASAP7_75t_L g366 ( .A(n_334), .B(n_304), .Y(n_366) );
AOI21xp33_ASAP7_75t_L g367 ( .A1(n_330), .A2(n_335), .B(n_304), .Y(n_367) );
CKINVDCx14_ASAP7_75t_R g368 ( .A(n_325), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_340), .B(n_263), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_308), .A2(n_282), .B1(n_279), .B2(n_295), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_322), .A2(n_242), .B1(n_239), .B2(n_235), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_308), .A2(n_282), .B1(n_246), .B2(n_237), .Y(n_372) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_321), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_355), .A2(n_237), .B1(n_246), .B2(n_255), .Y(n_374) );
BUFx3_ASAP7_75t_L g375 ( .A(n_332), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_312), .Y(n_376) );
O2A1O1Ixp5_ASAP7_75t_SL g377 ( .A1(n_307), .A2(n_135), .B(n_156), .C(n_142), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_332), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_340), .A2(n_242), .B1(n_304), .B2(n_294), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_340), .A2(n_294), .B1(n_306), .B2(n_268), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_316), .B(n_299), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_351), .A2(n_246), .B1(n_237), .B2(n_269), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_351), .A2(n_340), .B1(n_316), .B2(n_332), .Y(n_383) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_321), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_314), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_316), .A2(n_278), .B1(n_256), .B2(n_257), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_314), .B(n_291), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_312), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g389 ( .A1(n_338), .A2(n_270), .B1(n_245), .B2(n_250), .C(n_259), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_315), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_361), .B(n_291), .Y(n_391) );
OAI221xp5_ASAP7_75t_L g392 ( .A1(n_348), .A2(n_302), .B1(n_292), .B2(n_251), .C(n_249), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_332), .Y(n_393) );
INVx1_ASAP7_75t_SL g394 ( .A(n_332), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_315), .B(n_318), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_313), .Y(n_396) );
AOI211xp5_ASAP7_75t_L g397 ( .A1(n_360), .A2(n_261), .B(n_300), .C(n_293), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g398 ( .A1(n_325), .A2(n_264), .B1(n_283), .B2(n_306), .Y(n_398) );
OAI221xp5_ASAP7_75t_L g399 ( .A1(n_365), .A2(n_328), .B1(n_320), .B2(n_334), .C(n_324), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_395), .B(n_318), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_376), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_389), .A2(n_363), .B1(n_352), .B2(n_310), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_371), .A2(n_252), .B1(n_142), .B2(n_135), .C(n_156), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_364), .A2(n_363), .B1(n_352), .B2(n_310), .Y(n_404) );
OAI22xp33_ASAP7_75t_L g405 ( .A1(n_391), .A2(n_363), .B1(n_306), .B2(n_342), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_380), .A2(n_339), .B(n_341), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_398), .A2(n_306), .B1(n_147), .B2(n_141), .Y(n_407) );
BUFx12f_ASAP7_75t_L g408 ( .A(n_368), .Y(n_408) );
BUFx12f_ASAP7_75t_L g409 ( .A(n_378), .Y(n_409) );
OAI21x1_ASAP7_75t_L g410 ( .A1(n_377), .A2(n_356), .B(n_287), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_375), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_367), .A2(n_254), .B1(n_258), .B2(n_267), .Y(n_412) );
OAI21xp33_ASAP7_75t_L g413 ( .A1(n_391), .A2(n_164), .B(n_329), .Y(n_413) );
AO21x2_ASAP7_75t_L g414 ( .A1(n_380), .A2(n_164), .B(n_133), .Y(n_414) );
AOI222xp33_ASAP7_75t_L g415 ( .A1(n_374), .A2(n_370), .B1(n_371), .B2(n_372), .C1(n_369), .C2(n_385), .Y(n_415) );
INVx8_ASAP7_75t_L g416 ( .A(n_381), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_390), .A2(n_156), .B1(n_135), .B2(n_326), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_395), .B(n_336), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_397), .A2(n_156), .B1(n_297), .B2(n_285), .C(n_342), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_390), .A2(n_326), .B1(n_286), .B2(n_284), .Y(n_420) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_387), .A2(n_336), .B1(n_357), .B2(n_326), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_385), .B(n_357), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_369), .A2(n_267), .B1(n_254), .B2(n_258), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_397), .A2(n_133), .B1(n_163), .B2(n_161), .C(n_159), .Y(n_424) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_382), .A2(n_272), .B1(n_296), .B2(n_133), .C(n_254), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_408), .Y(n_426) );
OAI22xp33_ASAP7_75t_L g427 ( .A1(n_411), .A2(n_375), .B1(n_394), .B2(n_393), .Y(n_427) );
OAI211xp5_ASAP7_75t_L g428 ( .A1(n_415), .A2(n_383), .B(n_386), .C(n_392), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_407), .A2(n_366), .B1(n_387), .B2(n_379), .Y(n_429) );
OR2x6_ASAP7_75t_L g430 ( .A(n_407), .B(n_366), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_402), .A2(n_379), .B1(n_376), .B2(n_388), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_415), .A2(n_375), .B1(n_381), .B2(n_396), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_400), .B(n_388), .Y(n_433) );
OAI21x1_ASAP7_75t_L g434 ( .A1(n_406), .A2(n_377), .B(n_396), .Y(n_434) );
AOI222xp33_ASAP7_75t_L g435 ( .A1(n_408), .A2(n_161), .B1(n_159), .B2(n_158), .C1(n_163), .C2(n_381), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_401), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_400), .B(n_373), .Y(n_437) );
INVx1_ASAP7_75t_SL g438 ( .A(n_409), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_418), .B(n_129), .Y(n_439) );
INVx2_ASAP7_75t_SL g440 ( .A(n_409), .Y(n_440) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_404), .A2(n_163), .B1(n_159), .B2(n_161), .C(n_158), .Y(n_441) );
INVxp67_ASAP7_75t_L g442 ( .A(n_418), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_422), .B(n_381), .Y(n_443) );
OAI21xp5_ASAP7_75t_L g444 ( .A1(n_399), .A2(n_419), .B(n_424), .Y(n_444) );
OA21x2_ASAP7_75t_L g445 ( .A1(n_410), .A2(n_209), .B(n_171), .Y(n_445) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_410), .A2(n_209), .B(n_171), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_414), .A2(n_274), .B1(n_267), .B2(n_258), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_405), .A2(n_284), .B1(n_286), .B2(n_326), .Y(n_448) );
INVx5_ASAP7_75t_L g449 ( .A(n_416), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_422), .B(n_373), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_401), .B(n_313), .Y(n_451) );
INVxp67_ASAP7_75t_L g452 ( .A(n_411), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_414), .A2(n_274), .B1(n_344), .B2(n_349), .Y(n_453) );
AOI22xp33_ASAP7_75t_SL g454 ( .A1(n_416), .A2(n_331), .B1(n_384), .B2(n_373), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_417), .A2(n_326), .B1(n_344), .B2(n_349), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_414), .A2(n_274), .B1(n_331), .B2(n_307), .Y(n_456) );
NOR2xp67_ASAP7_75t_L g457 ( .A(n_420), .B(n_417), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_420), .Y(n_458) );
OAI221xp5_ASAP7_75t_SL g459 ( .A1(n_412), .A2(n_319), .B1(n_327), .B2(n_353), .C(n_347), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_432), .A2(n_416), .B1(n_425), .B2(n_413), .Y(n_460) );
OAI22xp5_ASAP7_75t_SL g461 ( .A1(n_426), .A2(n_416), .B1(n_423), .B2(n_326), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_436), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_442), .B(n_416), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_436), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_458), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_433), .B(n_421), .Y(n_466) );
OAI221xp5_ASAP7_75t_L g467 ( .A1(n_428), .A2(n_413), .B1(n_403), .B2(n_158), .C(n_159), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_458), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_445), .Y(n_469) );
AO31x2_ASAP7_75t_L g470 ( .A1(n_431), .A2(n_319), .A3(n_353), .B(n_347), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_457), .A2(n_430), .B1(n_429), .B2(n_444), .Y(n_471) );
BUFx3_ASAP7_75t_L g472 ( .A(n_449), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_433), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_450), .B(n_158), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_437), .B(n_373), .Y(n_475) );
OAI31xp33_ASAP7_75t_L g476 ( .A1(n_427), .A2(n_307), .A3(n_354), .B(n_309), .Y(n_476) );
BUFx2_ASAP7_75t_L g477 ( .A(n_450), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_457), .A2(n_158), .B1(n_159), .B2(n_161), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_450), .B(n_158), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_445), .Y(n_480) );
OAI22xp5_ASAP7_75t_SL g481 ( .A1(n_438), .A2(n_337), .B1(n_384), .B2(n_373), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_449), .A2(n_430), .B1(n_454), .B2(n_459), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_443), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_437), .B(n_159), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_430), .Y(n_485) );
OR2x2_ASAP7_75t_SL g486 ( .A(n_449), .B(n_373), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_451), .B(n_161), .Y(n_487) );
AOI21x1_ASAP7_75t_L g488 ( .A1(n_446), .A2(n_220), .B(n_181), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_449), .A2(n_384), .B1(n_311), .B2(n_317), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_451), .Y(n_490) );
OAI31xp33_ASAP7_75t_L g491 ( .A1(n_441), .A2(n_317), .A3(n_296), .B(n_345), .Y(n_491) );
OAI33xp33_ASAP7_75t_L g492 ( .A1(n_452), .A2(n_12), .A3(n_13), .B1(n_14), .B2(n_15), .B3(n_18), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_439), .B(n_161), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_449), .A2(n_317), .B(n_327), .C(n_346), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_430), .B(n_384), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_439), .B(n_161), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_434), .B(n_163), .Y(n_497) );
OAI221xp5_ASAP7_75t_SL g498 ( .A1(n_435), .A2(n_345), .B1(n_346), .B2(n_18), .C(n_19), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_440), .B(n_163), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_440), .B(n_13), .Y(n_500) );
AND2x2_ASAP7_75t_SL g501 ( .A(n_456), .B(n_384), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_448), .A2(n_384), .B1(n_337), .B2(n_274), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g503 ( .A1(n_455), .A2(n_331), .B1(n_337), .B2(n_343), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_453), .B(n_15), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_447), .B(n_20), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_434), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_445), .B(n_20), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_445), .B(n_22), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_473), .B(n_22), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_473), .B(n_23), .Y(n_510) );
OAI321xp33_ASAP7_75t_L g511 ( .A1(n_498), .A2(n_482), .A3(n_485), .B1(n_461), .B2(n_500), .C(n_504), .Y(n_511) );
OAI332xp33_ASAP7_75t_L g512 ( .A1(n_500), .A2(n_23), .A3(n_220), .B1(n_215), .B2(n_197), .B3(n_206), .C1(n_205), .C2(n_211), .Y(n_512) );
INVxp67_ASAP7_75t_L g513 ( .A(n_507), .Y(n_513) );
INVx3_ASAP7_75t_SL g514 ( .A(n_486), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_464), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_464), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_483), .B(n_446), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_490), .B(n_215), .Y(n_518) );
NOR3xp33_ASAP7_75t_L g519 ( .A(n_492), .B(n_193), .C(n_197), .Y(n_519) );
NAND3xp33_ASAP7_75t_L g520 ( .A(n_499), .B(n_168), .C(n_207), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_490), .B(n_25), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_462), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_477), .B(n_31), .Y(n_523) );
NAND4xp25_ASAP7_75t_L g524 ( .A(n_460), .B(n_205), .C(n_193), .D(n_206), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_474), .B(n_41), .Y(n_525) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_472), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_465), .B(n_210), .Y(n_527) );
NOR3xp33_ASAP7_75t_L g528 ( .A(n_467), .B(n_211), .C(n_216), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_469), .Y(n_529) );
OAI211xp5_ASAP7_75t_SL g530 ( .A1(n_499), .A2(n_227), .B(n_231), .C(n_222), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_469), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_465), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_481), .A2(n_362), .B(n_358), .Y(n_533) );
BUFx3_ASAP7_75t_L g534 ( .A(n_486), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_468), .Y(n_535) );
AOI221xp5_ASAP7_75t_L g536 ( .A1(n_468), .A2(n_222), .B1(n_216), .B2(n_227), .C(n_231), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_466), .B(n_44), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_506), .B(n_207), .C(n_210), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_479), .B(n_207), .Y(n_539) );
NOR3xp33_ASAP7_75t_L g540 ( .A(n_505), .B(n_224), .C(n_233), .Y(n_540) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_472), .B(n_362), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_479), .B(n_46), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_484), .B(n_207), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_507), .Y(n_544) );
OAI22xp5_ASAP7_75t_SL g545 ( .A1(n_485), .A2(n_362), .B1(n_358), .B2(n_343), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_463), .B(n_49), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_508), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_484), .B(n_51), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_493), .B(n_210), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_504), .B(n_54), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_508), .B(n_56), .Y(n_551) );
OAI21xp5_ASAP7_75t_L g552 ( .A1(n_478), .A2(n_331), .B(n_233), .Y(n_552) );
NAND3xp33_ASAP7_75t_SL g553 ( .A(n_476), .B(n_58), .C(n_59), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_466), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_496), .B(n_61), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_493), .Y(n_556) );
INVxp67_ASAP7_75t_L g557 ( .A(n_497), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_487), .B(n_168), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_487), .B(n_168), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_475), .B(n_62), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_475), .B(n_207), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_497), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_554), .B(n_506), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_544), .B(n_470), .Y(n_564) );
INVx6_ASAP7_75t_L g565 ( .A(n_526), .Y(n_565) );
OAI21xp33_ASAP7_75t_L g566 ( .A1(n_534), .A2(n_501), .B(n_495), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_547), .B(n_470), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_515), .B(n_470), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_516), .B(n_470), .Y(n_569) );
INVxp67_ASAP7_75t_SL g570 ( .A(n_557), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_532), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_535), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_522), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_513), .B(n_470), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_513), .B(n_495), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_514), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_534), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_550), .A2(n_501), .B1(n_503), .B2(n_502), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_557), .B(n_480), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_510), .B(n_480), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_556), .B(n_562), .Y(n_581) );
NAND2x1_ASAP7_75t_L g582 ( .A(n_511), .B(n_541), .Y(n_582) );
AND2x4_ASAP7_75t_L g583 ( .A(n_529), .B(n_488), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_512), .B(n_489), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_529), .B(n_488), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_509), .B(n_491), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_531), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_517), .B(n_494), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_537), .B(n_210), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_551), .B(n_168), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_523), .B(n_63), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_527), .B(n_168), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_550), .A2(n_331), .B1(n_210), .B2(n_343), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_539), .B(n_64), .Y(n_594) );
NAND4xp25_ASAP7_75t_L g595 ( .A(n_546), .B(n_224), .C(n_195), .D(n_213), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_538), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_518), .Y(n_597) );
NAND2xp33_ASAP7_75t_L g598 ( .A(n_521), .B(n_331), .Y(n_598) );
NOR3xp33_ASAP7_75t_L g599 ( .A(n_553), .B(n_234), .C(n_217), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_543), .B(n_65), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_546), .A2(n_362), .B1(n_358), .B2(n_321), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_561), .B(n_72), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_525), .B(n_230), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_542), .B(n_230), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_548), .B(n_230), .Y(n_605) );
OR2x6_ASAP7_75t_L g606 ( .A(n_545), .B(n_362), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_520), .Y(n_607) );
CKINVDCx16_ASAP7_75t_R g608 ( .A(n_553), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_558), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_570), .B(n_519), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_571), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_584), .A2(n_540), .B1(n_524), .B2(n_528), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_572), .Y(n_613) );
XOR2x2_ASAP7_75t_L g614 ( .A(n_576), .B(n_560), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_573), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_597), .B(n_540), .Y(n_616) );
INVxp67_ASAP7_75t_SL g617 ( .A(n_596), .Y(n_617) );
AOI211xp5_ASAP7_75t_SL g618 ( .A1(n_598), .A2(n_560), .B(n_533), .C(n_530), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_574), .B(n_559), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_608), .B(n_555), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_581), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_563), .Y(n_622) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_582), .A2(n_552), .B1(n_530), .B2(n_549), .C(n_536), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_565), .B(n_232), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_574), .B(n_230), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_577), .B(n_232), .Y(n_626) );
INVxp33_ASAP7_75t_L g627 ( .A(n_596), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_578), .A2(n_358), .B1(n_343), .B2(n_333), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_609), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_584), .A2(n_232), .B1(n_343), .B2(n_333), .Y(n_630) );
INVx3_ASAP7_75t_SL g631 ( .A(n_591), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_577), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_579), .Y(n_633) );
INVx2_ASAP7_75t_SL g634 ( .A(n_587), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_575), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_580), .B(n_232), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_564), .B(n_195), .Y(n_637) );
INVx1_ASAP7_75t_SL g638 ( .A(n_590), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_585), .Y(n_639) );
INVx2_ASAP7_75t_SL g640 ( .A(n_591), .Y(n_640) );
OAI22xp5_ASAP7_75t_SL g641 ( .A1(n_606), .A2(n_333), .B1(n_323), .B2(n_321), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_585), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g643 ( .A(n_599), .B(n_173), .C(n_333), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_567), .B(n_173), .Y(n_644) );
NOR3xp33_ASAP7_75t_L g645 ( .A(n_607), .B(n_217), .C(n_234), .Y(n_645) );
AOI211x1_ASAP7_75t_L g646 ( .A1(n_566), .A2(n_173), .B(n_213), .C(n_333), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_598), .A2(n_321), .B(n_323), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_568), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_569), .Y(n_649) );
AOI221xp5_ASAP7_75t_SL g650 ( .A1(n_586), .A2(n_323), .B1(n_217), .B2(n_234), .C(n_275), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_588), .Y(n_651) );
INVxp67_ASAP7_75t_L g652 ( .A(n_595), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_583), .B(n_280), .Y(n_653) );
XOR2x2_ASAP7_75t_L g654 ( .A(n_593), .B(n_601), .Y(n_654) );
O2A1O1Ixp33_ASAP7_75t_L g655 ( .A1(n_589), .A2(n_605), .B(n_604), .C(n_603), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_602), .Y(n_656) );
INVxp67_ASAP7_75t_SL g657 ( .A(n_583), .Y(n_657) );
AOI21xp33_ASAP7_75t_SL g658 ( .A1(n_606), .A2(n_594), .B(n_600), .Y(n_658) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_592), .B(n_471), .C(n_584), .D(n_360), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_629), .Y(n_660) );
AOI221xp5_ASAP7_75t_L g661 ( .A1(n_651), .A2(n_627), .B1(n_617), .B2(n_621), .C(n_659), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_622), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_627), .A2(n_635), .B1(n_649), .B2(n_648), .C(n_611), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_631), .A2(n_620), .B1(n_633), .B2(n_656), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_634), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_613), .A2(n_610), .B1(n_632), .B2(n_615), .C(n_612), .Y(n_666) );
OAI21xp5_ASAP7_75t_SL g667 ( .A1(n_618), .A2(n_658), .B(n_612), .Y(n_667) );
OAI321xp33_ASAP7_75t_L g668 ( .A1(n_628), .A2(n_640), .A3(n_652), .B1(n_623), .B2(n_616), .C(n_657), .Y(n_668) );
AOI321xp33_ASAP7_75t_L g669 ( .A1(n_655), .A2(n_619), .A3(n_625), .B1(n_642), .B2(n_639), .C(n_624), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_650), .B(n_645), .C(n_624), .Y(n_670) );
NAND2xp33_ASAP7_75t_SL g671 ( .A(n_614), .B(n_634), .Y(n_671) );
OAI211xp5_ASAP7_75t_L g672 ( .A1(n_667), .A2(n_646), .B(n_625), .C(n_643), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_671), .A2(n_654), .B1(n_638), .B2(n_644), .C(n_626), .Y(n_673) );
NOR3xp33_ASAP7_75t_L g674 ( .A(n_668), .B(n_626), .C(n_636), .Y(n_674) );
AOI211xp5_ASAP7_75t_SL g675 ( .A1(n_664), .A2(n_641), .B(n_637), .C(n_630), .Y(n_675) );
NAND2x1p5_ASAP7_75t_L g676 ( .A(n_662), .B(n_647), .Y(n_676) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_665), .Y(n_677) );
OAI222xp33_ASAP7_75t_L g678 ( .A1(n_673), .A2(n_665), .B1(n_669), .B2(n_660), .C1(n_661), .C2(n_666), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_677), .Y(n_679) );
NAND5xp2_ASAP7_75t_L g680 ( .A(n_675), .B(n_663), .C(n_670), .D(n_653), .E(n_592), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_676), .Y(n_681) );
NOR3xp33_ASAP7_75t_L g682 ( .A(n_678), .B(n_672), .C(n_674), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_679), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_682), .B(n_681), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_684), .Y(n_685) );
AND2x4_ASAP7_75t_L g686 ( .A(n_685), .B(n_683), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_686), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_687), .B(n_680), .Y(n_688) );
endmodule