module fake_aes_9835_n_33 (n_1, n_2, n_4, n_3, n_5, n_0, n_33);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_6;
wire n_7;
wire n_29;
INVx1_ASAP7_75t_L g6 ( .A(n_2), .Y(n_6) );
BUFx2_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_3), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_1), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_4), .Y(n_10) );
NAND2xp5_ASAP7_75t_SL g11 ( .A(n_7), .B(n_0), .Y(n_11) );
AOI21xp5_ASAP7_75t_L g12 ( .A1(n_6), .A2(n_0), .B(n_1), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_7), .B(n_0), .Y(n_13) );
OAI21x1_ASAP7_75t_L g14 ( .A1(n_6), .A2(n_1), .B(n_2), .Y(n_14) );
O2A1O1Ixp5_ASAP7_75t_L g15 ( .A1(n_10), .A2(n_2), .B(n_3), .C(n_4), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_13), .B(n_7), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
BUFx3_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_19), .B(n_9), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_17), .Y(n_22) );
AOI22xp33_ASAP7_75t_SL g23 ( .A1(n_20), .A2(n_19), .B1(n_16), .B2(n_8), .Y(n_23) );
OAI22xp33_ASAP7_75t_SL g24 ( .A1(n_21), .A2(n_19), .B1(n_8), .B2(n_9), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_20), .B(n_16), .Y(n_25) );
AOI22xp5_ASAP7_75t_L g26 ( .A1(n_23), .A2(n_16), .B1(n_21), .B2(n_11), .Y(n_26) );
AOI221xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_15), .B1(n_12), .B2(n_18), .C(n_17), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_18), .Y(n_28) );
CKINVDCx5p33_ASAP7_75t_R g29 ( .A(n_26), .Y(n_29) );
AOI32xp33_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_17), .A3(n_24), .B1(n_3), .B2(n_4), .Y(n_30) );
OAI22xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_27), .B1(n_22), .B2(n_5), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
AOI22xp5_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_22), .B1(n_30), .B2(n_31), .Y(n_33) );
endmodule