module fake_aes_5296_n_490 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_490);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_490;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g74 ( .A(n_46), .Y(n_74) );
INVxp67_ASAP7_75t_SL g75 ( .A(n_45), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_56), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_6), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_25), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_8), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_53), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_72), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_63), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_1), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_57), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_16), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_31), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_9), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_52), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_64), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_26), .Y(n_90) );
HB1xp67_ASAP7_75t_L g91 ( .A(n_44), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_17), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_42), .Y(n_93) );
INVxp33_ASAP7_75t_SL g94 ( .A(n_48), .Y(n_94) );
CKINVDCx14_ASAP7_75t_R g95 ( .A(n_21), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_10), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_15), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_49), .Y(n_98) );
BUFx3_ASAP7_75t_L g99 ( .A(n_73), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_0), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_20), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_22), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_39), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_38), .Y(n_104) );
CKINVDCx14_ASAP7_75t_R g105 ( .A(n_37), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_19), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_8), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_99), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_74), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_74), .Y(n_110) );
AND2x4_ASAP7_75t_L g111 ( .A(n_83), .B(n_0), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_91), .B(n_1), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_76), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_76), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_95), .B(n_2), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_78), .Y(n_116) );
AND2x6_ASAP7_75t_L g117 ( .A(n_99), .B(n_33), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_77), .B(n_2), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_78), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_80), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_80), .Y(n_121) );
INVx4_ASAP7_75t_L g122 ( .A(n_82), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_81), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_81), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_77), .B(n_3), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_84), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_88), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_88), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_90), .Y(n_130) );
BUFx3_ASAP7_75t_L g131 ( .A(n_117), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_111), .B(n_83), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_122), .B(n_89), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_108), .Y(n_134) );
BUFx3_ASAP7_75t_L g135 ( .A(n_117), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_111), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_122), .B(n_93), .Y(n_137) );
INVxp67_ASAP7_75t_L g138 ( .A(n_115), .Y(n_138) );
AO22x2_ASAP7_75t_L g139 ( .A1(n_111), .A2(n_98), .B1(n_90), .B2(n_101), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_114), .B(n_98), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_122), .B(n_101), .Y(n_141) );
INVx2_ASAP7_75t_SL g142 ( .A(n_114), .Y(n_142) );
INVx1_ASAP7_75t_SL g143 ( .A(n_115), .Y(n_143) );
OR2x2_ASAP7_75t_L g144 ( .A(n_112), .B(n_107), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_108), .Y(n_145) );
INVx4_ASAP7_75t_L g146 ( .A(n_117), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_114), .B(n_104), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_115), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_108), .Y(n_149) );
INVx1_ASAP7_75t_SL g150 ( .A(n_112), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_117), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_128), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_108), .Y(n_153) );
AND2x6_ASAP7_75t_L g154 ( .A(n_111), .B(n_103), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_111), .B(n_92), .Y(n_155) );
BUFx4f_ASAP7_75t_L g156 ( .A(n_154), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_150), .B(n_122), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_132), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_150), .B(n_118), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_132), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_132), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_144), .B(n_122), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_132), .Y(n_163) );
OR2x6_ASAP7_75t_L g164 ( .A(n_139), .B(n_118), .Y(n_164) );
NAND2xp33_ASAP7_75t_L g165 ( .A(n_154), .B(n_117), .Y(n_165) );
INVx2_ASAP7_75t_SL g166 ( .A(n_139), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_132), .Y(n_167) );
OAI221xp5_ASAP7_75t_L g168 ( .A1(n_138), .A2(n_125), .B1(n_109), .B2(n_110), .C(n_116), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_136), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_139), .A2(n_119), .B1(n_110), .B2(n_116), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_136), .Y(n_171) );
INVx2_ASAP7_75t_SL g172 ( .A(n_139), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_144), .B(n_109), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_144), .B(n_121), .Y(n_174) );
BUFx2_ASAP7_75t_L g175 ( .A(n_139), .Y(n_175) );
INVx8_ASAP7_75t_L g176 ( .A(n_154), .Y(n_176) );
INVxp67_ASAP7_75t_L g177 ( .A(n_143), .Y(n_177) );
INVx2_ASAP7_75t_SL g178 ( .A(n_139), .Y(n_178) );
INVx1_ASAP7_75t_SL g179 ( .A(n_148), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_138), .A2(n_154), .B1(n_143), .B2(n_141), .Y(n_181) );
BUFx2_ASAP7_75t_L g182 ( .A(n_154), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_142), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_155), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_131), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_155), .Y(n_186) );
CKINVDCx16_ASAP7_75t_R g187 ( .A(n_154), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_154), .A2(n_86), .B1(n_119), .B2(n_96), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_169), .Y(n_189) );
INVx5_ASAP7_75t_L g190 ( .A(n_176), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_176), .Y(n_191) );
AND2x2_ASAP7_75t_SL g192 ( .A(n_175), .B(n_155), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_169), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_176), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_159), .B(n_154), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_169), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g197 ( .A1(n_183), .A2(n_142), .B(n_141), .Y(n_197) );
BUFx2_ASAP7_75t_L g198 ( .A(n_175), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_171), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_166), .B(n_155), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_SL g201 ( .A1(n_173), .A2(n_142), .B(n_147), .C(n_140), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_171), .Y(n_202) );
INVx3_ASAP7_75t_L g203 ( .A(n_176), .Y(n_203) );
BUFx8_ASAP7_75t_SL g204 ( .A(n_164), .Y(n_204) );
CKINVDCx6p67_ASAP7_75t_R g205 ( .A(n_164), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_156), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_164), .A2(n_154), .B1(n_136), .B2(n_137), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_162), .A2(n_136), .B(n_140), .C(n_147), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_164), .A2(n_137), .B1(n_119), .B2(n_133), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_171), .Y(n_210) );
CKINVDCx6p67_ASAP7_75t_R g211 ( .A(n_187), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_159), .B(n_121), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_158), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_160), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_177), .B(n_159), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_166), .A2(n_126), .B1(n_123), .B2(n_124), .Y(n_216) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_179), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_174), .B(n_125), .Y(n_218) );
AND2x2_ASAP7_75t_SL g219 ( .A(n_156), .B(n_170), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_161), .Y(n_220) );
OAI211xp5_ASAP7_75t_L g221 ( .A1(n_215), .A2(n_188), .B(n_168), .C(n_181), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_189), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_190), .B(n_172), .Y(n_223) );
INVx3_ASAP7_75t_SL g224 ( .A(n_211), .Y(n_224) );
BUFx3_ASAP7_75t_L g225 ( .A(n_190), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_207), .A2(n_178), .B1(n_172), .B2(n_156), .Y(n_226) );
OAI22xp33_ASAP7_75t_L g227 ( .A1(n_205), .A2(n_178), .B1(n_182), .B2(n_157), .Y(n_227) );
NAND2xp33_ASAP7_75t_L g228 ( .A(n_190), .B(n_185), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_192), .A2(n_186), .B1(n_184), .B2(n_163), .Y(n_229) );
AND2x2_ASAP7_75t_SL g230 ( .A(n_219), .B(n_165), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_201), .A2(n_183), .B(n_165), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_190), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_213), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_218), .B(n_182), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_198), .Y(n_235) );
OAI22xp33_ASAP7_75t_L g236 ( .A1(n_205), .A2(n_180), .B1(n_167), .B2(n_126), .Y(n_236) );
BUFx2_ASAP7_75t_L g237 ( .A(n_198), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_189), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_190), .B(n_185), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_190), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_200), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_213), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_192), .A2(n_94), .B1(n_127), .B2(n_124), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_192), .A2(n_120), .B1(n_123), .B2(n_124), .Y(n_244) );
AOI21xp5_ASAP7_75t_R g245 ( .A1(n_204), .A2(n_105), .B(n_117), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_207), .A2(n_120), .B1(n_127), .B2(n_123), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_234), .B(n_212), .Y(n_247) );
AOI221xp5_ASAP7_75t_L g248 ( .A1(n_221), .A2(n_217), .B1(n_208), .B2(n_214), .C(n_220), .Y(n_248) );
OAI21xp33_ASAP7_75t_SL g249 ( .A1(n_230), .A2(n_219), .B(n_216), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_240), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_234), .B(n_200), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_229), .A2(n_219), .B1(n_216), .B2(n_209), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_230), .A2(n_200), .B1(n_195), .B2(n_211), .Y(n_253) );
OAI221xp5_ASAP7_75t_L g254 ( .A1(n_243), .A2(n_220), .B1(n_214), .B2(n_197), .C(n_193), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_244), .A2(n_200), .B1(n_191), .B2(n_194), .Y(n_255) );
OAI211xp5_ASAP7_75t_L g256 ( .A1(n_244), .A2(n_106), .B(n_79), .C(n_85), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_235), .B(n_193), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_229), .A2(n_191), .B1(n_194), .B2(n_199), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_235), .B(n_196), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_233), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_224), .Y(n_261) );
AOI221xp5_ASAP7_75t_L g262 ( .A1(n_236), .A2(n_97), .B1(n_124), .B2(n_123), .C(n_120), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_233), .Y(n_263) );
OAI221xp5_ASAP7_75t_L g264 ( .A1(n_237), .A2(n_202), .B1(n_199), .B2(n_196), .C(n_123), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_242), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_230), .A2(n_202), .B1(n_210), .B2(n_203), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_225), .Y(n_267) );
AOI221xp5_ASAP7_75t_L g268 ( .A1(n_248), .A2(n_246), .B1(n_242), .B2(n_237), .C(n_79), .Y(n_268) );
AOI221xp5_ASAP7_75t_L g269 ( .A1(n_256), .A2(n_107), .B1(n_106), .B2(n_85), .C(n_87), .Y(n_269) );
INVx1_ASAP7_75t_SL g270 ( .A(n_261), .Y(n_270) );
NAND3xp33_ASAP7_75t_L g271 ( .A(n_249), .B(n_231), .C(n_128), .Y(n_271) );
AOI221xp5_ASAP7_75t_L g272 ( .A1(n_262), .A2(n_252), .B1(n_249), .B2(n_260), .C(n_263), .Y(n_272) );
OAI211xp5_ASAP7_75t_L g273 ( .A1(n_260), .A2(n_87), .B(n_100), .C(n_92), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_252), .A2(n_226), .B1(n_227), .B2(n_241), .Y(n_274) );
OAI33xp33_ASAP7_75t_L g275 ( .A1(n_263), .A2(n_100), .A3(n_103), .B1(n_104), .B2(n_113), .B3(n_129), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_247), .B(n_224), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_265), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_265), .Y(n_278) );
INVxp67_ASAP7_75t_L g279 ( .A(n_261), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_247), .B(n_224), .Y(n_280) );
BUFx2_ASAP7_75t_L g281 ( .A(n_250), .Y(n_281) );
AOI21xp5_ASAP7_75t_SL g282 ( .A1(n_258), .A2(n_225), .B(n_240), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_254), .A2(n_130), .B1(n_129), .B2(n_113), .C(n_124), .Y(n_283) );
AO21x2_ASAP7_75t_L g284 ( .A1(n_266), .A2(n_113), .B(n_129), .Y(n_284) );
AOI211x1_ASAP7_75t_L g285 ( .A1(n_264), .A2(n_245), .B(n_4), .C(n_5), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_250), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_267), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_251), .B(n_222), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_251), .A2(n_241), .B1(n_225), .B2(n_120), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_286), .Y(n_290) );
OR2x6_ASAP7_75t_L g291 ( .A(n_282), .B(n_267), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_281), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_277), .B(n_250), .Y(n_293) );
AND2x2_ASAP7_75t_SL g294 ( .A(n_274), .B(n_223), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_276), .B(n_257), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_286), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_271), .B(n_240), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_272), .A2(n_268), .B1(n_274), .B2(n_275), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_278), .Y(n_299) );
NAND3xp33_ASAP7_75t_L g300 ( .A(n_285), .B(n_273), .C(n_269), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_277), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_278), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_281), .B(n_259), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_286), .Y(n_304) );
AOI33xp33_ASAP7_75t_L g305 ( .A1(n_270), .A2(n_113), .A3(n_129), .B1(n_130), .B2(n_253), .B3(n_152), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_284), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_288), .B(n_130), .Y(n_307) );
AOI211xp5_ASAP7_75t_L g308 ( .A1(n_282), .A2(n_255), .B(n_75), .C(n_102), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_288), .B(n_130), .Y(n_309) );
OAI221xp5_ASAP7_75t_L g310 ( .A1(n_271), .A2(n_241), .B1(n_127), .B2(n_120), .C(n_232), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_284), .B(n_222), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_284), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_287), .B(n_240), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_280), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_279), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_285), .B(n_240), .Y(n_316) );
OAI33xp33_ASAP7_75t_L g317 ( .A1(n_283), .A2(n_3), .A3(n_4), .B1(n_5), .B2(n_6), .B3(n_7), .Y(n_317) );
INVx3_ASAP7_75t_R g318 ( .A(n_289), .Y(n_318) );
NOR2xp67_ASAP7_75t_SL g319 ( .A(n_282), .B(n_240), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_272), .A2(n_241), .B1(n_128), .B2(n_238), .Y(n_320) );
NAND4xp25_ASAP7_75t_L g321 ( .A(n_308), .B(n_127), .C(n_134), .D(n_145), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_314), .B(n_7), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_302), .B(n_128), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_314), .B(n_9), .Y(n_324) );
OAI33xp33_ASAP7_75t_L g325 ( .A1(n_300), .A2(n_10), .A3(n_11), .B1(n_12), .B2(n_13), .B3(n_14), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_307), .B(n_128), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_294), .A2(n_128), .B1(n_238), .B2(n_127), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_302), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_299), .Y(n_329) );
INVx1_ASAP7_75t_SL g330 ( .A(n_315), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_299), .Y(n_331) );
OAI221xp5_ASAP7_75t_L g332 ( .A1(n_300), .A2(n_128), .B1(n_232), .B2(n_108), .C(n_210), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_294), .A2(n_128), .B1(n_232), .B2(n_108), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_303), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_307), .B(n_11), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_291), .B(n_108), .Y(n_337) );
INVx1_ASAP7_75t_SL g338 ( .A(n_315), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_294), .A2(n_108), .B1(n_223), .B2(n_117), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_307), .B(n_12), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_309), .B(n_13), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_293), .B(n_14), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_293), .B(n_15), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_293), .B(n_16), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_298), .A2(n_223), .B1(n_239), .B2(n_210), .Y(n_345) );
NOR2x1_ASAP7_75t_L g346 ( .A(n_315), .B(n_228), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_301), .Y(n_347) );
NOR4xp75_ASAP7_75t_L g348 ( .A(n_316), .B(n_18), .C(n_19), .D(n_203), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_309), .B(n_18), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_318), .B(n_23), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_292), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_311), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_309), .B(n_239), .Y(n_353) );
INVx1_ASAP7_75t_SL g354 ( .A(n_313), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_295), .B(n_239), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_298), .B(n_117), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_292), .B(n_153), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_311), .Y(n_358) );
NAND2x1p5_ASAP7_75t_L g359 ( .A(n_346), .B(n_319), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_329), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_332), .A2(n_310), .B(n_297), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_334), .B(n_306), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_330), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_331), .Y(n_364) );
NOR2xp67_ASAP7_75t_SL g365 ( .A(n_324), .B(n_310), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_352), .B(n_312), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_335), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_358), .B(n_313), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_338), .Y(n_369) );
NAND2xp33_ASAP7_75t_SL g370 ( .A(n_351), .B(n_319), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_328), .Y(n_371) );
OAI21xp5_ASAP7_75t_SL g372 ( .A1(n_322), .A2(n_320), .B(n_297), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_353), .B(n_304), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_322), .B(n_318), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_342), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_342), .B(n_304), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_343), .B(n_313), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_347), .B(n_297), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_354), .B(n_297), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_343), .B(n_313), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_344), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_323), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_323), .Y(n_383) );
INVx1_ASAP7_75t_SL g384 ( .A(n_355), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_325), .B(n_317), .Y(n_385) );
AO22x2_ASAP7_75t_L g386 ( .A1(n_337), .A2(n_297), .B1(n_296), .B2(n_290), .Y(n_386) );
XNOR2x2_ASAP7_75t_L g387 ( .A(n_348), .B(n_291), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_336), .B(n_320), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_340), .B(n_296), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_337), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_350), .B(n_317), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_341), .B(n_296), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_326), .B(n_296), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_333), .B(n_290), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_349), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_357), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_333), .B(n_290), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_327), .B(n_305), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_350), .B(n_291), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_327), .B(n_291), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_363), .B(n_291), .Y(n_401) );
OAI211xp5_ASAP7_75t_L g402 ( .A1(n_374), .A2(n_321), .B(n_339), .C(n_356), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_360), .Y(n_403) );
INVx3_ASAP7_75t_L g404 ( .A(n_386), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_364), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_369), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_375), .B(n_345), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_381), .B(n_339), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_396), .Y(n_409) );
XOR2x2_ASAP7_75t_L g410 ( .A(n_374), .B(n_24), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_370), .B(n_134), .Y(n_411) );
OAI222xp33_ASAP7_75t_L g412 ( .A1(n_365), .A2(n_203), .B1(n_149), .B2(n_145), .C1(n_134), .C2(n_206), .Y(n_412) );
INVx1_ASAP7_75t_SL g413 ( .A(n_376), .Y(n_413) );
XNOR2xp5_ASAP7_75t_L g414 ( .A(n_387), .B(n_27), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_386), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_370), .B(n_145), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_372), .A2(n_206), .B1(n_146), .B2(n_30), .Y(n_417) );
XOR2x2_ASAP7_75t_L g418 ( .A(n_387), .B(n_28), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_367), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_366), .B(n_395), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_391), .B(n_385), .Y(n_421) );
XOR2x2_ASAP7_75t_L g422 ( .A(n_391), .B(n_29), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_385), .B(n_32), .Y(n_423) );
XNOR2xp5_ASAP7_75t_L g424 ( .A(n_377), .B(n_34), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_362), .Y(n_425) );
O2A1O1Ixp33_ASAP7_75t_L g426 ( .A1(n_398), .A2(n_151), .B(n_135), .C(n_131), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_389), .B(n_35), .Y(n_427) );
XOR2x2_ASAP7_75t_SL g428 ( .A(n_359), .B(n_36), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_392), .B(n_40), .Y(n_429) );
AOI211xp5_ASAP7_75t_L g430 ( .A1(n_399), .A2(n_41), .B(n_43), .C(n_47), .Y(n_430) );
AND2x2_ASAP7_75t_SL g431 ( .A(n_399), .B(n_146), .Y(n_431) );
A2O1A1Ixp33_ASAP7_75t_L g432 ( .A1(n_361), .A2(n_50), .B(n_51), .C(n_54), .Y(n_432) );
AO22x1_ASAP7_75t_L g433 ( .A1(n_400), .A2(n_55), .B1(n_58), .B2(n_59), .Y(n_433) );
CKINVDCx14_ASAP7_75t_R g434 ( .A(n_373), .Y(n_434) );
AO22x2_ASAP7_75t_L g435 ( .A1(n_390), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_435) );
NAND5xp2_ASAP7_75t_L g436 ( .A(n_359), .B(n_65), .C(n_66), .D(n_67), .E(n_68), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_379), .B(n_69), .Y(n_437) );
AOI211xp5_ASAP7_75t_SL g438 ( .A1(n_388), .A2(n_70), .B(n_71), .C(n_131), .Y(n_438) );
OAI211xp5_ASAP7_75t_L g439 ( .A1(n_380), .A2(n_146), .B(n_135), .C(n_151), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_368), .Y(n_440) );
NAND3xp33_ASAP7_75t_L g441 ( .A(n_397), .B(n_185), .C(n_390), .Y(n_441) );
INVxp67_ASAP7_75t_L g442 ( .A(n_394), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_386), .A2(n_185), .B1(n_382), .B2(n_379), .Y(n_443) );
NOR2xp67_ASAP7_75t_SL g444 ( .A(n_393), .B(n_383), .Y(n_444) );
OAI21xp33_ASAP7_75t_SL g445 ( .A1(n_378), .A2(n_383), .B(n_371), .Y(n_445) );
AOI21xp33_ASAP7_75t_L g446 ( .A1(n_378), .A2(n_391), .B(n_385), .Y(n_446) );
AOI21xp33_ASAP7_75t_L g447 ( .A1(n_371), .A2(n_385), .B(n_391), .Y(n_447) );
AOI211xp5_ASAP7_75t_L g448 ( .A1(n_374), .A2(n_391), .B(n_372), .C(n_399), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_384), .B(n_375), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_360), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_384), .B(n_375), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_360), .Y(n_452) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_385), .A2(n_322), .B(n_391), .Y(n_453) );
AOI22x1_ASAP7_75t_SL g454 ( .A1(n_406), .A2(n_404), .B1(n_415), .B2(n_421), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_418), .A2(n_417), .B(n_411), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g456 ( .A1(n_421), .A2(n_453), .B(n_447), .C(n_446), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_440), .Y(n_457) );
INVxp67_ASAP7_75t_SL g458 ( .A(n_428), .Y(n_458) );
OAI211xp5_ASAP7_75t_L g459 ( .A1(n_448), .A2(n_447), .B(n_453), .C(n_423), .Y(n_459) );
NOR2x1_ASAP7_75t_L g460 ( .A(n_417), .B(n_414), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_423), .A2(n_422), .B1(n_408), .B2(n_410), .Y(n_461) );
NOR2x1_ASAP7_75t_L g462 ( .A(n_415), .B(n_404), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_409), .Y(n_463) );
OAI211xp5_ASAP7_75t_SL g464 ( .A1(n_445), .A2(n_402), .B(n_442), .C(n_443), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_425), .Y(n_465) );
NAND4xp25_ASAP7_75t_L g466 ( .A(n_436), .B(n_430), .C(n_438), .D(n_432), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_434), .A2(n_413), .B1(n_431), .B2(n_424), .Y(n_467) );
AOI22x1_ASAP7_75t_L g468 ( .A1(n_458), .A2(n_435), .B1(n_438), .B2(n_437), .Y(n_468) );
OAI22xp5_ASAP7_75t_SL g469 ( .A1(n_458), .A2(n_431), .B1(n_441), .B2(n_427), .Y(n_469) );
NAND4xp25_ASAP7_75t_L g470 ( .A(n_460), .B(n_432), .C(n_427), .D(n_429), .Y(n_470) );
INVxp67_ASAP7_75t_SL g471 ( .A(n_463), .Y(n_471) );
OAI22x1_ASAP7_75t_L g472 ( .A1(n_463), .A2(n_416), .B1(n_411), .B2(n_405), .Y(n_472) );
NAND5xp2_ASAP7_75t_L g473 ( .A(n_455), .B(n_429), .C(n_426), .D(n_407), .E(n_439), .Y(n_473) );
OAI211xp5_ASAP7_75t_SL g474 ( .A1(n_459), .A2(n_420), .B(n_416), .C(n_451), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_456), .A2(n_419), .B1(n_403), .B2(n_450), .C(n_452), .Y(n_475) );
BUFx2_ASAP7_75t_L g476 ( .A(n_462), .Y(n_476) );
NAND3xp33_ASAP7_75t_SL g477 ( .A(n_476), .B(n_461), .C(n_467), .Y(n_477) );
NAND3xp33_ASAP7_75t_L g478 ( .A(n_468), .B(n_454), .C(n_464), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_471), .Y(n_479) );
NAND4xp25_ASAP7_75t_L g480 ( .A(n_473), .B(n_470), .C(n_461), .D(n_466), .Y(n_480) );
OR3x1_ASAP7_75t_L g481 ( .A(n_474), .B(n_465), .C(n_457), .Y(n_481) );
NOR2x1_ASAP7_75t_L g482 ( .A(n_480), .B(n_412), .Y(n_482) );
AOI22xp5_ASAP7_75t_SL g483 ( .A1(n_479), .A2(n_472), .B1(n_433), .B2(n_469), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_477), .B(n_475), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_482), .Y(n_485) );
OAI222xp33_ASAP7_75t_L g486 ( .A1(n_484), .A2(n_481), .B1(n_478), .B2(n_444), .C1(n_449), .C2(n_401), .Y(n_486) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_485), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_487), .A2(n_485), .B(n_483), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_488), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_489), .A2(n_486), .B(n_487), .Y(n_490) );
endmodule