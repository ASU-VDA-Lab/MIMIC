module fake_jpeg_19373_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx11_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_11),
.B(n_23),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_0),
.B(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_68),
.Y(n_76)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_73),
.Y(n_90)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_59),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_70),
.A2(n_43),
.B1(n_62),
.B2(n_44),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_77),
.A2(n_81),
.B1(n_59),
.B2(n_60),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_52),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_52),
.B(n_55),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_47),
.B1(n_54),
.B2(n_51),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_68),
.C(n_64),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_87),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_94),
.B1(n_3),
.B2(n_4),
.Y(n_106)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_77),
.B1(n_79),
.B2(n_48),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_89),
.B1(n_50),
.B2(n_46),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_61),
.B1(n_49),
.B2(n_53),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_83),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_92),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_0),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_61),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_95),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_64),
.B1(n_50),
.B2(n_46),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_1),
.B(n_2),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_99),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_45),
.B1(n_17),
.B2(n_21),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_1),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_94),
.A2(n_14),
.B1(n_33),
.B2(n_31),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_104),
.Y(n_111)
);

AO22x2_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_30),
.B1(n_28),
.B2(n_27),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_102),
.A2(n_108),
.B(n_6),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_2),
.C(n_3),
.Y(n_104)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_4),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_109),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_38),
.B(n_25),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_117),
.Y(n_119)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

AO21x1_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_117),
.B(n_119),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_111),
.B1(n_116),
.B2(n_112),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_105),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_121),
.B1(n_103),
.B2(n_98),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_98),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_127),
.A2(n_115),
.B1(n_107),
.B2(n_102),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_102),
.A3(n_22),
.B1(n_12),
.B2(n_9),
.C1(n_6),
.C2(n_8),
.Y(n_129)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_129),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_7),
.Y(n_131)
);


endmodule