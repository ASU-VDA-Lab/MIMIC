module fake_netlist_1_5214_n_547 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_547);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_547;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_35), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_65), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_3), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_75), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_30), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_54), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_26), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_60), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_1), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_72), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_69), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_22), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_47), .Y(n_90) );
HB1xp67_ASAP7_75t_L g91 ( .A(n_41), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_70), .Y(n_92) );
BUFx3_ASAP7_75t_L g93 ( .A(n_8), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_44), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_5), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_38), .Y(n_96) );
OR2x2_ASAP7_75t_L g97 ( .A(n_34), .B(n_56), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_32), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_67), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_36), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_6), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_37), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_11), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_74), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_8), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_66), .Y(n_106) );
BUFx2_ASAP7_75t_L g107 ( .A(n_51), .Y(n_107) );
BUFx10_ASAP7_75t_L g108 ( .A(n_68), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_19), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_25), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_52), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_55), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_45), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
AND2x4_ASAP7_75t_L g115 ( .A(n_107), .B(n_0), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_81), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_85), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_85), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_88), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_107), .B(n_0), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_91), .B(n_1), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_96), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_86), .A2(n_103), .B1(n_80), .B2(n_114), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_81), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_96), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_87), .Y(n_126) );
BUFx8_ASAP7_75t_L g127 ( .A(n_97), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_88), .Y(n_128) );
NAND2xp33_ASAP7_75t_L g129 ( .A(n_79), .B(n_77), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_87), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_78), .B(n_2), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_89), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_89), .Y(n_133) );
BUFx8_ASAP7_75t_L g134 ( .A(n_97), .Y(n_134) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_90), .A2(n_29), .B(n_73), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_104), .Y(n_136) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_90), .A2(n_28), .B(n_71), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_127), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_117), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_117), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_118), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_118), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
AOI22xp33_ASAP7_75t_L g144 ( .A1(n_116), .A2(n_114), .B1(n_101), .B2(n_95), .Y(n_144) );
OR2x6_ASAP7_75t_L g145 ( .A(n_115), .B(n_95), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_122), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_116), .B(n_109), .Y(n_147) );
INVx4_ASAP7_75t_L g148 ( .A(n_115), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_135), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_122), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_119), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_121), .B(n_108), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_125), .Y(n_153) );
INVx4_ASAP7_75t_L g154 ( .A(n_115), .Y(n_154) );
INVx5_ASAP7_75t_L g155 ( .A(n_119), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_127), .B(n_108), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_119), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_125), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_127), .B(n_108), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_136), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_124), .B(n_109), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_119), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_136), .Y(n_163) );
NAND2xp33_ASAP7_75t_L g164 ( .A(n_143), .B(n_124), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_152), .B(n_134), .Y(n_165) );
O2A1O1Ixp5_ASAP7_75t_L g166 ( .A1(n_148), .A2(n_121), .B(n_120), .C(n_126), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_152), .B(n_134), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_138), .Y(n_169) );
NOR2x2_ASAP7_75t_L g170 ( .A(n_145), .B(n_134), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_151), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_148), .B(n_126), .Y(n_172) );
OAI22xp33_ASAP7_75t_L g173 ( .A1(n_145), .A2(n_103), .B1(n_133), .B2(n_132), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_151), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_148), .B(n_130), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_148), .B(n_130), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_154), .B(n_132), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_154), .B(n_133), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_154), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_154), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_145), .B(n_131), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_145), .A2(n_123), .B1(n_129), .B2(n_93), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_139), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_156), .B(n_79), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_141), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_159), .B(n_82), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_145), .B(n_82), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_144), .A2(n_93), .B1(n_105), .B2(n_112), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_147), .A2(n_137), .B(n_135), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_147), .B(n_105), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_151), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_144), .A2(n_128), .B1(n_119), .B2(n_94), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_141), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_143), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_161), .B(n_112), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_161), .B(n_84), .Y(n_196) );
NOR2xp67_ASAP7_75t_L g197 ( .A(n_140), .B(n_128), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_164), .A2(n_143), .B(n_149), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_173), .A2(n_146), .B1(n_140), .B2(n_160), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_172), .A2(n_143), .B(n_149), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_167), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_167), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_190), .B(n_142), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_170), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_183), .Y(n_205) );
OAI21xp33_ASAP7_75t_SL g206 ( .A1(n_183), .A2(n_163), .B(n_142), .Y(n_206) );
AOI22xp33_ASAP7_75t_SL g207 ( .A1(n_165), .A2(n_84), .B1(n_160), .B2(n_140), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_190), .B(n_150), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_181), .A2(n_168), .B1(n_182), .B2(n_195), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_185), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_196), .B(n_150), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_166), .A2(n_163), .B(n_153), .C(n_158), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_172), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_188), .B(n_153), .Y(n_214) );
BUFx12f_ASAP7_75t_L g215 ( .A(n_169), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_181), .A2(n_158), .B(n_160), .C(n_146), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_175), .A2(n_140), .B(n_160), .C(n_146), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_176), .A2(n_146), .B(n_92), .C(n_106), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_177), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_185), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_184), .B(n_149), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_193), .Y(n_222) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_193), .B(n_135), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_194), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_194), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_178), .A2(n_100), .B(n_92), .C(n_94), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_187), .A2(n_106), .B(n_100), .C(n_113), .Y(n_227) );
NAND2x1p5_ASAP7_75t_L g228 ( .A(n_179), .B(n_137), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_188), .B(n_149), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_194), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_SL g231 ( .A1(n_229), .A2(n_189), .B(n_186), .C(n_99), .Y(n_231) );
OAI22xp33_ASAP7_75t_L g232 ( .A1(n_204), .A2(n_169), .B1(n_179), .B2(n_180), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_213), .B(n_180), .Y(n_233) );
INVxp67_ASAP7_75t_L g234 ( .A(n_203), .Y(n_234) );
OAI22xp33_ASAP7_75t_SL g235 ( .A1(n_204), .A2(n_113), .B1(n_189), .B2(n_102), .Y(n_235) );
AOI21x1_ASAP7_75t_L g236 ( .A1(n_200), .A2(n_198), .B(n_225), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_201), .B(n_192), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_201), .Y(n_238) );
NOR2xp33_ASAP7_75t_SL g239 ( .A(n_224), .B(n_194), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_205), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_205), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_209), .B(n_143), .Y(n_242) );
AO31x2_ASAP7_75t_L g243 ( .A1(n_202), .A2(n_162), .A3(n_157), .B(n_104), .Y(n_243) );
OAI21x1_ASAP7_75t_L g244 ( .A1(n_228), .A2(n_137), .B(n_191), .Y(n_244) );
AOI31xp67_ASAP7_75t_L g245 ( .A1(n_225), .A2(n_157), .A3(n_162), .B(n_191), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_202), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_206), .A2(n_197), .B(n_149), .C(n_143), .Y(n_247) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_230), .A2(n_162), .B(n_157), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_210), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_227), .A2(n_197), .B(n_149), .C(n_83), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_210), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_220), .Y(n_252) );
BUFx2_ASAP7_75t_L g253 ( .A(n_208), .Y(n_253) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_230), .A2(n_98), .B(n_110), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_220), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_219), .B(n_194), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_222), .A2(n_111), .B(n_171), .C(n_174), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_249), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_234), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_239), .A2(n_224), .B(n_221), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_246), .B(n_222), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_238), .A2(n_216), .B(n_226), .C(n_218), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_240), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_246), .B(n_214), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_249), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_253), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_240), .Y(n_267) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_238), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_253), .B(n_207), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_251), .B(n_211), .Y(n_270) );
OA21x2_ASAP7_75t_L g271 ( .A1(n_247), .A2(n_199), .B(n_171), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_239), .A2(n_224), .B(n_217), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_235), .A2(n_215), .B1(n_228), .B2(n_128), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_251), .B(n_212), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_242), .A2(n_224), .B(n_228), .Y(n_275) );
INVx1_ASAP7_75t_SL g276 ( .A(n_241), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_255), .B(n_223), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_255), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_241), .B(n_215), .Y(n_279) );
OAI221xp5_ASAP7_75t_L g280 ( .A1(n_250), .A2(n_223), .B1(n_128), .B2(n_137), .C(n_174), .Y(n_280) );
INVx3_ASAP7_75t_L g281 ( .A(n_268), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_266), .A2(n_235), .B1(n_252), .B2(n_232), .Y(n_282) );
AO21x2_ASAP7_75t_L g283 ( .A1(n_280), .A2(n_231), .B(n_236), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_258), .B(n_252), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_276), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_276), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_258), .B(n_243), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_266), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_265), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_259), .B(n_233), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_269), .A2(n_233), .B1(n_237), .B2(n_256), .Y(n_291) );
OA21x2_ASAP7_75t_L g292 ( .A1(n_275), .A2(n_244), .B(n_236), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_265), .Y(n_293) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_260), .A2(n_244), .B(n_223), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_278), .Y(n_295) );
OA21x2_ASAP7_75t_L g296 ( .A1(n_272), .A2(n_245), .B(n_237), .Y(n_296) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_274), .A2(n_257), .B(n_245), .Y(n_297) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_274), .A2(n_254), .B(n_243), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_278), .Y(n_299) );
AO21x2_ASAP7_75t_L g300 ( .A1(n_264), .A2(n_254), .B(n_243), .Y(n_300) );
INVxp67_ASAP7_75t_L g301 ( .A(n_266), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_261), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_290), .B(n_264), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_289), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_289), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_282), .B(n_273), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_289), .B(n_261), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_293), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_290), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_294), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_287), .B(n_277), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_293), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_281), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_287), .B(n_277), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_292), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_293), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_288), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_281), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_299), .B(n_270), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_299), .B(n_279), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_295), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_282), .A2(n_262), .B1(n_268), .B2(n_267), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_295), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_295), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_286), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_292), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_287), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_284), .B(n_267), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_284), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_284), .B(n_267), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_281), .B(n_243), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_302), .B(n_267), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_305), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_304), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_327), .B(n_298), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_303), .B(n_302), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_331), .B(n_281), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_305), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_309), .B(n_291), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_308), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_304), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_327), .B(n_291), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_312), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_311), .B(n_285), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_320), .B(n_288), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_317), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_331), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_308), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_311), .B(n_314), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_331), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_314), .B(n_298), .Y(n_351) );
AND2x4_ASAP7_75t_SL g352 ( .A(n_328), .B(n_285), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_314), .B(n_298), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_312), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_314), .B(n_298), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_329), .B(n_298), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_321), .B(n_286), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_316), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_329), .B(n_288), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_316), .B(n_328), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_321), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_323), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_323), .Y(n_363) );
NAND2x1_ASAP7_75t_L g364 ( .A(n_324), .B(n_281), .Y(n_364) );
CKINVDCx16_ASAP7_75t_R g365 ( .A(n_330), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_324), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_325), .Y(n_367) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_307), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_330), .B(n_286), .Y(n_369) );
NOR2x1_ASAP7_75t_L g370 ( .A(n_307), .B(n_300), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_325), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_319), .B(n_301), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_315), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_332), .B(n_301), .Y(n_374) );
NAND2x1_ASAP7_75t_L g375 ( .A(n_331), .B(n_268), .Y(n_375) );
NAND2xp33_ASAP7_75t_L g376 ( .A(n_322), .B(n_268), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_365), .B(n_332), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_344), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_365), .Y(n_379) );
NAND2xp33_ASAP7_75t_L g380 ( .A(n_370), .B(n_306), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_344), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_373), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_368), .B(n_326), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_349), .B(n_326), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_349), .B(n_318), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_334), .Y(n_386) );
INVx2_ASAP7_75t_SL g387 ( .A(n_346), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_376), .A2(n_300), .B(n_326), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_336), .B(n_315), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_339), .B(n_315), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_373), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_334), .Y(n_392) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_346), .B(n_310), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_351), .B(n_318), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_335), .B(n_300), .Y(n_395) );
NAND2xp33_ASAP7_75t_L g396 ( .A(n_370), .B(n_268), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_360), .B(n_318), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_351), .B(n_318), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_335), .B(n_300), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_353), .B(n_313), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_353), .B(n_313), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_355), .B(n_313), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_341), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_355), .B(n_360), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_372), .B(n_313), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_341), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_345), .B(n_300), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_374), .B(n_296), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_356), .B(n_297), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_343), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_361), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_343), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_356), .B(n_297), .Y(n_413) );
NAND2x1_ASAP7_75t_L g414 ( .A(n_350), .B(n_310), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_359), .B(n_296), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_361), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_362), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_354), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_364), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_350), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_342), .B(n_297), .Y(n_421) );
NOR2x2_ASAP7_75t_L g422 ( .A(n_362), .B(n_310), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_369), .B(n_296), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_354), .Y(n_424) );
AND2x4_ASAP7_75t_SL g425 ( .A(n_337), .B(n_268), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_369), .B(n_297), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_363), .B(n_297), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_363), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_378), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_381), .B(n_366), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_379), .B(n_347), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_404), .B(n_352), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_420), .A2(n_347), .B1(n_352), .B2(n_375), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_387), .Y(n_434) );
INVx2_ASAP7_75t_SL g435 ( .A(n_387), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_420), .B(n_394), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_390), .B(n_366), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_386), .Y(n_438) );
INVxp67_ASAP7_75t_L g439 ( .A(n_389), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_384), .B(n_352), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_408), .B(n_367), .Y(n_441) );
AOI222xp33_ASAP7_75t_L g442 ( .A1(n_380), .A2(n_347), .B1(n_371), .B2(n_367), .C1(n_337), .C2(n_333), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_407), .B(n_371), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_416), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_385), .B(n_337), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_392), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_415), .B(n_338), .Y(n_447) );
AOI222xp33_ASAP7_75t_L g448 ( .A1(n_380), .A2(n_337), .B1(n_333), .B2(n_358), .C1(n_338), .C2(n_340), .Y(n_448) );
NOR2x1_ASAP7_75t_L g449 ( .A(n_393), .B(n_364), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_398), .B(n_375), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_383), .B(n_357), .Y(n_451) );
INVx1_ASAP7_75t_SL g452 ( .A(n_422), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_400), .B(n_358), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_401), .B(n_402), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_419), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_377), .B(n_348), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_395), .B(n_348), .Y(n_457) );
NOR2xp67_ASAP7_75t_L g458 ( .A(n_419), .B(n_357), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_405), .B(n_2), .Y(n_459) );
NOR2x1_ASAP7_75t_L g460 ( .A(n_393), .B(n_340), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_403), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_423), .B(n_296), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_405), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_397), .B(n_310), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_406), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_399), .B(n_410), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_412), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_416), .B(n_296), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_428), .B(n_296), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_428), .B(n_310), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_418), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_424), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_422), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_441), .Y(n_474) );
OAI22xp33_ASAP7_75t_L g475 ( .A1(n_452), .A2(n_419), .B1(n_414), .B2(n_388), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_430), .Y(n_476) );
NAND2xp33_ASAP7_75t_L g477 ( .A(n_452), .B(n_426), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_437), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_437), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_438), .Y(n_480) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_466), .A2(n_409), .B1(n_413), .B2(n_421), .C(n_427), .Y(n_481) );
AND4x1_ASAP7_75t_L g482 ( .A(n_442), .B(n_3), .C(n_4), .D(n_5), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_439), .B(n_417), .Y(n_483) );
AOI21xp33_ASAP7_75t_L g484 ( .A1(n_459), .A2(n_396), .B(n_382), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_463), .A2(n_396), .B1(n_417), .B2(n_411), .Y(n_485) );
INVxp67_ASAP7_75t_SL g486 ( .A(n_444), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_429), .B(n_411), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_446), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_468), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_443), .B(n_391), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_458), .A2(n_391), .B(n_382), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_461), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_462), .B(n_425), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_431), .A2(n_425), .B1(n_263), .B2(n_292), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_465), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_467), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_471), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_457), .B(n_283), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_442), .A2(n_254), .B(n_263), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_457), .B(n_283), .Y(n_500) );
AOI211xp5_ASAP7_75t_L g501 ( .A1(n_433), .A2(n_128), .B(n_294), .C(n_263), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_447), .B(n_451), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_469), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_478), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_475), .A2(n_435), .B(n_434), .C(n_455), .Y(n_505) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_486), .A2(n_473), .B1(n_433), .B2(n_455), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_481), .B(n_448), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_474), .B(n_436), .Y(n_508) );
AOI322xp5_ASAP7_75t_L g509 ( .A1(n_475), .A2(n_431), .A3(n_432), .B1(n_436), .B2(n_456), .C1(n_440), .C2(n_454), .Y(n_509) );
OAI222xp33_ASAP7_75t_L g510 ( .A1(n_493), .A2(n_449), .B1(n_450), .B2(n_460), .C1(n_445), .C2(n_472), .Y(n_510) );
AOI322xp5_ASAP7_75t_L g511 ( .A1(n_477), .A2(n_453), .A3(n_464), .B1(n_448), .B2(n_263), .C1(n_470), .C2(n_11), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g512 ( .A1(n_481), .A2(n_283), .B1(n_155), .B2(n_7), .C(n_9), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g513 ( .A1(n_479), .A2(n_283), .B1(n_155), .B2(n_7), .C(n_9), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_476), .B(n_283), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_489), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_486), .A2(n_292), .B1(n_254), .B2(n_271), .Y(n_516) );
OAI221xp5_ASAP7_75t_L g517 ( .A1(n_482), .A2(n_292), .B1(n_271), .B2(n_155), .C(n_12), .Y(n_517) );
AOI222xp33_ASAP7_75t_L g518 ( .A1(n_498), .A2(n_4), .B1(n_6), .B2(n_10), .C1(n_12), .C2(n_13), .Y(n_518) );
AOI322xp5_ASAP7_75t_L g519 ( .A1(n_502), .A2(n_10), .A3(n_13), .B1(n_14), .B2(n_292), .C1(n_271), .C2(n_243), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_503), .B(n_271), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_501), .A2(n_248), .B1(n_155), .B2(n_294), .Y(n_521) );
AOI221xp5_ASAP7_75t_L g522 ( .A1(n_507), .A2(n_492), .B1(n_480), .B2(n_497), .C(n_496), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_509), .B(n_483), .Y(n_523) );
INVx1_ASAP7_75t_SL g524 ( .A(n_508), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g525 ( .A1(n_505), .A2(n_488), .B1(n_495), .B2(n_484), .C(n_494), .Y(n_525) );
NOR2xp33_ASAP7_75t_R g526 ( .A(n_504), .B(n_490), .Y(n_526) );
AOI221xp5_ASAP7_75t_L g527 ( .A1(n_506), .A2(n_491), .B1(n_487), .B2(n_500), .C(n_499), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_511), .B(n_485), .Y(n_528) );
NAND4xp75_ASAP7_75t_L g529 ( .A(n_512), .B(n_248), .C(n_16), .D(n_17), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_SL g530 ( .A1(n_517), .A2(n_15), .B(n_18), .C(n_20), .Y(n_530) );
OAI211xp5_ASAP7_75t_L g531 ( .A1(n_518), .A2(n_155), .B(n_248), .C(n_224), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_522), .B(n_518), .Y(n_532) );
NAND5xp2_ASAP7_75t_L g533 ( .A(n_531), .B(n_513), .C(n_519), .D(n_510), .E(n_514), .Y(n_533) );
NAND5xp2_ASAP7_75t_L g534 ( .A(n_523), .B(n_520), .C(n_521), .D(n_516), .E(n_27), .Y(n_534) );
NAND4xp25_ASAP7_75t_L g535 ( .A(n_528), .B(n_515), .C(n_23), .D(n_24), .Y(n_535) );
NAND5xp2_ASAP7_75t_L g536 ( .A(n_527), .B(n_21), .C(n_31), .D(n_33), .E(n_39), .Y(n_536) );
NAND4xp75_ASAP7_75t_L g537 ( .A(n_532), .B(n_525), .C(n_530), .D(n_526), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_533), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_535), .Y(n_539) );
OAI22xp5_ASAP7_75t_SL g540 ( .A1(n_538), .A2(n_524), .B1(n_534), .B2(n_536), .Y(n_540) );
OR3x2_ASAP7_75t_L g541 ( .A(n_537), .B(n_529), .C(n_42), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_540), .Y(n_542) );
OAI31xp33_ASAP7_75t_SL g543 ( .A1(n_542), .A2(n_541), .A3(n_539), .B(n_46), .Y(n_543) );
AOI222xp33_ASAP7_75t_L g544 ( .A1(n_543), .A2(n_539), .B1(n_155), .B2(n_48), .C1(n_49), .C2(n_50), .Y(n_544) );
AOI222xp33_ASAP7_75t_L g545 ( .A1(n_544), .A2(n_155), .B1(n_43), .B2(n_53), .C1(n_57), .C2(n_58), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_545), .A2(n_248), .B1(n_59), .B2(n_61), .Y(n_546) );
AOI222xp33_ASAP7_75t_L g547 ( .A1(n_546), .A2(n_40), .B1(n_62), .B2(n_63), .C1(n_64), .C2(n_76), .Y(n_547) );
endmodule