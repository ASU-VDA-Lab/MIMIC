module fake_jpeg_2753_n_158 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_36),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_62),
.Y(n_66)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_48),
.B1(n_56),
.B2(n_43),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_72),
.B1(n_74),
.B2(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_55),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_42),
.B(n_45),
.C(n_46),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_54),
.B(n_46),
.C(n_45),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_48),
.B1(n_47),
.B2(n_56),
.Y(n_72)
);

OR2x4_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_41),
.Y(n_73)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_59),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_52),
.B1(n_41),
.B2(n_42),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_77),
.B(n_80),
.Y(n_105)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_84),
.C(n_85),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_75),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_83),
.B1(n_60),
.B2(n_50),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_73),
.A2(n_63),
.B1(n_60),
.B2(n_47),
.Y(n_83)
);

BUFx4f_ASAP7_75t_SL g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_90),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_53),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_69),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_74),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_17),
.C(n_38),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_0),
.B(n_1),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_10),
.B(n_11),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_2),
.C(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_106),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_2),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_100),
.B(n_18),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_103),
.B1(n_7),
.B2(n_8),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_118),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_16),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_112),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_91),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_39),
.C(n_34),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_116),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_117),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_98),
.B(n_32),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_7),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_9),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_114),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_124),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_125),
.B1(n_92),
.B2(n_15),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_24),
.C(n_28),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_97),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_134),
.Y(n_141)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_120),
.A2(n_92),
.B(n_20),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_128),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_27),
.B1(n_30),
.B2(n_14),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_135),
.B1(n_131),
.B2(n_126),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_121),
.Y(n_134)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_116),
.Y(n_138)
);

A2O1A1O1Ixp25_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_110),
.B(n_124),
.C(n_133),
.D(n_130),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_143),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_128),
.C(n_131),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_147),
.Y(n_149)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_140),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_141),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_144),
.B1(n_147),
.B2(n_145),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_146),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_150),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_149),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_136),
.B(n_132),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g157 ( 
.A(n_156),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_129),
.Y(n_158)
);


endmodule