module fake_jpeg_22001_n_282 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_282);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_282;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_37),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_41),
.Y(n_53)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_26),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_61),
.Y(n_77)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_64),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_27),
.B1(n_33),
.B2(n_32),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_46),
.A2(n_47),
.B1(n_26),
.B2(n_22),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_39),
.B1(n_43),
.B2(n_42),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_27),
.B1(n_34),
.B2(n_29),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_58),
.B1(n_60),
.B2(n_42),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_27),
.B1(n_34),
.B2(n_29),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_51),
.B1(n_26),
.B2(n_22),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_27),
.B1(n_34),
.B2(n_29),
.Y(n_51)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_38),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_19),
.B1(n_22),
.B2(n_28),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_32),
.B(n_19),
.C(n_28),
.Y(n_60)
);

NAND2x1_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_23),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_65),
.B1(n_41),
.B2(n_38),
.Y(n_69)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_70),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_69),
.B(n_92),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

NOR4xp25_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_0),
.C(n_1),
.D(n_2),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_1),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_42),
.B1(n_19),
.B2(n_28),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_86),
.B1(n_101),
.B2(n_59),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_76),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_85),
.Y(n_102)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx2_ASAP7_75t_SL g126 ( 
.A(n_75),
.Y(n_126)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_78),
.B(n_81),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_79),
.B(n_87),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_88),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_41),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_89),
.B1(n_47),
.B2(n_55),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_38),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_65),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_24),
.B1(n_17),
.B2(n_25),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_95),
.B1(n_98),
.B2(n_100),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_21),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_94),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_44),
.B(n_37),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_46),
.A2(n_37),
.B1(n_23),
.B2(n_18),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_31),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_97),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_31),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_23),
.B1(n_18),
.B2(n_30),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_50),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_1),
.Y(n_127)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_23),
.B1(n_18),
.B2(n_21),
.Y(n_101)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_0),
.Y(n_104)
);

AOI221xp5_ASAP7_75t_L g154 ( 
.A1(n_104),
.A2(n_125),
.B1(n_99),
.B2(n_68),
.C(n_5),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_105),
.A2(n_113),
.B1(n_75),
.B2(n_68),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_90),
.B1(n_95),
.B2(n_88),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_54),
.C(n_2),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_123),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_54),
.A3(n_64),
.B1(n_62),
.B2(n_45),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_116),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_64),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_121),
.C(n_67),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_62),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_81),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_62),
.C(n_21),
.Y(n_121)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_70),
.B1(n_83),
.B2(n_73),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_129),
.A2(n_134),
.B1(n_153),
.B2(n_155),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_131),
.B1(n_145),
.B2(n_154),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_77),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_137),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_136),
.Y(n_183)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_94),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_140),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_158),
.B(n_103),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_116),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_141),
.Y(n_185)
);

BUFx8_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_142),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_78),
.Y(n_143)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_111),
.A2(n_98),
.B1(n_84),
.B2(n_81),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_92),
.Y(n_146)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_106),
.B(n_87),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_148),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_112),
.B(n_97),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_110),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_112),
.B(n_96),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_151),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_119),
.A2(n_67),
.B1(n_4),
.B2(n_5),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_125),
.C(n_108),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_123),
.B1(n_107),
.B2(n_7),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_122),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_121),
.B(n_115),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_174),
.B(n_175),
.Y(n_188)
);

XOR2x2_ASAP7_75t_SL g200 ( 
.A(n_164),
.B(n_186),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_166),
.A2(n_177),
.B1(n_155),
.B2(n_147),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_169),
.C(n_179),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_108),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_128),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_173),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_3),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_107),
.B(n_6),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_130),
.A2(n_107),
.B1(n_7),
.B2(n_8),
.Y(n_177)
);

A2O1A1O1Ixp25_ASAP7_75t_L g179 ( 
.A1(n_142),
.A2(n_137),
.B(n_144),
.C(n_153),
.D(n_145),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_142),
.A2(n_3),
.B(n_7),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_151),
.B(n_148),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_8),
.C(n_9),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_182),
.C(n_133),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_10),
.Y(n_182)
);

NAND2xp33_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_10),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_190),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_192),
.Y(n_217)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_135),
.Y(n_193)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_198),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_133),
.C(n_141),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_205),
.C(n_175),
.Y(n_227)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_150),
.B1(n_136),
.B2(n_138),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_204),
.B1(n_208),
.B2(n_209),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_185),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_202),
.Y(n_210)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_176),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_146),
.C(n_134),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_149),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_197),
.Y(n_214)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_178),
.B(n_165),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_220),
.C(n_226),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_173),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_168),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_208),
.B1(n_166),
.B2(n_177),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_199),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_179),
.B1(n_159),
.B2(n_162),
.Y(n_222)
);

XOR2x2_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_164),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_189),
.B(n_172),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_226),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_182),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_172),
.C(n_194),
.Y(n_236)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_228),
.B(n_229),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_210),
.B(n_184),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_188),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_232),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_213),
.B(n_184),
.Y(n_233)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_234),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_242),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_237),
.C(n_238),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_194),
.C(n_204),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_194),
.C(n_196),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_239),
.B(n_241),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_187),
.B1(n_198),
.B2(n_200),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_240),
.A2(n_222),
.B1(n_219),
.B2(n_227),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_181),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_218),
.Y(n_242)
);

NAND4xp25_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_223),
.C(n_221),
.D(n_200),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_243),
.A2(n_246),
.B1(n_14),
.B2(n_15),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_236),
.A2(n_225),
.B(n_219),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_216),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_254),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_253),
.B(n_232),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_173),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_231),
.C(n_212),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_258),
.Y(n_268)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_231),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_260),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_247),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_11),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_14),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_SL g267 ( 
.A(n_263),
.B(n_14),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_244),
.B(n_243),
.C(n_246),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_267),
.B1(n_263),
.B2(n_257),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_270),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_264),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_271),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_251),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_273),
.C(n_274),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_244),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_258),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_255),
.C(n_271),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_278),
.B(n_279),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_254),
.C(n_253),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_280),
.A2(n_275),
.B1(n_15),
.B2(n_16),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_16),
.Y(n_282)
);


endmodule