module real_aes_7935_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_725;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_385;
wire n_214;
wire n_275;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_103;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_168;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_1), .A2(n_132), .B(n_136), .C(n_217), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_2), .A2(n_166), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g492 ( .A(n_3), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_4), .B(n_233), .Y(n_252) );
AOI21xp33_ASAP7_75t_L g457 ( .A1(n_5), .A2(n_166), .B(n_458), .Y(n_457) );
AND2x6_ASAP7_75t_L g132 ( .A(n_6), .B(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g207 ( .A(n_7), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_8), .B(n_42), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_9), .A2(n_165), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_10), .B(n_144), .Y(n_219) );
INVx1_ASAP7_75t_L g462 ( .A(n_11), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_12), .B(n_247), .Y(n_517) );
INVx1_ASAP7_75t_L g152 ( .A(n_13), .Y(n_152) );
INVx1_ASAP7_75t_L g529 ( .A(n_14), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_15), .A2(n_142), .B(n_229), .C(n_231), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_16), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_17), .B(n_480), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_18), .B(n_166), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_19), .B(n_178), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_20), .A2(n_247), .B(n_262), .C(n_264), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_21), .B(n_233), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_22), .B(n_144), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_23), .A2(n_174), .B(n_231), .C(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_24), .B(n_144), .Y(n_143) );
CKINVDCx16_ASAP7_75t_R g183 ( .A(n_25), .Y(n_183) );
INVx1_ASAP7_75t_L g140 ( .A(n_26), .Y(n_140) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_27), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_28), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_29), .B(n_144), .Y(n_493) );
OAI22xp5_ASAP7_75t_SL g723 ( .A1(n_30), .A2(n_31), .B1(n_724), .B2(n_725), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_30), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_31), .Y(n_724) );
INVx1_ASAP7_75t_L g172 ( .A(n_32), .Y(n_172) );
INVx1_ASAP7_75t_L g471 ( .A(n_33), .Y(n_471) );
AOI222xp33_ASAP7_75t_L g115 ( .A1(n_34), .A2(n_116), .B1(n_723), .B2(n_726), .C1(n_729), .C2(n_730), .Y(n_115) );
INVx2_ASAP7_75t_L g130 ( .A(n_35), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_36), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_37), .A2(n_247), .B(n_248), .C(n_250), .Y(n_246) );
INVxp67_ASAP7_75t_L g173 ( .A(n_38), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_39), .A2(n_136), .B(n_139), .C(n_147), .Y(n_135) );
CKINVDCx14_ASAP7_75t_R g245 ( .A(n_40), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_41), .A2(n_132), .B(n_136), .C(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g470 ( .A(n_43), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_44), .A2(n_191), .B(n_205), .C(n_206), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_45), .B(n_144), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_46), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_47), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_48), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g260 ( .A(n_49), .Y(n_260) );
CKINVDCx16_ASAP7_75t_R g472 ( .A(n_50), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_51), .B(n_166), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_52), .A2(n_136), .B1(n_264), .B2(n_469), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_53), .Y(n_508) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_54), .Y(n_489) );
CKINVDCx14_ASAP7_75t_R g203 ( .A(n_55), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_56), .A2(n_205), .B(n_250), .C(n_461), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_57), .Y(n_545) );
INVx1_ASAP7_75t_L g459 ( .A(n_58), .Y(n_459) );
AOI222xp33_ASAP7_75t_SL g100 ( .A1(n_59), .A2(n_101), .B1(n_114), .B2(n_733), .C1(n_738), .C2(n_749), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_59), .A2(n_87), .B1(n_741), .B2(n_742), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_59), .Y(n_742) );
INVx1_ASAP7_75t_L g133 ( .A(n_60), .Y(n_133) );
INVx1_ASAP7_75t_L g151 ( .A(n_61), .Y(n_151) );
INVx1_ASAP7_75t_SL g249 ( .A(n_62), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_63), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_64), .B(n_233), .Y(n_266) );
INVx1_ASAP7_75t_L g186 ( .A(n_65), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_SL g479 ( .A1(n_66), .A2(n_250), .B(n_480), .C(n_481), .Y(n_479) );
INVxp67_ASAP7_75t_L g482 ( .A(n_67), .Y(n_482) );
INVx1_ASAP7_75t_L g105 ( .A(n_68), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_69), .A2(n_166), .B(n_202), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_70), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_71), .A2(n_166), .B(n_226), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_72), .Y(n_474) );
INVx1_ASAP7_75t_L g539 ( .A(n_73), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_74), .A2(n_165), .B(n_167), .Y(n_164) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_75), .Y(n_134) );
INVx1_ASAP7_75t_L g227 ( .A(n_76), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_77), .A2(n_132), .B(n_136), .C(n_541), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_78), .A2(n_166), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g230 ( .A(n_79), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_80), .B(n_141), .Y(n_505) );
INVx2_ASAP7_75t_L g149 ( .A(n_81), .Y(n_149) );
INVx1_ASAP7_75t_L g218 ( .A(n_82), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_83), .B(n_480), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_84), .A2(n_132), .B(n_136), .C(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_L g109 ( .A(n_85), .B(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g119 ( .A(n_85), .B(n_111), .Y(n_119) );
INVx2_ASAP7_75t_L g448 ( .A(n_85), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_86), .A2(n_136), .B(n_185), .C(n_193), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_87), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_88), .B(n_148), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_89), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_90), .A2(n_132), .B(n_136), .C(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_91), .Y(n_521) );
INVx1_ASAP7_75t_L g478 ( .A(n_92), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_93), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_94), .B(n_141), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_95), .B(n_156), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_96), .B(n_156), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_97), .B(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g263 ( .A(n_98), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_99), .A2(n_166), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
NAND2xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_107), .Y(n_102) );
NOR2xp33_ASAP7_75t_SL g103 ( .A(n_104), .B(n_106), .Y(n_103) );
INVx1_ASAP7_75t_SL g737 ( .A(n_104), .Y(n_737) );
INVx1_ASAP7_75t_L g736 ( .A(n_106), .Y(n_736) );
OA21x2_ASAP7_75t_L g750 ( .A1(n_106), .A2(n_737), .B(n_748), .Y(n_750) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_109), .Y(n_744) );
BUFx2_ASAP7_75t_L g748 ( .A(n_109), .Y(n_748) );
NOR2x2_ASAP7_75t_L g732 ( .A(n_110), .B(n_448), .Y(n_732) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g447 ( .A(n_111), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_120), .B1(n_445), .B2(n_449), .Y(n_116) );
OAI22x1_ASAP7_75t_L g726 ( .A1(n_117), .A2(n_445), .B1(n_727), .B2(n_728), .Y(n_726) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g727 ( .A(n_120), .Y(n_727) );
XOR2xp5_ASAP7_75t_L g739 ( .A(n_120), .B(n_740), .Y(n_739) );
OR4x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_335), .C(n_382), .D(n_422), .Y(n_120) );
NAND3xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_281), .C(n_310), .Y(n_121) );
AOI211xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_196), .B(n_234), .C(n_274), .Y(n_122) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_123), .A2(n_294), .B(n_311), .C(n_315), .Y(n_310) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_158), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_125), .B(n_273), .Y(n_272) );
INVx3_ASAP7_75t_SL g277 ( .A(n_125), .Y(n_277) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_125), .Y(n_289) );
AND2x4_ASAP7_75t_L g293 ( .A(n_125), .B(n_241), .Y(n_293) );
AND2x2_ASAP7_75t_L g304 ( .A(n_125), .B(n_181), .Y(n_304) );
OR2x2_ASAP7_75t_L g328 ( .A(n_125), .B(n_237), .Y(n_328) );
AND2x2_ASAP7_75t_L g341 ( .A(n_125), .B(n_242), .Y(n_341) );
AND2x2_ASAP7_75t_L g381 ( .A(n_125), .B(n_367), .Y(n_381) );
AND2x2_ASAP7_75t_L g388 ( .A(n_125), .B(n_351), .Y(n_388) );
AND2x2_ASAP7_75t_L g418 ( .A(n_125), .B(n_159), .Y(n_418) );
OR2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_153), .Y(n_125) );
O2A1O1Ixp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_134), .B(n_135), .C(n_148), .Y(n_126) );
OAI21xp5_ASAP7_75t_L g182 ( .A1(n_127), .A2(n_183), .B(n_184), .Y(n_182) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_127), .A2(n_215), .B(n_216), .Y(n_214) );
OAI22xp33_ASAP7_75t_L g467 ( .A1(n_127), .A2(n_176), .B1(n_468), .B2(n_472), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_127), .A2(n_489), .B(n_490), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_127), .A2(n_539), .B(n_540), .Y(n_538) );
NAND2x1p5_ASAP7_75t_L g127 ( .A(n_128), .B(n_132), .Y(n_127) );
AND2x4_ASAP7_75t_L g166 ( .A(n_128), .B(n_132), .Y(n_166) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
INVx1_ASAP7_75t_L g146 ( .A(n_129), .Y(n_146) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g137 ( .A(n_130), .Y(n_137) );
INVx1_ASAP7_75t_L g265 ( .A(n_130), .Y(n_265) );
INVx1_ASAP7_75t_L g138 ( .A(n_131), .Y(n_138) );
INVx3_ASAP7_75t_L g142 ( .A(n_131), .Y(n_142) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_131), .Y(n_144) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_131), .Y(n_175) );
INVx1_ASAP7_75t_L g480 ( .A(n_131), .Y(n_480) );
BUFx3_ASAP7_75t_L g147 ( .A(n_132), .Y(n_147) );
INVx4_ASAP7_75t_SL g176 ( .A(n_132), .Y(n_176) );
INVx5_ASAP7_75t_L g169 ( .A(n_136), .Y(n_169) );
AND2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx3_ASAP7_75t_L g192 ( .A(n_137), .Y(n_192) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_137), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_141), .B(n_143), .C(n_145), .Y(n_139) );
OAI22xp33_ASAP7_75t_L g171 ( .A1(n_141), .A2(n_172), .B1(n_173), .B2(n_174), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_141), .A2(n_492), .B(n_493), .C(n_494), .Y(n_491) );
INVx5_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_142), .B(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_142), .B(n_462), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_142), .B(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g205 ( .A(n_144), .Y(n_205) );
INVx4_ASAP7_75t_L g247 ( .A(n_144), .Y(n_247) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_146), .B(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g179 ( .A(n_148), .Y(n_179) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_148), .A2(n_201), .B(n_208), .Y(n_200) );
INVx1_ASAP7_75t_L g213 ( .A(n_148), .Y(n_213) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_148), .A2(n_524), .B(n_530), .Y(n_523) );
AND2x2_ASAP7_75t_SL g148 ( .A(n_149), .B(n_150), .Y(n_148) );
AND2x2_ASAP7_75t_L g157 ( .A(n_149), .B(n_150), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_155), .A2(n_182), .B(n_194), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_155), .B(n_221), .Y(n_220) );
INVx3_ASAP7_75t_L g233 ( .A(n_155), .Y(n_233) );
NOR2xp33_ASAP7_75t_SL g507 ( .A(n_155), .B(n_508), .Y(n_507) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_156), .Y(n_224) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_156), .A2(n_476), .B(n_483), .Y(n_475) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g163 ( .A(n_157), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_158), .B(n_345), .Y(n_357) );
AND2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_180), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_159), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g295 ( .A(n_159), .B(n_180), .Y(n_295) );
BUFx3_ASAP7_75t_L g303 ( .A(n_159), .Y(n_303) );
OR2x2_ASAP7_75t_L g324 ( .A(n_159), .B(n_199), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_159), .B(n_345), .Y(n_435) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_164), .B(n_177), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_161), .A2(n_238), .B(n_239), .Y(n_237) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_161), .A2(n_538), .B(n_544), .Y(n_537) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AOI21xp5_ASAP7_75t_SL g501 ( .A1(n_162), .A2(n_502), .B(n_503), .Y(n_501) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AO21x2_ASAP7_75t_L g466 ( .A1(n_163), .A2(n_467), .B(n_473), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_163), .B(n_474), .Y(n_473) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_163), .A2(n_488), .B(n_495), .Y(n_487) );
INVx1_ASAP7_75t_L g238 ( .A(n_164), .Y(n_238) );
BUFx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_SL g167 ( .A1(n_168), .A2(n_169), .B(n_170), .C(n_176), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_SL g202 ( .A1(n_169), .A2(n_176), .B(n_203), .C(n_204), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_SL g226 ( .A1(n_169), .A2(n_176), .B(n_227), .C(n_228), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_169), .A2(n_176), .B(n_245), .C(n_246), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_SL g259 ( .A1(n_169), .A2(n_176), .B(n_260), .C(n_261), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g458 ( .A1(n_169), .A2(n_176), .B(n_459), .C(n_460), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_169), .A2(n_176), .B(n_478), .C(n_479), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_169), .A2(n_176), .B(n_526), .C(n_527), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_174), .B(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_174), .B(n_263), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_174), .B(n_529), .Y(n_528) );
INVx4_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g188 ( .A(n_175), .Y(n_188) );
OAI22xp5_ASAP7_75t_SL g469 ( .A1(n_175), .A2(n_188), .B1(n_470), .B2(n_471), .Y(n_469) );
INVx1_ASAP7_75t_L g193 ( .A(n_176), .Y(n_193) );
INVx1_ASAP7_75t_L g239 ( .A(n_177), .Y(n_239) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_179), .B(n_195), .Y(n_194) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_179), .A2(n_513), .B(n_520), .Y(n_512) );
AND2x2_ASAP7_75t_L g240 ( .A(n_180), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g288 ( .A(n_180), .Y(n_288) );
AND2x2_ASAP7_75t_L g351 ( .A(n_180), .B(n_242), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g353 ( .A1(n_180), .A2(n_354), .B1(n_356), .B2(n_358), .C(n_359), .Y(n_353) );
AND2x2_ASAP7_75t_L g367 ( .A(n_180), .B(n_237), .Y(n_367) );
AND2x2_ASAP7_75t_L g393 ( .A(n_180), .B(n_277), .Y(n_393) );
INVx2_ASAP7_75t_SL g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g273 ( .A(n_181), .B(n_242), .Y(n_273) );
BUFx2_ASAP7_75t_L g407 ( .A(n_181), .Y(n_407) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_189), .C(n_190), .Y(n_185) );
O2A1O1Ixp5_ASAP7_75t_L g217 ( .A1(n_187), .A2(n_190), .B(n_218), .C(n_219), .Y(n_217) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_190), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_190), .A2(n_542), .B(n_543), .Y(n_541) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g231 ( .A(n_192), .Y(n_231) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OAI32xp33_ASAP7_75t_L g373 ( .A1(n_197), .A2(n_334), .A3(n_348), .B1(n_374), .B2(n_375), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_209), .Y(n_197) );
AND2x2_ASAP7_75t_L g314 ( .A(n_198), .B(n_256), .Y(n_314) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
OR2x2_ASAP7_75t_L g296 ( .A(n_199), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_199), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g368 ( .A(n_199), .B(n_256), .Y(n_368) );
AND2x2_ASAP7_75t_L g379 ( .A(n_199), .B(n_271), .Y(n_379) );
BUFx3_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
OR2x2_ASAP7_75t_L g280 ( .A(n_200), .B(n_257), .Y(n_280) );
AND2x2_ASAP7_75t_L g284 ( .A(n_200), .B(n_257), .Y(n_284) );
AND2x2_ASAP7_75t_L g319 ( .A(n_200), .B(n_270), .Y(n_319) );
AND2x2_ASAP7_75t_L g326 ( .A(n_200), .B(n_222), .Y(n_326) );
OAI211xp5_ASAP7_75t_L g331 ( .A1(n_200), .A2(n_277), .B(n_288), .C(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g385 ( .A(n_200), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_200), .B(n_211), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_209), .B(n_268), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_209), .B(n_284), .Y(n_374) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g279 ( .A(n_210), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_222), .Y(n_210) );
AND2x2_ASAP7_75t_L g271 ( .A(n_211), .B(n_223), .Y(n_271) );
OR2x2_ASAP7_75t_L g286 ( .A(n_211), .B(n_223), .Y(n_286) );
AND2x2_ASAP7_75t_L g309 ( .A(n_211), .B(n_270), .Y(n_309) );
INVx1_ASAP7_75t_L g313 ( .A(n_211), .Y(n_313) );
AND2x2_ASAP7_75t_L g332 ( .A(n_211), .B(n_269), .Y(n_332) );
OAI22xp33_ASAP7_75t_L g342 ( .A1(n_211), .A2(n_297), .B1(n_343), .B2(n_344), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_211), .B(n_385), .Y(n_409) );
AND2x2_ASAP7_75t_L g424 ( .A(n_211), .B(n_284), .Y(n_424) );
INVx4_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
BUFx3_ASAP7_75t_L g254 ( .A(n_212), .Y(n_254) );
AND2x2_ASAP7_75t_L g298 ( .A(n_212), .B(n_223), .Y(n_298) );
AND2x2_ASAP7_75t_L g300 ( .A(n_212), .B(n_256), .Y(n_300) );
AND3x2_ASAP7_75t_L g362 ( .A(n_212), .B(n_326), .C(n_363), .Y(n_362) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_220), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_213), .B(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_213), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_213), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g397 ( .A(n_222), .B(n_269), .Y(n_397) );
INVx1_ASAP7_75t_SL g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g256 ( .A(n_223), .B(n_257), .Y(n_256) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_223), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_223), .B(n_268), .Y(n_330) );
NAND3xp33_ASAP7_75t_L g437 ( .A(n_223), .B(n_309), .C(n_385), .Y(n_437) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_232), .Y(n_223) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_224), .A2(n_243), .B(n_252), .Y(n_242) );
OA21x2_ASAP7_75t_L g257 ( .A1(n_224), .A2(n_258), .B(n_266), .Y(n_257) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_233), .A2(n_457), .B(n_463), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_253), .B1(n_267), .B2(n_272), .Y(n_234) );
INVx1_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_240), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_237), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g349 ( .A(n_237), .Y(n_349) );
OAI31xp33_ASAP7_75t_L g365 ( .A1(n_240), .A2(n_366), .A3(n_367), .B(n_368), .Y(n_365) );
AND2x2_ASAP7_75t_L g390 ( .A(n_240), .B(n_277), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_240), .B(n_303), .Y(n_436) );
AND2x2_ASAP7_75t_L g345 ( .A(n_241), .B(n_277), .Y(n_345) );
AND2x2_ASAP7_75t_L g406 ( .A(n_241), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g276 ( .A(n_242), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g334 ( .A(n_242), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_247), .B(n_249), .Y(n_248) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_251), .Y(n_518) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
CKINVDCx16_ASAP7_75t_R g355 ( .A(n_254), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_255), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
AOI221x1_ASAP7_75t_SL g322 ( .A1(n_256), .A2(n_323), .B1(n_325), .B2(n_327), .C(n_329), .Y(n_322) );
INVx2_ASAP7_75t_L g270 ( .A(n_257), .Y(n_270) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_257), .Y(n_364) );
INVx2_ASAP7_75t_L g494 ( .A(n_264), .Y(n_494) );
INVx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g352 ( .A(n_267), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_271), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_268), .B(n_285), .Y(n_377) );
INVx1_ASAP7_75t_SL g440 ( .A(n_268), .Y(n_440) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g358 ( .A(n_271), .B(n_284), .Y(n_358) );
INVx1_ASAP7_75t_L g426 ( .A(n_272), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_272), .B(n_355), .Y(n_439) );
INVx2_ASAP7_75t_SL g278 ( .A(n_273), .Y(n_278) );
AND2x2_ASAP7_75t_L g321 ( .A(n_273), .B(n_277), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_273), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_273), .B(n_348), .Y(n_375) );
AOI21xp33_ASAP7_75t_SL g274 ( .A1(n_275), .A2(n_278), .B(n_279), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_276), .B(n_348), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_276), .B(n_303), .Y(n_444) );
OR2x2_ASAP7_75t_L g316 ( .A(n_277), .B(n_295), .Y(n_316) );
AND2x2_ASAP7_75t_L g415 ( .A(n_277), .B(n_406), .Y(n_415) );
OAI22xp5_ASAP7_75t_SL g290 ( .A1(n_278), .A2(n_291), .B1(n_296), .B2(n_299), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_278), .B(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g338 ( .A(n_280), .B(n_286), .Y(n_338) );
INVx1_ASAP7_75t_L g402 ( .A(n_280), .Y(n_402) );
AOI311xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_287), .A3(n_289), .B(n_290), .C(n_301), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_285), .A2(n_417), .B1(n_429), .B2(n_432), .C(n_434), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_285), .B(n_440), .Y(n_442) );
INVx2_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g339 ( .A(n_287), .Y(n_339) );
AOI211xp5_ASAP7_75t_L g329 ( .A1(n_288), .A2(n_330), .B(n_331), .C(n_333), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
O2A1O1Ixp33_ASAP7_75t_SL g398 ( .A1(n_292), .A2(n_294), .B(n_399), .C(n_400), .Y(n_398) );
INVx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_293), .B(n_367), .Y(n_433) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
OAI221xp5_ASAP7_75t_L g315 ( .A1(n_296), .A2(n_316), .B1(n_317), .B2(n_320), .C(n_322), .Y(n_315) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g318 ( .A(n_298), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g401 ( .A(n_298), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_305), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g359 ( .A1(n_302), .A2(n_360), .B(n_361), .C(n_365), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_303), .B(n_304), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_303), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_303), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g325 ( .A(n_309), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_313), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g427 ( .A(n_316), .Y(n_427) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_319), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g354 ( .A(n_319), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_SL g431 ( .A(n_319), .Y(n_431) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g372 ( .A(n_321), .B(n_348), .Y(n_372) );
INVx1_ASAP7_75t_SL g366 ( .A(n_328), .Y(n_366) );
INVx1_ASAP7_75t_L g343 ( .A(n_334), .Y(n_343) );
NAND3xp33_ASAP7_75t_SL g335 ( .A(n_336), .B(n_353), .C(n_369), .Y(n_335) );
AOI322xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_339), .A3(n_340), .B1(n_342), .B2(n_346), .C1(n_350), .C2(n_352), .Y(n_336) );
AOI211xp5_ASAP7_75t_L g389 ( .A1(n_337), .A2(n_390), .B(n_391), .C(n_398), .Y(n_389) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_340), .A2(n_361), .B1(n_392), .B2(n_394), .Y(n_391) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g350 ( .A(n_348), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g387 ( .A(n_348), .B(n_388), .Y(n_387) );
AOI32xp33_ASAP7_75t_L g438 ( .A1(n_348), .A2(n_439), .A3(n_440), .B1(n_441), .B2(n_443), .Y(n_438) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g360 ( .A(n_351), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_351), .A2(n_404), .B1(n_408), .B2(n_410), .C(n_413), .Y(n_403) );
AND2x2_ASAP7_75t_L g417 ( .A(n_351), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g420 ( .A(n_355), .B(n_421), .Y(n_420) );
OR2x2_ASAP7_75t_L g430 ( .A(n_355), .B(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVxp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g421 ( .A(n_364), .B(n_385), .Y(n_421) );
AOI211xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_372), .B(n_373), .C(n_376), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AOI21xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B(n_380), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI211xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_386), .B(n_389), .C(n_403), .Y(n_382) );
INVxp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_397), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g412 ( .A(n_409), .Y(n_412) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI21xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .B(n_419), .Y(n_413) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI211xp5_ASAP7_75t_SL g422 ( .A1(n_423), .A2(n_425), .B(n_428), .C(n_438), .Y(n_422) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_424), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI21xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B(n_437), .Y(n_434) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVxp67_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx2_ASAP7_75t_L g728 ( .A(n_450), .Y(n_728) );
BUFx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND3x1_ASAP7_75t_L g451 ( .A(n_452), .B(n_645), .C(n_690), .Y(n_451) );
NOR4xp25_ASAP7_75t_L g452 ( .A(n_453), .B(n_568), .C(n_609), .D(n_626), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_484), .B(n_498), .C(n_531), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_464), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_455), .B(n_485), .Y(n_484) );
NOR4xp25_ASAP7_75t_L g592 ( .A(n_455), .B(n_586), .C(n_593), .D(n_599), .Y(n_592) );
AND2x2_ASAP7_75t_L g665 ( .A(n_455), .B(n_554), .Y(n_665) );
AND2x2_ASAP7_75t_L g684 ( .A(n_455), .B(n_630), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_455), .B(n_679), .Y(n_693) );
AND2x2_ASAP7_75t_L g706 ( .A(n_455), .B(n_497), .Y(n_706) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_SL g551 ( .A(n_456), .Y(n_551) );
AND2x2_ASAP7_75t_L g558 ( .A(n_456), .B(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g608 ( .A(n_456), .B(n_465), .Y(n_608) );
AND2x2_ASAP7_75t_SL g619 ( .A(n_456), .B(n_554), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_456), .B(n_465), .Y(n_623) );
AND2x2_ASAP7_75t_L g632 ( .A(n_456), .B(n_557), .Y(n_632) );
BUFx2_ASAP7_75t_L g655 ( .A(n_456), .Y(n_655) );
AND2x2_ASAP7_75t_L g659 ( .A(n_456), .B(n_475), .Y(n_659) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_475), .Y(n_464) );
AND2x2_ASAP7_75t_L g497 ( .A(n_465), .B(n_475), .Y(n_497) );
BUFx2_ASAP7_75t_L g561 ( .A(n_465), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_465), .A2(n_594), .B1(n_596), .B2(n_597), .Y(n_593) );
OR2x2_ASAP7_75t_L g615 ( .A(n_465), .B(n_487), .Y(n_615) );
AND2x2_ASAP7_75t_L g679 ( .A(n_465), .B(n_557), .Y(n_679) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g547 ( .A(n_466), .B(n_487), .Y(n_547) );
AND2x2_ASAP7_75t_L g554 ( .A(n_466), .B(n_475), .Y(n_554) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_466), .Y(n_596) );
OR2x2_ASAP7_75t_L g631 ( .A(n_466), .B(n_486), .Y(n_631) );
INVx1_ASAP7_75t_L g550 ( .A(n_475), .Y(n_550) );
INVx3_ASAP7_75t_L g559 ( .A(n_475), .Y(n_559) );
BUFx2_ASAP7_75t_L g583 ( .A(n_475), .Y(n_583) );
AND2x2_ASAP7_75t_L g616 ( .A(n_475), .B(n_551), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_484), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_701) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_497), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_486), .B(n_559), .Y(n_563) );
INVx1_ASAP7_75t_L g591 ( .A(n_486), .Y(n_591) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_L g557 ( .A(n_487), .Y(n_557) );
INVx1_ASAP7_75t_L g569 ( .A(n_497), .Y(n_569) );
NAND2x1_ASAP7_75t_SL g498 ( .A(n_499), .B(n_509), .Y(n_498) );
AND2x2_ASAP7_75t_L g567 ( .A(n_499), .B(n_522), .Y(n_567) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_499), .Y(n_641) );
AND2x2_ASAP7_75t_L g668 ( .A(n_499), .B(n_588), .Y(n_668) );
AND2x2_ASAP7_75t_L g676 ( .A(n_499), .B(n_638), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_499), .B(n_534), .Y(n_703) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g535 ( .A(n_500), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g552 ( .A(n_500), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g573 ( .A(n_500), .Y(n_573) );
INVx1_ASAP7_75t_L g579 ( .A(n_500), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_500), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g612 ( .A(n_500), .B(n_537), .Y(n_612) );
OR2x2_ASAP7_75t_L g650 ( .A(n_500), .B(n_605), .Y(n_650) );
AOI32xp33_ASAP7_75t_L g662 ( .A1(n_500), .A2(n_663), .A3(n_666), .B1(n_667), .B2(n_668), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_500), .B(n_638), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_500), .B(n_598), .Y(n_713) );
OR2x6_ASAP7_75t_L g500 ( .A(n_501), .B(n_507), .Y(n_500) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_L g624 ( .A(n_510), .B(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_522), .Y(n_510) );
INVx1_ASAP7_75t_L g586 ( .A(n_511), .Y(n_586) );
AND2x2_ASAP7_75t_L g588 ( .A(n_511), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_511), .B(n_536), .Y(n_605) );
AND2x2_ASAP7_75t_L g638 ( .A(n_511), .B(n_614), .Y(n_638) );
AND2x2_ASAP7_75t_L g675 ( .A(n_511), .B(n_537), .Y(n_675) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g534 ( .A(n_512), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_512), .B(n_536), .Y(n_565) );
AND2x2_ASAP7_75t_L g572 ( .A(n_512), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g613 ( .A(n_512), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_519), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B(n_518), .Y(n_515) );
INVx2_ASAP7_75t_L g589 ( .A(n_522), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_522), .B(n_536), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_522), .B(n_580), .Y(n_661) );
INVx1_ASAP7_75t_L g683 ( .A(n_522), .Y(n_683) );
INVx1_ASAP7_75t_L g700 ( .A(n_522), .Y(n_700) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g553 ( .A(n_523), .B(n_536), .Y(n_553) );
AND2x2_ASAP7_75t_L g575 ( .A(n_523), .B(n_537), .Y(n_575) );
INVx1_ASAP7_75t_L g614 ( .A(n_523), .Y(n_614) );
AOI221x1_ASAP7_75t_SL g531 ( .A1(n_532), .A2(n_546), .B1(n_552), .B2(n_554), .C(n_555), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_532), .A2(n_619), .B1(n_686), .B2(n_687), .Y(n_685) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
AND2x2_ASAP7_75t_L g577 ( .A(n_533), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g672 ( .A(n_533), .B(n_552), .Y(n_672) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g628 ( .A(n_534), .B(n_553), .Y(n_628) );
INVx1_ASAP7_75t_L g640 ( .A(n_535), .Y(n_640) );
AND2x2_ASAP7_75t_L g651 ( .A(n_535), .B(n_638), .Y(n_651) );
AND2x2_ASAP7_75t_L g718 ( .A(n_535), .B(n_613), .Y(n_718) );
INVx2_ASAP7_75t_L g580 ( .A(n_536), .Y(n_580) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_547), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g670 ( .A(n_547), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_548), .B(n_631), .Y(n_634) );
INVx3_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_549), .A2(n_670), .B(n_715), .Y(n_714) );
AND2x4_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NOR2xp33_ASAP7_75t_SL g692 ( .A(n_552), .B(n_578), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_553), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g644 ( .A(n_553), .B(n_572), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_553), .B(n_579), .Y(n_721) );
AND2x2_ASAP7_75t_L g590 ( .A(n_554), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g657 ( .A(n_554), .Y(n_657) );
AOI21xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_560), .B(n_564), .Y(n_555) );
NAND2x1_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_557), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g606 ( .A(n_557), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g618 ( .A(n_557), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_557), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g642 ( .A(n_558), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_558), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_558), .B(n_561), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
AOI211xp5_ASAP7_75t_L g629 ( .A1(n_561), .A2(n_600), .B(n_630), .C(n_632), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_561), .A2(n_648), .B1(n_651), .B2(n_652), .C(n_656), .Y(n_647) );
AND2x2_ASAP7_75t_L g643 ( .A(n_562), .B(n_596), .Y(n_643) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g603 ( .A(n_567), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g674 ( .A(n_567), .B(n_675), .Y(n_674) );
OAI211xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B(n_576), .C(n_601), .Y(n_568) );
NAND3xp33_ASAP7_75t_SL g687 ( .A(n_569), .B(n_688), .C(n_689), .Y(n_687) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_574), .Y(n_570) );
OR2x2_ASAP7_75t_L g660 ( .A(n_571), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_581), .B1(n_584), .B2(n_590), .C(n_592), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_578), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_578), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g600 ( .A(n_583), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_583), .A2(n_640), .B1(n_641), .B2(n_642), .Y(n_639) );
OR2x2_ASAP7_75t_L g720 ( .A(n_583), .B(n_631), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_585), .B(n_587), .Y(n_584) );
INVxp67_ASAP7_75t_L g694 ( .A(n_586), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_588), .B(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_L g595 ( .A(n_589), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_591), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_591), .B(n_638), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_591), .B(n_658), .Y(n_697) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_595), .Y(n_621) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g711 ( .A(n_600), .B(n_631), .Y(n_711) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_606), .Y(n_602) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_SL g689 ( .A(n_606), .Y(n_689) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OAI322xp33_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_615), .A3(n_616), .B1(n_617), .B2(n_620), .C1(n_622), .C2(n_624), .Y(n_609) );
OAI322xp33_ASAP7_75t_L g691 ( .A1(n_610), .A2(n_692), .A3(n_693), .B1(n_694), .B2(n_695), .C1(n_696), .C2(n_698), .Y(n_691) );
CKINVDCx16_ASAP7_75t_R g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx4_ASAP7_75t_L g625 ( .A(n_612), .Y(n_625) );
AND2x2_ASAP7_75t_L g686 ( .A(n_612), .B(n_638), .Y(n_686) );
AND2x2_ASAP7_75t_L g699 ( .A(n_612), .B(n_700), .Y(n_699) );
CKINVDCx16_ASAP7_75t_R g710 ( .A(n_615), .Y(n_710) );
INVx1_ASAP7_75t_L g688 ( .A(n_616), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
OR2x2_ASAP7_75t_L g622 ( .A(n_618), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g705 ( .A(n_618), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_618), .B(n_659), .Y(n_716) );
OR2x2_ASAP7_75t_L g649 ( .A(n_621), .B(n_650), .Y(n_649) );
INVxp33_ASAP7_75t_L g666 ( .A(n_621), .Y(n_666) );
OAI221xp5_ASAP7_75t_SL g626 ( .A1(n_625), .A2(n_627), .B1(n_629), .B2(n_633), .C(n_635), .Y(n_626) );
NOR2xp67_ASAP7_75t_L g682 ( .A(n_625), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g709 ( .A(n_625), .Y(n_709) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
INVx3_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
AOI322xp5_ASAP7_75t_L g673 ( .A1(n_632), .A2(n_657), .A3(n_674), .B1(n_676), .B2(n_677), .C1(n_680), .C2(n_684), .Y(n_673) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_639), .B1(n_643), .B2(n_644), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_646), .B(n_669), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_647), .B(n_662), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_650), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
NAND2xp33_ASAP7_75t_SL g667 ( .A(n_653), .B(n_664), .Y(n_667) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
OAI322xp33_ASAP7_75t_L g707 ( .A1(n_655), .A2(n_708), .A3(n_710), .B1(n_711), .B2(n_712), .C1(n_714), .C2(n_717), .Y(n_707) );
AOI21xp33_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_658), .B(n_660), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_665), .B(n_713), .Y(n_722) );
OAI211xp5_ASAP7_75t_SL g669 ( .A1(n_670), .A2(n_671), .B(n_673), .C(n_685), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NOR4xp25_ASAP7_75t_L g690 ( .A(n_691), .B(n_701), .C(n_707), .D(n_719), .Y(n_690) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
INVxp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
CKINVDCx14_ASAP7_75t_R g717 ( .A(n_718), .Y(n_717) );
OAI21xp5_ASAP7_75t_SL g719 ( .A1(n_720), .A2(n_721), .B(n_722), .Y(n_719) );
INVx1_ASAP7_75t_L g729 ( .A(n_723), .Y(n_729) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_737), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OAI21xp5_ASAP7_75t_SL g738 ( .A1(n_739), .A2(n_743), .B(n_745), .Y(n_738) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
BUFx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_750), .Y(n_749) );
endmodule