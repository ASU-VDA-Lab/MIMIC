module fake_jpeg_29251_n_295 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_295);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx6_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_1),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx12_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_67),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_69),
.Y(n_87)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_70),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_72),
.Y(n_83)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_43),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_39),
.B1(n_23),
.B2(n_24),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_75),
.A2(n_27),
.B1(n_31),
.B2(n_28),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_36),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_21),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_24),
.B1(n_21),
.B2(n_25),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_81),
.B1(n_68),
.B2(n_40),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_23),
.B1(n_25),
.B2(n_27),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_102),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_73),
.B1(n_69),
.B2(n_51),
.Y(n_81)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_26),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_105),
.B(n_115),
.Y(n_149)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_107),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_82),
.B(n_26),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_113),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_136),
.B1(n_98),
.B2(n_91),
.Y(n_138)
);

BUFx2_ASAP7_75t_SL g110 ( 
.A(n_78),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

HAxp5_ASAP7_75t_SL g111 ( 
.A(n_80),
.B(n_37),
.CON(n_111),
.SN(n_111)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_119),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_83),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_35),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_116),
.B(n_122),
.Y(n_158)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_118),
.A2(n_131),
.B1(n_86),
.B2(n_103),
.Y(n_150)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_121),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_155)
);

AO22x1_ASAP7_75t_SL g122 ( 
.A1(n_88),
.A2(n_45),
.B1(n_49),
.B2(n_40),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_88),
.A2(n_30),
.B1(n_38),
.B2(n_28),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_38),
.Y(n_124)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_124),
.B(n_127),
.CI(n_132),
.CON(n_153),
.SN(n_153)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_78),
.A2(n_30),
.B1(n_31),
.B2(n_44),
.Y(n_126)
);

INVx6_ASAP7_75t_SL g127 ( 
.A(n_86),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_129),
.B(n_130),
.Y(n_146)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_101),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_84),
.A2(n_36),
.B1(n_35),
.B2(n_43),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_92),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_134),
.B(n_135),
.Y(n_145)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_117),
.B1(n_133),
.B2(n_106),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_91),
.B1(n_85),
.B2(n_93),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_142),
.B1(n_130),
.B2(n_131),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_85),
.B1(n_90),
.B2(n_95),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_154),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_123),
.B1(n_111),
.B2(n_122),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_122),
.A2(n_92),
.B1(n_103),
.B2(n_43),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_126),
.A2(n_43),
.B1(n_3),
.B2(n_5),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_159),
.A2(n_163),
.B1(n_154),
.B2(n_137),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_146),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_164),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_155),
.A2(n_121),
.B1(n_134),
.B2(n_114),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_146),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_165),
.Y(n_192)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_168),
.B(n_171),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_124),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_170),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_104),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVxp33_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_172),
.Y(n_180)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_173),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_170),
.C(n_153),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_189),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_167),
.A2(n_158),
.B1(n_138),
.B2(n_139),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_185),
.B1(n_193),
.B2(n_196),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_167),
.A2(n_158),
.B1(n_160),
.B2(n_164),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_151),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_176),
.B(n_157),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_149),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_175),
.A2(n_139),
.B1(n_141),
.B2(n_152),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_162),
.A2(n_139),
.B(n_150),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_142),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_186),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_187),
.A2(n_137),
.B(n_171),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_210),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_187),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_204),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_178),
.A2(n_166),
.B1(n_165),
.B2(n_168),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_213),
.B1(n_180),
.B2(n_179),
.Y(n_222)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_208),
.B(n_195),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_192),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_209),
.Y(n_214)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_191),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_212),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_148),
.B(n_149),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_208),
.B(n_188),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_148),
.C(n_194),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_198),
.A2(n_196),
.B1(n_189),
.B2(n_180),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_219),
.A2(n_222),
.B1(n_201),
.B2(n_206),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_183),
.B1(n_185),
.B2(n_193),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_223),
.A2(n_203),
.B1(n_211),
.B2(n_194),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_228),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_225),
.A2(n_198),
.B(n_202),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_229),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_227),
.A2(n_213),
.B1(n_212),
.B2(n_205),
.Y(n_230)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_231),
.A2(n_223),
.B1(n_225),
.B2(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_233),
.A2(n_144),
.B1(n_5),
.B2(n_7),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_203),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_236),
.Y(n_249)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_238),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_184),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_144),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_191),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_241),
.Y(n_253)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_140),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_214),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_215),
.C(n_221),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_247),
.C(n_254),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_245),
.A2(n_231),
.B1(n_236),
.B2(n_237),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_217),
.C(n_220),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_255),
.B1(n_251),
.B2(n_253),
.Y(n_258)
);

INVxp33_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_250),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_2),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_250),
.A2(n_239),
.B(n_237),
.Y(n_257)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_264),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_252),
.A2(n_16),
.B(n_15),
.Y(n_260)
);

AOI21x1_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_2),
.B(n_7),
.Y(n_275)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_263),
.Y(n_274)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_14),
.C(n_5),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_244),
.C(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_266),
.B(n_12),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_267),
.B(n_271),
.Y(n_279)
);

OAI21x1_ASAP7_75t_SL g268 ( 
.A1(n_261),
.A2(n_249),
.B(n_14),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_268),
.A2(n_272),
.B1(n_274),
.B2(n_270),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_260),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_265),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_275),
.A2(n_259),
.B(n_257),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_278),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_277),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_262),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_280),
.B(n_281),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_256),
.B1(n_262),
.B2(n_9),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_279),
.B(n_267),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_283),
.A2(n_278),
.B(n_276),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_287),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_285),
.A2(n_275),
.B(n_8),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_284),
.Y(n_288)
);

O2A1O1Ixp33_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_282),
.B(n_8),
.C(n_9),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_289),
.A2(n_7),
.B(n_8),
.Y(n_291)
);

AO21x1_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_290),
.B(n_11),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_10),
.C(n_12),
.Y(n_293)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_293),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_10),
.B1(n_12),
.B2(n_282),
.Y(n_295)
);


endmodule