module fake_jpeg_30632_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_41),
.Y(n_52)
);

CKINVDCx11_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_44),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_17),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_35),
.B1(n_22),
.B2(n_17),
.Y(n_59)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

HAxp5_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_32),
.CON(n_51),
.SN(n_51)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_51),
.A2(n_26),
.B(n_38),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_76),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_28),
.B1(n_36),
.B2(n_23),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_74),
.B1(n_75),
.B2(n_22),
.Y(n_78)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_64),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_32),
.B1(n_34),
.B2(n_30),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_42),
.B1(n_48),
.B2(n_24),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_77),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_42),
.A2(n_33),
.B1(n_23),
.B2(n_20),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_23),
.B1(n_36),
.B2(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_38),
.B(n_30),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_78),
.A2(n_25),
.B1(n_21),
.B2(n_4),
.Y(n_150)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_77),
.B(n_24),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_82),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_43),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_83),
.B(n_87),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_36),
.B1(n_20),
.B2(n_19),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_109),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_37),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_90),
.A2(n_101),
.B(n_26),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_51),
.B(n_37),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_96),
.B(n_99),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_18),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_39),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_68),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_102),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_18),
.Y(n_103)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_44),
.Y(n_104)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_26),
.B(n_48),
.C(n_25),
.Y(n_141)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_41),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_66),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_113),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_SL g112 ( 
.A(n_66),
.B(n_31),
.C(n_43),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_117),
.B1(n_118),
.B2(n_17),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_41),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_73),
.B(n_19),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_58),
.A2(n_20),
.B1(n_33),
.B2(n_26),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_33),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_119),
.B(n_121),
.C(n_125),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_49),
.C(n_46),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_91),
.A2(n_70),
.B1(n_48),
.B2(n_42),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_124),
.A2(n_140),
.B1(n_144),
.B2(n_111),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_49),
.C(n_46),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_129),
.B(n_141),
.Y(n_180)
);

AOI32xp33_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_49),
.A3(n_46),
.B1(n_35),
.B2(n_22),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_90),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_46),
.C(n_49),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_152),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_96),
.A2(n_35),
.B(n_15),
.C(n_11),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_139),
.B(n_149),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_85),
.A2(n_48),
.B1(n_69),
.B2(n_65),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_101),
.A2(n_70),
.B1(n_58),
.B2(n_26),
.Y(n_144)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_150),
.A2(n_101),
.B1(n_90),
.B2(n_93),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_80),
.C(n_85),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_153),
.A2(n_94),
.B1(n_115),
.B2(n_134),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_155),
.A2(n_158),
.B(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_85),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_166),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_97),
.B(n_92),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_122),
.B(n_89),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_165),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_92),
.B(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_95),
.B(n_98),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_163),
.A2(n_182),
.B(n_123),
.Y(n_197)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_78),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_126),
.B(n_81),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_168),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_148),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_81),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_173),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_171),
.A2(n_150),
.B1(n_147),
.B2(n_142),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_130),
.A2(n_78),
.B1(n_95),
.B2(n_98),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_172),
.A2(n_26),
.B1(n_25),
.B2(n_21),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_119),
.B(n_78),
.Y(n_173)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_130),
.A2(n_81),
.B1(n_94),
.B2(n_88),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_132),
.B(n_100),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_152),
.Y(n_194)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g186 ( 
.A(n_157),
.B(n_148),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_202),
.B1(n_205),
.B2(n_207),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_211),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_161),
.A2(n_139),
.B(n_149),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_195),
.A2(n_212),
.B(n_169),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_180),
.A2(n_153),
.B1(n_154),
.B2(n_168),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_196),
.A2(n_197),
.B(n_175),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_125),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_201),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_137),
.C(n_121),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_166),
.A2(n_144),
.B1(n_141),
.B2(n_116),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_173),
.B(n_100),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_209),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_171),
.A2(n_79),
.B1(n_88),
.B2(n_114),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_180),
.A2(n_115),
.B1(n_94),
.B2(n_114),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_174),
.B(n_138),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_107),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_154),
.A2(n_108),
.B(n_134),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_214),
.A2(n_216),
.B1(n_156),
.B2(n_165),
.Y(n_234)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_217),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_211),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_219),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_180),
.B1(n_158),
.B2(n_163),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_224),
.A2(n_227),
.B1(n_214),
.B2(n_189),
.Y(n_252)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_205),
.A2(n_184),
.B1(n_174),
.B2(n_160),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_197),
.A2(n_160),
.B1(n_176),
.B2(n_179),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_239),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_178),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_201),
.C(n_209),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_199),
.Y(n_233)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_243),
.B1(n_186),
.B2(n_188),
.Y(n_257)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_192),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_236),
.Y(n_254)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_237),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_193),
.B(n_177),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_245),
.Y(n_247)
);

INVxp67_ASAP7_75t_R g239 ( 
.A(n_195),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_240),
.A2(n_212),
.B(n_190),
.Y(n_250)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_244),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_196),
.A2(n_105),
.B1(n_9),
.B2(n_12),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_187),
.Y(n_244)
);

NAND3xp33_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_7),
.C(n_16),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_220),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_250),
.A2(n_256),
.B(n_259),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_252),
.A2(n_15),
.B1(n_13),
.B2(n_9),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_224),
.A2(n_185),
.B1(n_189),
.B2(n_186),
.Y(n_255)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_257),
.A2(n_259),
.B1(n_261),
.B2(n_263),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_222),
.A2(n_185),
.B1(n_190),
.B2(n_203),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_221),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_188),
.B1(n_217),
.B2(n_208),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_243),
.A2(n_239),
.B1(n_234),
.B2(n_241),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_210),
.B1(n_206),
.B2(n_200),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_222),
.A2(n_225),
.B1(n_227),
.B2(n_231),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_264),
.A2(n_192),
.B1(n_105),
.B2(n_4),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_220),
.B(n_200),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_221),
.C(n_223),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_274),
.Y(n_298)
);

AND2x2_ASAP7_75t_SL g270 ( 
.A(n_249),
.B(n_230),
.Y(n_270)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_270),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_232),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_277),
.C(n_283),
.Y(n_292)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_266),
.Y(n_273)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_252),
.Y(n_299)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_278),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_218),
.C(n_236),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_282),
.Y(n_291)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_246),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_281),
.B(n_285),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_1),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_105),
.C(n_9),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_284),
.A2(n_250),
.B(n_256),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_16),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_287),
.B1(n_15),
.B2(n_13),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_247),
.B(n_255),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_265),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_265),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_293),
.A2(n_295),
.B(n_270),
.Y(n_314)
);

AO221x1_ASAP7_75t_L g295 ( 
.A1(n_280),
.A2(n_260),
.B1(n_251),
.B2(n_262),
.C(n_247),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_284),
.A2(n_256),
.B1(n_254),
.B2(n_261),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_300),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_272),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_263),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_264),
.C(n_257),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_299),
.C(n_292),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_303),
.A2(n_279),
.B1(n_272),
.B2(n_286),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_294),
.B(n_270),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_297),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_310),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_269),
.C(n_274),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_309),
.B(n_311),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_302),
.A2(n_275),
.B(n_283),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_313),
.A2(n_291),
.B1(n_300),
.B2(n_298),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_293),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_304),
.A2(n_271),
.B1(n_3),
.B2(n_4),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_304),
.B1(n_290),
.B2(n_4),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_308),
.B(n_301),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_318),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_309),
.B(n_289),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_320),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_324),
.B1(n_312),
.B2(n_313),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_323),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_305),
.A2(n_291),
.B1(n_298),
.B2(n_5),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_316),
.A2(n_312),
.B(n_307),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_328),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_324),
.A2(n_315),
.B1(n_310),
.B2(n_5),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_329),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_321),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_331),
.B(n_334),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_321),
.C(n_3),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_325),
.C(n_327),
.Y(n_335)
);

OAI211xp5_ASAP7_75t_L g337 ( 
.A1(n_335),
.A2(n_330),
.B(n_333),
.C(n_5),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_337),
.Y(n_338)
);

AO21x2_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_336),
.B(n_3),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_1),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_6),
.B(n_339),
.Y(n_341)
);


endmodule