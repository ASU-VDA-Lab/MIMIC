module fake_ariane_3028_n_96 (n_8, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_10, n_96);

input n_8;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_10;

output n_96;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_74;
wire n_33;
wire n_40;
wire n_53;
wire n_66;
wire n_71;
wire n_24;
wire n_49;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_44;
wire n_30;
wire n_82;
wire n_42;
wire n_31;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_88;
wire n_68;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_35;
wire n_54;
wire n_25;

INVx4_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_5),
.B(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2x1_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

OA21x2_ASAP7_75t_L g29 ( 
.A1(n_14),
.A2(n_9),
.B(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

OAI21x1_ASAP7_75t_L g31 ( 
.A1(n_18),
.A2(n_19),
.B(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

AND2x4_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_13),
.Y(n_34)
);

CKINVDCx11_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

AND2x6_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_3),
.A2(n_7),
.B1(n_10),
.B2(n_6),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_8),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_25),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_34),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_24),
.B(n_34),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_24),
.B(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

AOI21x1_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_53),
.B(n_49),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_50),
.B(n_45),
.Y(n_62)
);

OAI21x1_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_29),
.B(n_41),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_35),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

OR2x2_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_33),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_38),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_62),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_74),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_74),
.Y(n_78)
);

AOI211xp5_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_67),
.B(n_71),
.C(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_75),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_63),
.B(n_67),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_27),
.C(n_72),
.Y(n_82)
);

NOR4xp25_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_58),
.C(n_65),
.D(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

NAND4xp25_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_72),
.C(n_65),
.D(n_32),
.Y(n_85)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_73),
.B(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

OAI22x1_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_78),
.B1(n_82),
.B2(n_29),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_63),
.C(n_60),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_76),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_32),
.B1(n_26),
.B2(n_39),
.Y(n_93)
);

NOR4xp25_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_36),
.C(n_65),
.D(n_90),
.Y(n_94)
);

OAI21x1_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_91),
.B(n_93),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_36),
.Y(n_96)
);


endmodule