module real_aes_7505_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_0), .B(n_109), .C(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g457 ( .A(n_0), .Y(n_457) );
INVx1_ASAP7_75t_L g490 ( .A(n_1), .Y(n_490) );
INVx1_ASAP7_75t_L g199 ( .A(n_2), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_3), .A2(n_37), .B1(n_160), .B2(n_520), .Y(n_535) );
AOI21xp33_ASAP7_75t_L g167 ( .A1(n_4), .A2(n_141), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_5), .B(n_134), .Y(n_503) );
AND2x6_ASAP7_75t_L g146 ( .A(n_6), .B(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_7), .A2(n_249), .B(n_250), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_8), .B(n_38), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_8), .B(n_38), .Y(n_458) );
INVx1_ASAP7_75t_L g174 ( .A(n_9), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_10), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g139 ( .A(n_11), .Y(n_139) );
INVx1_ASAP7_75t_L g484 ( .A(n_12), .Y(n_484) );
INVx1_ASAP7_75t_L g255 ( .A(n_13), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_14), .B(n_182), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_15), .B(n_135), .Y(n_561) );
AO32x2_ASAP7_75t_L g533 ( .A1(n_16), .A2(n_134), .A3(n_179), .B1(n_512), .B2(n_534), .Y(n_533) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_17), .A2(n_62), .B1(n_123), .B2(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g124 ( .A(n_17), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_18), .B(n_160), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_19), .B(n_155), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_20), .B(n_135), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_21), .A2(n_50), .B1(n_160), .B2(n_520), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_22), .B(n_141), .Y(n_211) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_23), .A2(n_78), .B1(n_160), .B2(n_182), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_24), .B(n_160), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_25), .B(n_163), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_26), .A2(n_253), .B(n_254), .C(n_256), .Y(n_252) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_27), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_28), .B(n_176), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_29), .B(n_172), .Y(n_201) );
INVx1_ASAP7_75t_L g188 ( .A(n_30), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g118 ( .A1(n_31), .A2(n_119), .B1(n_120), .B2(n_451), .Y(n_118) );
INVx1_ASAP7_75t_L g451 ( .A(n_31), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_32), .B(n_176), .Y(n_550) );
INVx2_ASAP7_75t_L g144 ( .A(n_33), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_34), .B(n_160), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_35), .B(n_176), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_36), .A2(n_146), .B(n_150), .C(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g186 ( .A(n_39), .Y(n_186) );
OAI22xp5_ASAP7_75t_SL g764 ( .A1(n_40), .A2(n_765), .B1(n_768), .B2(n_769), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_40), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_41), .B(n_172), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_42), .B(n_160), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_43), .A2(n_89), .B1(n_218), .B2(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_44), .B(n_160), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_45), .B(n_160), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g189 ( .A(n_46), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_47), .A2(n_71), .B1(n_766), .B2(n_767), .Y(n_765) );
CKINVDCx16_ASAP7_75t_R g767 ( .A(n_47), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_48), .B(n_489), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_49), .B(n_141), .Y(n_243) );
AOI22xp33_ASAP7_75t_SL g559 ( .A1(n_51), .A2(n_60), .B1(n_160), .B2(n_182), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_52), .A2(n_150), .B1(n_182), .B2(n_184), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_53), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_54), .B(n_160), .Y(n_511) );
CKINVDCx16_ASAP7_75t_R g196 ( .A(n_55), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_56), .B(n_160), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_57), .A2(n_159), .B(n_171), .C(n_173), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_58), .Y(n_231) );
INVx1_ASAP7_75t_L g169 ( .A(n_59), .Y(n_169) );
INVx1_ASAP7_75t_L g147 ( .A(n_61), .Y(n_147) );
INVx1_ASAP7_75t_L g123 ( .A(n_62), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_63), .A2(n_104), .B1(n_113), .B2(n_777), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_64), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_65), .B(n_160), .Y(n_491) );
INVx1_ASAP7_75t_L g138 ( .A(n_66), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_67), .Y(n_116) );
AO32x2_ASAP7_75t_L g517 ( .A1(n_68), .A2(n_134), .A3(n_235), .B1(n_512), .B2(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g510 ( .A(n_69), .Y(n_510) );
INVx1_ASAP7_75t_L g545 ( .A(n_70), .Y(n_545) );
INVx1_ASAP7_75t_L g766 ( .A(n_71), .Y(n_766) );
A2O1A1Ixp33_ASAP7_75t_SL g154 ( .A1(n_72), .A2(n_155), .B(n_156), .C(n_159), .Y(n_154) );
INVxp67_ASAP7_75t_L g157 ( .A(n_73), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_74), .B(n_182), .Y(n_546) );
INVx1_ASAP7_75t_L g112 ( .A(n_75), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_76), .Y(n_192) );
INVx1_ASAP7_75t_L g224 ( .A(n_77), .Y(n_224) );
AOI222xp33_ASAP7_75t_L g462 ( .A1(n_79), .A2(n_463), .B1(n_763), .B2(n_764), .C1(n_770), .C2(n_771), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_80), .A2(n_146), .B(n_150), .C(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_81), .B(n_520), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_82), .B(n_182), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_83), .B(n_200), .Y(n_214) );
INVx2_ASAP7_75t_L g136 ( .A(n_84), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_85), .B(n_155), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_86), .B(n_182), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_87), .A2(n_146), .B(n_150), .C(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g109 ( .A(n_88), .Y(n_109) );
OR2x2_ASAP7_75t_L g454 ( .A(n_88), .B(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g468 ( .A(n_88), .B(n_456), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_90), .A2(n_102), .B1(n_182), .B2(n_183), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_91), .B(n_176), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_92), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_93), .A2(n_146), .B(n_150), .C(n_238), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_94), .Y(n_245) );
INVx1_ASAP7_75t_L g153 ( .A(n_95), .Y(n_153) );
CKINVDCx16_ASAP7_75t_R g251 ( .A(n_96), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_97), .B(n_200), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_98), .B(n_182), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_99), .B(n_134), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_100), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_101), .A2(n_141), .B(n_148), .Y(n_140) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g778 ( .A(n_105), .Y(n_778) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
OR2x2_ASAP7_75t_L g470 ( .A(n_109), .B(n_456), .Y(n_470) );
NOR2x2_ASAP7_75t_L g770 ( .A(n_109), .B(n_455), .Y(n_770) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AO21x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_117), .B(n_461), .Y(n_113) );
INVx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g776 ( .A(n_115), .Y(n_776) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OAI21xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_452), .B(n_459), .Y(n_117) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_122), .B1(n_125), .B2(n_450), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g450 ( .A(n_125), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_125), .A2(n_465), .B1(n_469), .B2(n_471), .Y(n_464) );
INVx1_ASAP7_75t_SL g773 ( .A(n_125), .Y(n_773) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND4x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_368), .C(n_415), .D(n_435), .Y(n_126) );
NOR3xp33_ASAP7_75t_SL g127 ( .A(n_128), .B(n_298), .C(n_323), .Y(n_127) );
OAI211xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_206), .B(n_258), .C(n_288), .Y(n_128) );
INVxp67_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_177), .Y(n_130) );
INVx3_ASAP7_75t_SL g340 ( .A(n_131), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_131), .B(n_271), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_131), .B(n_193), .Y(n_421) );
AND2x2_ASAP7_75t_L g444 ( .A(n_131), .B(n_310), .Y(n_444) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_165), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g262 ( .A(n_133), .B(n_166), .Y(n_262) );
INVx3_ASAP7_75t_L g275 ( .A(n_133), .Y(n_275) );
AND2x2_ASAP7_75t_L g280 ( .A(n_133), .B(n_165), .Y(n_280) );
OR2x2_ASAP7_75t_L g331 ( .A(n_133), .B(n_272), .Y(n_331) );
BUFx2_ASAP7_75t_L g351 ( .A(n_133), .Y(n_351) );
AND2x2_ASAP7_75t_L g361 ( .A(n_133), .B(n_272), .Y(n_361) );
AND2x2_ASAP7_75t_L g367 ( .A(n_133), .B(n_178), .Y(n_367) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_140), .B(n_162), .Y(n_133) );
INVx4_ASAP7_75t_L g164 ( .A(n_134), .Y(n_164) );
OA21x2_ASAP7_75t_L g495 ( .A1(n_134), .A2(n_496), .B(n_503), .Y(n_495) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g179 ( .A(n_135), .Y(n_179) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g176 ( .A(n_136), .B(n_137), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
BUFx2_ASAP7_75t_L g249 ( .A(n_141), .Y(n_249) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_146), .Y(n_141) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_142), .B(n_146), .Y(n_190) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
INVx1_ASAP7_75t_L g489 ( .A(n_143), .Y(n_489) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g151 ( .A(n_144), .Y(n_151) );
INVx1_ASAP7_75t_L g183 ( .A(n_144), .Y(n_183) );
INVx1_ASAP7_75t_L g152 ( .A(n_145), .Y(n_152) );
INVx1_ASAP7_75t_L g155 ( .A(n_145), .Y(n_155) );
INVx3_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_145), .Y(n_185) );
INVx4_ASAP7_75t_SL g161 ( .A(n_146), .Y(n_161) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_146), .A2(n_483), .B(n_487), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_146), .A2(n_497), .B(n_500), .Y(n_496) );
BUFx3_ASAP7_75t_L g512 ( .A(n_146), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_146), .A2(n_525), .B(n_529), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_146), .A2(n_544), .B(n_547), .Y(n_543) );
O2A1O1Ixp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_153), .B(n_154), .C(n_161), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g168 ( .A1(n_149), .A2(n_161), .B(n_169), .C(n_170), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_149), .A2(n_161), .B(n_251), .C(n_252), .Y(n_250) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x6_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_151), .Y(n_160) );
BUFx3_ASAP7_75t_L g218 ( .A(n_151), .Y(n_218) );
INVx1_ASAP7_75t_L g520 ( .A(n_151), .Y(n_520) );
INVx1_ASAP7_75t_L g528 ( .A(n_155), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_158), .B(n_174), .Y(n_173) );
INVx5_ASAP7_75t_L g200 ( .A(n_158), .Y(n_200) );
OAI22xp5_ASAP7_75t_SL g518 ( .A1(n_158), .A2(n_172), .B1(n_519), .B2(n_521), .Y(n_518) );
O2A1O1Ixp5_ASAP7_75t_SL g544 ( .A1(n_159), .A2(n_200), .B(n_545), .C(n_546), .Y(n_544) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_160), .Y(n_242) );
OAI22xp33_ASAP7_75t_L g180 ( .A1(n_161), .A2(n_181), .B1(n_189), .B2(n_190), .Y(n_180) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_163), .A2(n_167), .B(n_175), .Y(n_166) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_SL g220 ( .A(n_164), .B(n_221), .Y(n_220) );
AO21x1_ASAP7_75t_L g556 ( .A1(n_164), .A2(n_557), .B(n_560), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g575 ( .A(n_164), .B(n_512), .C(n_557), .Y(n_575) );
INVx1_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_166), .B(n_272), .Y(n_286) );
INVx2_ASAP7_75t_L g296 ( .A(n_166), .Y(n_296) );
AND2x2_ASAP7_75t_L g309 ( .A(n_166), .B(n_275), .Y(n_309) );
OR2x2_ASAP7_75t_L g320 ( .A(n_166), .B(n_272), .Y(n_320) );
AND2x2_ASAP7_75t_SL g366 ( .A(n_166), .B(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_L g378 ( .A(n_166), .Y(n_378) );
AND2x2_ASAP7_75t_L g424 ( .A(n_166), .B(n_178), .Y(n_424) );
O2A1O1Ixp5_ASAP7_75t_L g509 ( .A1(n_171), .A2(n_488), .B(n_510), .C(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_171), .A2(n_530), .B(n_531), .Y(n_529) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx4_ASAP7_75t_L g241 ( .A(n_172), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_172), .A2(n_492), .B1(n_535), .B2(n_536), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_172), .A2(n_492), .B1(n_558), .B2(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g205 ( .A(n_176), .Y(n_205) );
INVx2_ASAP7_75t_L g235 ( .A(n_176), .Y(n_235) );
OA21x2_ASAP7_75t_L g247 ( .A1(n_176), .A2(n_248), .B(n_257), .Y(n_247) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_176), .A2(n_524), .B(n_532), .Y(n_523) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_176), .A2(n_543), .B(n_550), .Y(n_542) );
INVx3_ASAP7_75t_SL g297 ( .A(n_177), .Y(n_297) );
OR2x2_ASAP7_75t_L g350 ( .A(n_177), .B(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_193), .Y(n_177) );
INVx3_ASAP7_75t_L g272 ( .A(n_178), .Y(n_272) );
AND2x2_ASAP7_75t_L g339 ( .A(n_178), .B(n_194), .Y(n_339) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_178), .Y(n_407) );
AOI33xp33_ASAP7_75t_L g411 ( .A1(n_178), .A2(n_340), .A3(n_347), .B1(n_356), .B2(n_412), .B3(n_413), .Y(n_411) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_191), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_179), .B(n_192), .Y(n_191) );
AO21x2_ASAP7_75t_L g194 ( .A1(n_179), .A2(n_195), .B(n_203), .Y(n_194) );
INVx2_ASAP7_75t_L g219 ( .A(n_179), .Y(n_219) );
INVx2_ASAP7_75t_L g202 ( .A(n_182), .Y(n_202) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
OAI22xp5_ASAP7_75t_SL g184 ( .A1(n_185), .A2(n_186), .B1(n_187), .B2(n_188), .Y(n_184) );
INVx2_ASAP7_75t_L g187 ( .A(n_185), .Y(n_187) );
INVx4_ASAP7_75t_L g253 ( .A(n_185), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g195 ( .A1(n_190), .A2(n_196), .B(n_197), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_190), .A2(n_224), .B(n_225), .Y(n_223) );
INVx1_ASAP7_75t_L g260 ( .A(n_193), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_193), .B(n_275), .Y(n_274) );
NOR3xp33_ASAP7_75t_L g334 ( .A(n_193), .B(n_335), .C(n_337), .Y(n_334) );
AND2x2_ASAP7_75t_L g360 ( .A(n_193), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_193), .B(n_367), .Y(n_370) );
AND2x2_ASAP7_75t_L g423 ( .A(n_193), .B(n_424), .Y(n_423) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx3_ASAP7_75t_L g279 ( .A(n_194), .Y(n_279) );
OR2x2_ASAP7_75t_L g373 ( .A(n_194), .B(n_272), .Y(n_373) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_201), .C(n_202), .Y(n_198) );
INVx2_ASAP7_75t_L g492 ( .A(n_200), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_200), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_200), .A2(n_507), .B(n_508), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_202), .A2(n_484), .B(n_485), .C(n_486), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_205), .B(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_205), .B(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_232), .Y(n_206) );
AOI32xp33_ASAP7_75t_L g324 ( .A1(n_207), .A2(n_325), .A3(n_327), .B1(n_329), .B2(n_332), .Y(n_324) );
NOR2xp67_ASAP7_75t_L g397 ( .A(n_207), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g427 ( .A(n_207), .Y(n_427) );
INVx4_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g359 ( .A(n_208), .B(n_343), .Y(n_359) );
AND2x2_ASAP7_75t_L g379 ( .A(n_208), .B(n_305), .Y(n_379) );
AND2x2_ASAP7_75t_L g447 ( .A(n_208), .B(n_365), .Y(n_447) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_222), .Y(n_208) );
INVx3_ASAP7_75t_L g268 ( .A(n_209), .Y(n_268) );
AND2x2_ASAP7_75t_L g282 ( .A(n_209), .B(n_266), .Y(n_282) );
OR2x2_ASAP7_75t_L g287 ( .A(n_209), .B(n_265), .Y(n_287) );
INVx1_ASAP7_75t_L g294 ( .A(n_209), .Y(n_294) );
AND2x2_ASAP7_75t_L g302 ( .A(n_209), .B(n_276), .Y(n_302) );
AND2x2_ASAP7_75t_L g304 ( .A(n_209), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_209), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g357 ( .A(n_209), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_209), .B(n_442), .Y(n_441) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_220), .Y(n_209) );
AOI21xp5_ASAP7_75t_SL g210 ( .A1(n_211), .A2(n_212), .B(n_219), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_216), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_216), .A2(n_227), .B(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g256 ( .A(n_218), .Y(n_256) );
INVx1_ASAP7_75t_L g229 ( .A(n_219), .Y(n_229) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_219), .A2(n_482), .B(n_493), .Y(n_481) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_219), .A2(n_505), .B(n_513), .Y(n_504) );
INVx2_ASAP7_75t_L g266 ( .A(n_222), .Y(n_266) );
AND2x2_ASAP7_75t_L g312 ( .A(n_222), .B(n_233), .Y(n_312) );
AND2x2_ASAP7_75t_L g322 ( .A(n_222), .B(n_247), .Y(n_322) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_229), .B(n_230), .Y(n_222) );
INVx2_ASAP7_75t_L g442 ( .A(n_232), .Y(n_442) );
OR2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_246), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_233), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g283 ( .A(n_233), .Y(n_283) );
AND2x2_ASAP7_75t_L g327 ( .A(n_233), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g343 ( .A(n_233), .B(n_306), .Y(n_343) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g291 ( .A(n_234), .Y(n_291) );
AND2x2_ASAP7_75t_L g305 ( .A(n_234), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g356 ( .A(n_234), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_234), .B(n_266), .Y(n_388) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_244), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_243), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_242), .Y(n_238) );
AND2x2_ASAP7_75t_L g267 ( .A(n_246), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g328 ( .A(n_246), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_246), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g365 ( .A(n_246), .Y(n_365) );
INVx1_ASAP7_75t_L g398 ( .A(n_246), .Y(n_398) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g276 ( .A(n_247), .B(n_266), .Y(n_276) );
INVx1_ASAP7_75t_L g306 ( .A(n_247), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_253), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g486 ( .A(n_253), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_253), .A2(n_548), .B(n_549), .Y(n_547) );
AOI221xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_263), .B1(n_269), .B2(n_276), .C(n_277), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_260), .B(n_280), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_260), .B(n_343), .Y(n_420) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_262), .B(n_310), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_262), .B(n_271), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_262), .B(n_285), .Y(n_414) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g336 ( .A(n_266), .Y(n_336) );
AND2x2_ASAP7_75t_L g311 ( .A(n_267), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g389 ( .A(n_267), .Y(n_389) );
AND2x2_ASAP7_75t_L g321 ( .A(n_268), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_268), .B(n_291), .Y(n_337) );
AND2x2_ASAP7_75t_L g401 ( .A(n_268), .B(n_327), .Y(n_401) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g310 ( .A(n_272), .B(n_279), .Y(n_310) );
AND2x2_ASAP7_75t_L g406 ( .A(n_273), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_275), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_276), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_276), .B(n_283), .Y(n_371) );
AND2x2_ASAP7_75t_L g391 ( .A(n_276), .B(n_291), .Y(n_391) );
AND2x2_ASAP7_75t_L g412 ( .A(n_276), .B(n_356), .Y(n_412) );
OAI32xp33_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_281), .A3(n_283), .B1(n_284), .B2(n_287), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_SL g285 ( .A(n_279), .Y(n_285) );
NAND2x1_ASAP7_75t_L g326 ( .A(n_279), .B(n_309), .Y(n_326) );
OR2x2_ASAP7_75t_L g330 ( .A(n_279), .B(n_331), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_279), .B(n_378), .Y(n_431) );
INVx1_ASAP7_75t_L g299 ( .A(n_280), .Y(n_299) );
OAI221xp5_ASAP7_75t_SL g417 ( .A1(n_281), .A2(n_372), .B1(n_418), .B2(n_421), .C(n_422), .Y(n_417) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g289 ( .A(n_282), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g332 ( .A(n_282), .B(n_305), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_282), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g410 ( .A(n_282), .B(n_343), .Y(n_410) );
INVxp67_ASAP7_75t_L g346 ( .A(n_283), .Y(n_346) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AND2x2_ASAP7_75t_L g416 ( .A(n_285), .B(n_403), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_285), .B(n_366), .Y(n_439) );
INVx1_ASAP7_75t_L g314 ( .A(n_287), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_287), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g432 ( .A(n_287), .B(n_433), .Y(n_432) );
OAI21xp5_ASAP7_75t_SL g288 ( .A1(n_289), .A2(n_292), .B(n_295), .Y(n_288) );
AND2x2_ASAP7_75t_L g301 ( .A(n_290), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g385 ( .A(n_294), .B(n_305), .Y(n_385) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x2_ASAP7_75t_L g403 ( .A(n_296), .B(n_361), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_296), .B(n_360), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_297), .B(n_309), .Y(n_383) );
OAI211xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_303), .C(n_313), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g333 ( .A1(n_299), .A2(n_334), .B1(n_338), .B2(n_341), .C(n_344), .Y(n_333) );
AOI31xp33_ASAP7_75t_L g428 ( .A1(n_299), .A2(n_429), .A3(n_430), .B(n_432), .Y(n_428) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_307), .B1(n_309), .B2(n_311), .Y(n_303) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g429 ( .A(n_309), .Y(n_429) );
INVx1_ASAP7_75t_L g392 ( .A(n_310), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_L g435 ( .A1(n_312), .A2(n_436), .B(n_438), .C(n_440), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B1(n_317), .B2(n_321), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_318), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OAI221xp5_ASAP7_75t_SL g408 ( .A1(n_320), .A2(n_354), .B1(n_373), .B2(n_409), .C(n_411), .Y(n_408) );
INVx1_ASAP7_75t_L g404 ( .A(n_321), .Y(n_404) );
INVx1_ASAP7_75t_L g358 ( .A(n_322), .Y(n_358) );
NAND3xp33_ASAP7_75t_SL g323 ( .A(n_324), .B(n_333), .C(n_348), .Y(n_323) );
OAI21xp33_ASAP7_75t_L g374 ( .A1(n_325), .A2(n_375), .B(n_379), .Y(n_374) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_327), .B(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g434 ( .A(n_328), .Y(n_434) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g372 ( .A(n_335), .B(n_355), .Y(n_372) );
INVx1_ASAP7_75t_L g347 ( .A(n_336), .Y(n_347) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g345 ( .A(n_339), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_339), .B(n_377), .Y(n_376) );
NOR4xp25_ASAP7_75t_L g344 ( .A(n_340), .B(n_345), .C(n_346), .D(n_347), .Y(n_344) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI222xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_353), .B1(n_359), .B2(n_360), .C1(n_362), .C2(n_366), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_350), .B(n_352), .Y(n_349) );
INVx1_ASAP7_75t_L g446 ( .A(n_350), .Y(n_446) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_358), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_362), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI21xp5_ASAP7_75t_SL g422 ( .A1(n_367), .A2(n_423), .B(n_425), .Y(n_422) );
NOR4xp25_ASAP7_75t_L g368 ( .A(n_369), .B(n_380), .C(n_393), .D(n_408), .Y(n_368) );
OAI221xp5_ASAP7_75t_SL g369 ( .A1(n_370), .A2(n_371), .B1(n_372), .B2(n_373), .C(n_374), .Y(n_369) );
INVx1_ASAP7_75t_L g449 ( .A(n_370), .Y(n_449) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_377), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
OAI222xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_384), .B1(n_386), .B2(n_387), .C1(n_390), .C2(n_392), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI211xp5_ASAP7_75t_L g415 ( .A1(n_385), .A2(n_416), .B(n_417), .C(n_428), .Y(n_415) );
OR2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
OAI222xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_399), .B1(n_400), .B2(n_402), .C1(n_404), .C2(n_405), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_410), .A2(n_413), .B1(n_446), .B2(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI211xp5_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_443), .B(n_445), .C(n_448), .Y(n_440) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g460 ( .A(n_453), .Y(n_460) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
AOI21xp33_ASAP7_75t_L g461 ( .A1(n_459), .A2(n_462), .B(n_775), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_467), .A2(n_472), .B1(n_773), .B2(n_774), .Y(n_772) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx6_ASAP7_75t_L g774 ( .A(n_470), .Y(n_774) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_SL g472 ( .A(n_473), .B(n_729), .Y(n_472) );
NOR3xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_633), .C(n_717), .Y(n_473) );
NAND4xp25_ASAP7_75t_L g474 ( .A(n_475), .B(n_576), .C(n_598), .D(n_614), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_514), .B1(n_537), .B2(n_555), .C(n_562), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_494), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_478), .B(n_555), .Y(n_588) );
NAND4xp25_ASAP7_75t_L g628 ( .A(n_478), .B(n_616), .C(n_629), .D(n_631), .Y(n_628) );
INVxp67_ASAP7_75t_L g745 ( .A(n_478), .Y(n_745) );
INVx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OR2x2_ASAP7_75t_L g627 ( .A(n_479), .B(n_565), .Y(n_627) );
AND2x2_ASAP7_75t_L g651 ( .A(n_479), .B(n_494), .Y(n_651) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g618 ( .A(n_480), .B(n_554), .Y(n_618) );
AND2x2_ASAP7_75t_L g658 ( .A(n_480), .B(n_639), .Y(n_658) );
AND2x2_ASAP7_75t_L g675 ( .A(n_480), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_480), .B(n_495), .Y(n_699) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g553 ( .A(n_481), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g570 ( .A(n_481), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g582 ( .A(n_481), .B(n_495), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_481), .B(n_504), .Y(n_604) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_490), .B(n_491), .C(n_492), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_492), .A2(n_501), .B(n_502), .Y(n_500) );
AND2x2_ASAP7_75t_L g585 ( .A(n_494), .B(n_586), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_494), .A2(n_635), .B1(n_638), .B2(n_640), .C(n_644), .Y(n_634) );
AND2x2_ASAP7_75t_L g693 ( .A(n_494), .B(n_658), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_494), .B(n_675), .Y(n_727) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_504), .Y(n_494) );
INVx3_ASAP7_75t_L g554 ( .A(n_495), .Y(n_554) );
AND2x2_ASAP7_75t_L g602 ( .A(n_495), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g656 ( .A(n_495), .B(n_571), .Y(n_656) );
AND2x2_ASAP7_75t_L g714 ( .A(n_495), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g555 ( .A(n_504), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g571 ( .A(n_504), .Y(n_571) );
INVx1_ASAP7_75t_L g626 ( .A(n_504), .Y(n_626) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_504), .Y(n_632) );
AND2x2_ASAP7_75t_L g677 ( .A(n_504), .B(n_554), .Y(n_677) );
OR2x2_ASAP7_75t_L g716 ( .A(n_504), .B(n_556), .Y(n_716) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_509), .B(n_512), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_514), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_522), .Y(n_514) );
AND2x2_ASAP7_75t_L g712 ( .A(n_515), .B(n_709), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_515), .B(n_694), .Y(n_744) );
BUFx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g643 ( .A(n_516), .B(n_567), .Y(n_643) );
AND2x2_ASAP7_75t_L g692 ( .A(n_516), .B(n_540), .Y(n_692) );
INVx1_ASAP7_75t_L g738 ( .A(n_516), .Y(n_738) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_517), .Y(n_552) );
AND2x2_ASAP7_75t_L g593 ( .A(n_517), .B(n_567), .Y(n_593) );
INVx1_ASAP7_75t_L g610 ( .A(n_517), .Y(n_610) );
AND2x2_ASAP7_75t_L g616 ( .A(n_517), .B(n_533), .Y(n_616) );
AND2x2_ASAP7_75t_L g684 ( .A(n_522), .B(n_592), .Y(n_684) );
INVx2_ASAP7_75t_L g749 ( .A(n_522), .Y(n_749) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_533), .Y(n_522) );
AND2x2_ASAP7_75t_L g566 ( .A(n_523), .B(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g579 ( .A(n_523), .B(n_541), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_523), .B(n_540), .Y(n_607) );
INVx1_ASAP7_75t_L g613 ( .A(n_523), .Y(n_613) );
INVx1_ASAP7_75t_L g630 ( .A(n_523), .Y(n_630) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_523), .Y(n_642) );
INVx2_ASAP7_75t_L g710 ( .A(n_523), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B(n_528), .Y(n_525) );
INVx2_ASAP7_75t_L g567 ( .A(n_533), .Y(n_567) );
BUFx2_ASAP7_75t_L g664 ( .A(n_533), .Y(n_664) );
AND2x2_ASAP7_75t_L g709 ( .A(n_533), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_551), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_539), .B(n_646), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_539), .A2(n_708), .B(n_722), .Y(n_732) );
AND2x2_ASAP7_75t_L g757 ( .A(n_539), .B(n_643), .Y(n_757) );
BUFx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g679 ( .A(n_541), .Y(n_679) );
AND2x2_ASAP7_75t_L g708 ( .A(n_541), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_542), .Y(n_592) );
INVx2_ASAP7_75t_L g611 ( .A(n_542), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_542), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx2_ASAP7_75t_L g565 ( .A(n_552), .Y(n_565) );
OR2x2_ASAP7_75t_L g578 ( .A(n_552), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g646 ( .A(n_552), .B(n_642), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_552), .B(n_742), .Y(n_741) );
OR2x2_ASAP7_75t_L g747 ( .A(n_552), .B(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_552), .B(n_684), .Y(n_759) );
AND2x2_ASAP7_75t_L g638 ( .A(n_553), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g661 ( .A(n_553), .B(n_555), .Y(n_661) );
INVx2_ASAP7_75t_L g573 ( .A(n_554), .Y(n_573) );
AND2x2_ASAP7_75t_L g601 ( .A(n_554), .B(n_574), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_554), .B(n_626), .Y(n_682) );
AND2x2_ASAP7_75t_L g596 ( .A(n_555), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g743 ( .A(n_555), .Y(n_743) );
AND2x2_ASAP7_75t_L g755 ( .A(n_555), .B(n_618), .Y(n_755) );
AND2x2_ASAP7_75t_L g581 ( .A(n_556), .B(n_571), .Y(n_581) );
INVx1_ASAP7_75t_L g676 ( .A(n_556), .Y(n_676) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x4_ASAP7_75t_L g574 ( .A(n_561), .B(n_575), .Y(n_574) );
INVxp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_568), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_565), .B(n_612), .Y(n_621) );
OR2x2_ASAP7_75t_L g753 ( .A(n_565), .B(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g670 ( .A(n_566), .B(n_611), .Y(n_670) );
AND2x2_ASAP7_75t_L g678 ( .A(n_566), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g737 ( .A(n_566), .B(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g761 ( .A(n_566), .B(n_608), .Y(n_761) );
NOR2xp67_ASAP7_75t_L g719 ( .A(n_567), .B(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g748 ( .A(n_567), .B(n_611), .Y(n_748) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2x1p5_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
AND2x2_ASAP7_75t_L g600 ( .A(n_570), .B(n_601), .Y(n_600) );
INVxp67_ASAP7_75t_L g762 ( .A(n_570), .Y(n_762) );
NOR2x1_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g597 ( .A(n_573), .Y(n_597) );
AND2x2_ASAP7_75t_L g648 ( .A(n_573), .B(n_581), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_573), .B(n_716), .Y(n_742) );
INVx2_ASAP7_75t_L g587 ( .A(n_574), .Y(n_587) );
INVx3_ASAP7_75t_L g639 ( .A(n_574), .Y(n_639) );
OR2x2_ASAP7_75t_L g667 ( .A(n_574), .B(n_668), .Y(n_667) );
AOI311xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_580), .A3(n_582), .B(n_583), .C(n_594), .Y(n_576) );
O2A1O1Ixp33_ASAP7_75t_L g614 ( .A1(n_577), .A2(n_615), .B(n_617), .C(n_619), .Y(n_614) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_SL g599 ( .A(n_579), .Y(n_599) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g617 ( .A(n_581), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_581), .B(n_597), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_581), .B(n_582), .Y(n_750) );
AND2x2_ASAP7_75t_L g672 ( .A(n_582), .B(n_586), .Y(n_672) );
AOI21xp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_588), .B(n_589), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g730 ( .A(n_586), .B(n_618), .Y(n_730) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_587), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g624 ( .A(n_587), .Y(n_624) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
AND2x2_ASAP7_75t_L g615 ( .A(n_591), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g660 ( .A(n_593), .Y(n_660) );
AND2x4_ASAP7_75t_L g722 ( .A(n_593), .B(n_691), .Y(n_722) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AOI222xp33_ASAP7_75t_L g673 ( .A1(n_596), .A2(n_662), .B1(n_674), .B2(n_678), .C1(n_680), .C2(n_684), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_600), .B(n_602), .C(n_605), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_599), .B(n_643), .Y(n_666) );
INVx1_ASAP7_75t_L g688 ( .A(n_601), .Y(n_688) );
INVx1_ASAP7_75t_L g622 ( .A(n_603), .Y(n_622) );
OR2x2_ASAP7_75t_L g687 ( .A(n_604), .B(n_688), .Y(n_687) );
OAI21xp33_ASAP7_75t_SL g605 ( .A1(n_606), .A2(n_608), .B(n_612), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_606), .B(n_624), .C(n_625), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_606), .A2(n_643), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_610), .Y(n_663) );
AND2x2_ASAP7_75t_SL g629 ( .A(n_611), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g720 ( .A(n_611), .Y(n_720) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_611), .Y(n_736) );
INVx2_ASAP7_75t_L g694 ( .A(n_612), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_616), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g668 ( .A(n_618), .Y(n_668) );
OAI221xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_622), .B1(n_623), .B2(n_627), .C(n_628), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_622), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g756 ( .A(n_622), .Y(n_756) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g637 ( .A(n_629), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_629), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g695 ( .A(n_629), .B(n_643), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_629), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g728 ( .A(n_629), .B(n_663), .Y(n_728) );
BUFx3_ASAP7_75t_L g691 ( .A(n_630), .Y(n_691) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND5xp2_ASAP7_75t_L g633 ( .A(n_634), .B(n_652), .C(n_673), .D(n_685), .E(n_700), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AOI32xp33_ASAP7_75t_L g725 ( .A1(n_637), .A2(n_664), .A3(n_680), .B1(n_726), .B2(n_728), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_639), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g649 ( .A(n_643), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_647), .B1(n_649), .B2(n_650), .Y(n_644) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_659), .B1(n_661), .B2(n_662), .C(n_665), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g724 ( .A(n_656), .B(n_675), .Y(n_724) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g739 ( .A1(n_661), .A2(n_722), .B1(n_740), .B2(n_745), .C(n_746), .Y(n_739) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx2_ASAP7_75t_L g705 ( .A(n_664), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B1(n_669), .B2(n_671), .Y(n_665) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
INVx1_ASAP7_75t_L g683 ( .A(n_675), .Y(n_683) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
AOI222xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_689), .B1(n_693), .B2(n_694), .C1(n_695), .C2(n_696), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_692), .Y(n_689) );
INVxp67_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OAI22xp33_ASAP7_75t_L g740 ( .A1(n_694), .A2(n_741), .B1(n_743), .B2(n_744), .Y(n_740) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_703), .B(n_706), .Y(n_700) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI21xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_711), .B(n_713), .Y(n_706) );
INVx2_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g754 ( .A(n_709), .Y(n_754) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_721), .B(n_723), .C(n_725), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AOI211xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B(n_733), .C(n_758), .Y(n_729) );
CKINVDCx16_ASAP7_75t_R g734 ( .A(n_730), .Y(n_734) );
INVxp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI211xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B(n_739), .C(n_751), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
AOI21xp33_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_749), .B(n_750), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AOI21xp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B(n_762), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g768 ( .A(n_765), .Y(n_768) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
endmodule