module real_aes_12853_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_919;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_961;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_938;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_656;
wire n_316;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_936;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_713;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_649;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_155;
wire n_653;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_949;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx2_ASAP7_75t_SL g171 ( .A(n_0), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_1), .Y(n_333) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_2), .A2(n_51), .B(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g179 ( .A(n_2), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_3), .B(n_166), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_4), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_5), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_6), .B(n_198), .Y(n_659) );
AND2x2_ASAP7_75t_L g272 ( .A(n_7), .B(n_189), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_8), .B(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_9), .B(n_220), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_10), .B(n_220), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g958 ( .A(n_11), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_12), .B(n_631), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_13), .B(n_152), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_14), .B(n_284), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_15), .B(n_169), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_16), .Y(n_678) );
BUFx3_ASAP7_75t_L g148 ( .A(n_17), .Y(n_148) );
INVx1_ASAP7_75t_L g154 ( .A(n_17), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_18), .B(n_188), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_19), .B(n_260), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_20), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g656 ( .A(n_21), .Y(n_656) );
BUFx10_ASAP7_75t_L g581 ( .A(n_22), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_23), .B(n_228), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_24), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_25), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_26), .B(n_619), .Y(n_643) );
NAND3xp33_ASAP7_75t_L g248 ( .A(n_27), .B(n_246), .C(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_28), .B(n_228), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_29), .B(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_30), .B(n_260), .Y(n_711) );
NAND2xp33_ASAP7_75t_L g622 ( .A(n_31), .B(n_147), .Y(n_622) );
INVx1_ASAP7_75t_L g183 ( .A(n_32), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g669 ( .A1(n_33), .A2(n_262), .B(n_338), .C(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_34), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_35), .B(n_335), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_36), .B(n_166), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_37), .A2(n_58), .B1(n_940), .B2(n_941), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_37), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_38), .B(n_311), .Y(n_649) );
INVx1_ASAP7_75t_L g112 ( .A(n_39), .Y(n_112) );
AND3x2_ASAP7_75t_L g956 ( .A(n_39), .B(n_948), .C(n_949), .Y(n_956) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_40), .B(n_222), .Y(n_221) );
AO221x1_ASAP7_75t_L g628 ( .A1(n_41), .A2(n_84), .B1(n_146), .B2(n_228), .C(n_310), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_42), .B(n_646), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_43), .B(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_L g182 ( .A(n_44), .B(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_45), .B(n_188), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g952 ( .A(n_46), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_47), .B(n_161), .Y(n_160) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_48), .B(n_337), .C(n_338), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_49), .B(n_188), .Y(n_187) );
AOI22x1_ASAP7_75t_SL g568 ( .A1(n_50), .A2(n_89), .B1(n_569), .B2(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_50), .Y(n_570) );
INVx1_ASAP7_75t_L g178 ( .A(n_51), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_52), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_53), .A2(n_165), .B(n_168), .C(n_172), .Y(n_164) );
INVx1_ASAP7_75t_L g163 ( .A(n_54), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g675 ( .A(n_55), .Y(n_675) );
A2O1A1Ixp33_ASAP7_75t_L g682 ( .A1(n_56), .A2(n_683), .B(n_684), .C(n_686), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_57), .B(n_188), .Y(n_339) );
INVx1_ASAP7_75t_L g941 ( .A(n_58), .Y(n_941) );
INVx2_ASAP7_75t_L g685 ( .A(n_59), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_60), .B(n_161), .Y(n_661) );
AND2x4_ASAP7_75t_L g109 ( .A(n_61), .B(n_110), .Y(n_109) );
INVx3_ASAP7_75t_L g294 ( .A(n_62), .Y(n_294) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_63), .Y(n_117) );
NOR2xp67_ASAP7_75t_L g127 ( .A(n_63), .B(n_75), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_64), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g110 ( .A(n_65), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_66), .B(n_194), .Y(n_203) );
INVx1_ASAP7_75t_L g309 ( .A(n_67), .Y(n_309) );
AND2x2_ASAP7_75t_L g651 ( .A(n_68), .B(n_161), .Y(n_651) );
INVx1_ASAP7_75t_L g634 ( .A(n_69), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_70), .B(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g125 ( .A(n_70), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_71), .B(n_241), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_72), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g330 ( .A(n_73), .B(n_249), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g630 ( .A1(n_74), .A2(n_77), .B1(n_619), .B2(n_631), .Y(n_630) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_75), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_76), .B(n_338), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_78), .B(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g149 ( .A(n_79), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_80), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_81), .B(n_315), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g936 ( .A1(n_82), .A2(n_937), .B1(n_938), .B2(n_939), .Y(n_936) );
CKINVDCx5p33_ASAP7_75t_R g937 ( .A(n_82), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_83), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g692 ( .A(n_85), .B(n_189), .Y(n_692) );
INVx1_ASAP7_75t_L g158 ( .A(n_86), .Y(n_158) );
INVx1_ASAP7_75t_L g174 ( .A(n_86), .Y(n_174) );
BUFx3_ASAP7_75t_L g284 ( .A(n_86), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_87), .B(n_241), .Y(n_331) );
INVx1_ASAP7_75t_L g292 ( .A(n_88), .Y(n_292) );
INVx1_ASAP7_75t_L g569 ( .A(n_89), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_90), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_91), .B(n_176), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_92), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_93), .B(n_189), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_94), .B(n_646), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_95), .B(n_161), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_96), .B(n_201), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_97), .Y(n_287) );
INVx1_ASAP7_75t_L g282 ( .A(n_98), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g716 ( .A(n_99), .Y(n_716) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_100), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_101), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_102), .B(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_118), .B(n_957), .Y(n_103) );
BUFx4f_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND3x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_113), .C(n_116), .Y(n_105) );
AND3x4_ASAP7_75t_L g961 ( .A(n_106), .B(n_113), .C(n_116), .Y(n_961) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_111), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g587 ( .A(n_111), .Y(n_587) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_112), .B(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OR2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_128), .Y(n_118) );
INVxp67_ASAP7_75t_L g580 ( .A(n_119), .Y(n_580) );
NOR2xp67_ASAP7_75t_SL g119 ( .A(n_120), .B(n_121), .Y(n_119) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_SL g574 ( .A(n_123), .Y(n_574) );
NOR2x1p5_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx2_ASAP7_75t_L g949 ( .A(n_125), .Y(n_949) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_127), .Y(n_948) );
OAI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_581), .B(n_582), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_131), .B(n_575), .Y(n_129) );
OAI31xp33_ASAP7_75t_L g575 ( .A1(n_130), .A2(n_132), .A3(n_576), .B(n_580), .Y(n_575) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_572), .Y(n_131) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_134), .B1(n_568), .B2(n_571), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g588 ( .A(n_134), .Y(n_588) );
AND3x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_472), .C(n_518), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_416), .Y(n_135) );
NAND3xp33_ASAP7_75t_SL g136 ( .A(n_137), .B(n_353), .C(n_388), .Y(n_136) );
AOI22xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_211), .B1(n_340), .B2(n_347), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_184), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g468 ( .A(n_141), .B(n_214), .Y(n_468) );
AND2x4_ASAP7_75t_L g481 ( .A(n_141), .B(n_376), .Y(n_481) );
AND2x2_ASAP7_75t_L g512 ( .A(n_141), .B(n_397), .Y(n_512) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_141), .Y(n_545) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OR2x6_ASAP7_75t_L g365 ( .A(n_142), .B(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_SL g377 ( .A(n_142), .B(n_344), .Y(n_377) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g343 ( .A(n_143), .Y(n_343) );
OAI21x1_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_159), .B(n_175), .Y(n_143) );
AOI21x1_ASAP7_75t_SL g144 ( .A1(n_145), .A2(n_150), .B(n_155), .Y(n_144) );
OR2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_149), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g220 ( .A(n_147), .Y(n_220) );
INVx2_ASAP7_75t_L g241 ( .A(n_147), .Y(n_241) );
INVx3_ASAP7_75t_L g260 ( .A(n_147), .Y(n_260) );
INVx2_ASAP7_75t_L g266 ( .A(n_147), .Y(n_266) );
INVx2_ASAP7_75t_L g335 ( .A(n_147), .Y(n_335) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_148), .Y(n_170) );
INVx2_ASAP7_75t_L g250 ( .A(n_148), .Y(n_250) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g222 ( .A(n_152), .Y(n_222) );
INVx2_ASAP7_75t_L g225 ( .A(n_152), .Y(n_225) );
INVx2_ASAP7_75t_L g243 ( .A(n_152), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_152), .B(n_678), .Y(n_677) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_153), .Y(n_228) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_154), .Y(n_167) );
AOI22x1_ASAP7_75t_L g257 ( .A1(n_155), .A2(n_173), .B1(n_258), .B2(n_264), .Y(n_257) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_156), .A2(n_193), .B(n_196), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_156), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g289 ( .A(n_157), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_157), .A2(n_617), .B(n_618), .Y(n_616) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx3_ASAP7_75t_L g205 ( .A(n_158), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_164), .Y(n_159) );
OAI21xp33_ASAP7_75t_L g175 ( .A1(n_160), .A2(n_176), .B(n_181), .Y(n_175) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_161), .Y(n_207) );
INVx1_ASAP7_75t_L g346 ( .A(n_161), .Y(n_346) );
INVxp67_ASAP7_75t_SL g602 ( .A(n_161), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_161), .B(n_285), .Y(n_612) );
INVx2_ASAP7_75t_L g641 ( .A(n_161), .Y(n_641) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g190 ( .A(n_162), .Y(n_190) );
BUFx2_ASAP7_75t_L g302 ( .A(n_162), .Y(n_302) );
INVx1_ASAP7_75t_L g180 ( .A(n_163), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_165), .A2(n_265), .B1(n_267), .B2(n_268), .Y(n_264) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g198 ( .A(n_167), .Y(n_198) );
INVx1_ASAP7_75t_L g202 ( .A(n_167), .Y(n_202) );
INVx2_ASAP7_75t_L g337 ( .A(n_167), .Y(n_337) );
INVx1_ASAP7_75t_L g676 ( .A(n_167), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_171), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g195 ( .A(n_170), .Y(n_195) );
INVx1_ASAP7_75t_L g315 ( .A(n_170), .Y(n_315) );
INVx2_ASAP7_75t_L g631 ( .A(n_170), .Y(n_631) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AOI21x1_ASAP7_75t_L g239 ( .A1(n_173), .A2(n_240), .B(n_242), .Y(n_239) );
AOI21xp5_ASAP7_75t_SL g642 ( .A1(n_173), .A2(n_643), .B(n_644), .Y(n_642) );
BUFx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g230 ( .A(n_174), .Y(n_230) );
INVxp67_ASAP7_75t_L g269 ( .A(n_176), .Y(n_269) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_177), .B(n_209), .Y(n_667) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_180), .Y(n_177) );
AOI21x1_ASAP7_75t_L g278 ( .A1(n_178), .A2(n_179), .B(n_180), .Y(n_278) );
INVx1_ASAP7_75t_L g271 ( .A(n_181), .Y(n_271) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g210 ( .A(n_182), .Y(n_210) );
BUFx6f_ASAP7_75t_SL g231 ( .A(n_182), .Y(n_231) );
INVx3_ASAP7_75t_L g285 ( .A(n_182), .Y(n_285) );
OR2x2_ASAP7_75t_L g457 ( .A(n_184), .B(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g478 ( .A(n_184), .B(n_365), .Y(n_478) );
BUFx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g385 ( .A(n_185), .Y(n_385) );
AND2x2_ASAP7_75t_L g392 ( .A(n_185), .B(n_344), .Y(n_392) );
INVx2_ASAP7_75t_L g397 ( .A(n_185), .Y(n_397) );
AND2x2_ASAP7_75t_L g412 ( .A(n_185), .B(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g422 ( .A(n_185), .B(n_234), .Y(n_422) );
OR2x2_ASAP7_75t_L g438 ( .A(n_185), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g467 ( .A(n_185), .Y(n_467) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NAND2x1_ASAP7_75t_L g186 ( .A(n_187), .B(n_191), .Y(n_186) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_188), .Y(n_237) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OAI21x1_ASAP7_75t_SL g191 ( .A1(n_192), .A2(n_199), .B(n_206), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_194), .A2(n_291), .B1(n_293), .B2(n_295), .Y(n_290) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_195), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_203), .B(n_204), .Y(n_199) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_205), .A2(n_219), .B(n_221), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_205), .A2(n_621), .B(n_622), .Y(n_620) );
INVx1_ASAP7_75t_L g686 ( .A(n_205), .Y(n_686) );
NOR2x1_ASAP7_75t_SL g206 ( .A(n_207), .B(n_208), .Y(n_206) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_207), .Y(n_216) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g251 ( .A(n_210), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_253), .B1(n_317), .B2(n_321), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
OR2x2_ASAP7_75t_L g505 ( .A(n_213), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_233), .Y(n_213) );
BUFx3_ASAP7_75t_L g319 ( .A(n_214), .Y(n_319) );
AND2x2_ASAP7_75t_L g410 ( .A(n_214), .B(n_385), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_214), .Y(n_413) );
AND2x2_ASAP7_75t_L g527 ( .A(n_214), .B(n_343), .Y(n_527) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_215), .Y(n_449) );
OAI21x1_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_232), .Y(n_215) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_216), .A2(n_257), .B(n_351), .Y(n_350) );
OAI21x1_ASAP7_75t_L g376 ( .A1(n_216), .A2(n_217), .B(n_232), .Y(n_376) );
OAI21x1_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_223), .B(n_231), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_226), .B(n_229), .Y(n_223) );
INVx2_ASAP7_75t_L g262 ( .A(n_225), .Y(n_262) );
INVxp67_ASAP7_75t_L g247 ( .A(n_227), .Y(n_247) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_228), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g295 ( .A(n_228), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_229), .A2(n_313), .B(n_314), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_229), .A2(n_330), .B(n_331), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_229), .A2(n_649), .B(n_650), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_229), .A2(n_659), .B(n_660), .Y(n_658) );
INVx1_ASAP7_75t_L g691 ( .A(n_229), .Y(n_691) );
BUFx10_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g246 ( .A(n_230), .Y(n_246) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_231), .A2(n_304), .B(n_312), .Y(n_303) );
OAI21x1_ASAP7_75t_L g654 ( .A1(n_231), .A2(n_655), .B(n_658), .Y(n_654) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_233), .Y(n_425) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_234), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_234), .B(n_343), .Y(n_458) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g366 ( .A(n_235), .Y(n_366) );
INVxp67_ASAP7_75t_SL g439 ( .A(n_235), .Y(n_439) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OAI21x1_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_252), .Y(n_236) );
OA21x2_ASAP7_75t_L g344 ( .A1(n_238), .A2(n_252), .B(n_345), .Y(n_344) );
OAI21x1_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_244), .B(n_251), .Y(n_238) );
O2A1O1Ixp5_ASAP7_75t_L g655 ( .A1(n_243), .A2(n_611), .B(n_656), .C(n_657), .Y(n_655) );
OAI21xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_247), .B(n_248), .Y(n_244) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g311 ( .A(n_250), .Y(n_311) );
INVx2_ASAP7_75t_L g619 ( .A(n_250), .Y(n_619) );
INVx2_ASAP7_75t_L g646 ( .A(n_250), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g328 ( .A1(n_251), .A2(n_329), .B(n_332), .Y(n_328) );
INVx2_ASAP7_75t_L g418 ( .A(n_253), .Y(n_418) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_273), .Y(n_253) );
INVx1_ASAP7_75t_L g383 ( .A(n_254), .Y(n_383) );
INVx1_ASAP7_75t_L g415 ( .A(n_254), .Y(n_415) );
BUFx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g401 ( .A(n_255), .Y(n_401) );
AO31x2_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_269), .A3(n_270), .B(n_272), .Y(n_255) );
AO31x2_ASAP7_75t_L g433 ( .A1(n_256), .A2(n_269), .A3(n_270), .B(n_272), .Y(n_433) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OAI22x1_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_261), .B1(n_262), .B2(n_263), .Y(n_258) );
INVxp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVxp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVxp67_ASAP7_75t_L g305 ( .A(n_266), .Y(n_305) );
BUFx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g351 ( .A(n_272), .Y(n_351) );
INVx1_ASAP7_75t_L g551 ( .A(n_273), .Y(n_551) );
INVxp67_ASAP7_75t_SL g562 ( .A(n_273), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_298), .Y(n_273) );
NOR2x1_ASAP7_75t_L g324 ( .A(n_274), .B(n_325), .Y(n_324) );
BUFx2_ASAP7_75t_L g387 ( .A(n_274), .Y(n_387) );
INVx1_ASAP7_75t_L g429 ( .A(n_274), .Y(n_429) );
AND2x2_ASAP7_75t_L g488 ( .A(n_274), .B(n_299), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_274), .B(n_352), .Y(n_510) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g348 ( .A(n_275), .B(n_299), .Y(n_348) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_279), .B(n_296), .Y(n_275) );
AO21x1_ASAP7_75t_L g361 ( .A1(n_276), .A2(n_279), .B(n_296), .Y(n_361) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_SL g296 ( .A(n_277), .B(n_297), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_277), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_R g632 ( .A(n_278), .B(n_285), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_290), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_283), .B1(n_286), .B2(n_288), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
NOR3xp33_ASAP7_75t_L g291 ( .A(n_284), .B(n_285), .C(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g310 ( .A(n_284), .Y(n_310) );
INVx2_ASAP7_75t_L g338 ( .A(n_284), .Y(n_338) );
INVx1_ASAP7_75t_L g611 ( .A(n_284), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_285), .B(n_289), .Y(n_288) );
NOR3xp33_ASAP7_75t_L g293 ( .A(n_285), .B(n_289), .C(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g623 ( .A(n_285), .Y(n_623) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_299), .Y(n_323) );
INVx3_ASAP7_75t_L g357 ( .A(n_299), .Y(n_357) );
INVx2_ASAP7_75t_L g370 ( .A(n_299), .Y(n_370) );
AND2x2_ASAP7_75t_L g374 ( .A(n_299), .B(n_350), .Y(n_374) );
INVx1_ASAP7_75t_L g398 ( .A(n_299), .Y(n_398) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_303), .B(n_316), .Y(n_300) );
OAI21x1_ASAP7_75t_L g327 ( .A1(n_301), .A2(n_328), .B(n_339), .Y(n_327) );
OAI21x1_ASAP7_75t_L g653 ( .A1(n_301), .A2(n_654), .B(n_661), .Y(n_653) );
BUFx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVxp67_ASAP7_75t_L g694 ( .A(n_302), .Y(n_694) );
OAI21xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_306), .B(n_307), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_311), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g607 ( .A(n_310), .Y(n_607) );
INVxp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_319), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g436 ( .A(n_319), .Y(n_436) );
OR2x2_ASAP7_75t_L g477 ( .A(n_319), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
OR2x2_ASAP7_75t_L g557 ( .A(n_322), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g373 ( .A(n_325), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_325), .B(n_357), .Y(n_406) );
NOR2xp67_ASAP7_75t_L g516 ( .A(n_325), .B(n_356), .Y(n_516) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx3_ASAP7_75t_L g352 ( .A(n_326), .Y(n_352) );
AND2x2_ASAP7_75t_L g359 ( .A(n_326), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g471 ( .A(n_326), .B(n_350), .Y(n_471) );
INVx1_ASAP7_75t_L g494 ( .A(n_326), .Y(n_494) );
INVx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
O2A1O1Ixp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_334), .B(n_336), .C(n_338), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g712 ( .A1(n_334), .A2(n_713), .B(n_714), .Y(n_712) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI211xp5_ASAP7_75t_L g353 ( .A1(n_342), .A2(n_354), .B(n_362), .C(n_378), .Y(n_353) );
AND2x2_ASAP7_75t_L g502 ( .A(n_342), .B(n_466), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_342), .B(n_397), .Y(n_555) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g381 ( .A(n_343), .Y(n_381) );
AND2x4_ASAP7_75t_L g391 ( .A(n_343), .B(n_376), .Y(n_391) );
OA21x2_ASAP7_75t_L g614 ( .A1(n_345), .A2(n_615), .B(n_624), .Y(n_614) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
AOI32xp33_ASAP7_75t_L g479 ( .A1(n_347), .A2(n_421), .A3(n_480), .B1(n_482), .B2(n_484), .Y(n_479) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
AND2x2_ASAP7_75t_L g470 ( .A(n_348), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g371 ( .A(n_349), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_349), .B(n_429), .Y(n_445) );
AND2x2_ASAP7_75t_L g498 ( .A(n_349), .B(n_387), .Y(n_498) );
AND2x2_ASAP7_75t_L g561 ( .A(n_349), .B(n_562), .Y(n_561) );
AND2x4_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
INVx1_ASAP7_75t_L g408 ( .A(n_350), .Y(n_408) );
OR2x2_ASAP7_75t_L g432 ( .A(n_352), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
AOI21xp33_ASAP7_75t_SL g451 ( .A1(n_355), .A2(n_409), .B(n_450), .Y(n_451) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
BUFx2_ASAP7_75t_L g496 ( .A(n_356), .Y(n_496) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_357), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g461 ( .A(n_357), .B(n_433), .Y(n_461) );
INVx1_ASAP7_75t_L g395 ( .A(n_358), .Y(n_395) );
OR2x2_ASAP7_75t_L g441 ( .A(n_358), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g400 ( .A(n_359), .Y(n_400) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_359), .Y(n_462) );
AND2x2_ASAP7_75t_L g503 ( .A(n_359), .B(n_401), .Y(n_503) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g369 ( .A(n_361), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_361), .B(n_408), .Y(n_407) );
OAI22xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_367), .B1(n_372), .B2(n_375), .Y(n_362) );
INVxp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2x1p5_ASAP7_75t_L g411 ( .A(n_364), .B(n_412), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_364), .A2(n_534), .B1(n_536), .B2(n_538), .Y(n_533) );
INVx2_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g454 ( .A(n_365), .B(n_397), .Y(n_454) );
AND2x2_ASAP7_75t_L g382 ( .A(n_366), .B(n_376), .Y(n_382) );
INVx2_ASAP7_75t_L g567 ( .A(n_367), .Y(n_567) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_371), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g475 ( .A(n_369), .B(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g484 ( .A(n_369), .B(n_471), .Y(n_484) );
AND2x2_ASAP7_75t_L g523 ( .A(n_369), .B(n_415), .Y(n_523) );
AND2x2_ASAP7_75t_L g542 ( .A(n_369), .B(n_506), .Y(n_542) );
INVx1_ASAP7_75t_L g389 ( .A(n_371), .Y(n_389) );
OAI321xp33_ASAP7_75t_L g559 ( .A1(n_372), .A2(n_448), .A3(n_482), .B1(n_560), .B2(n_563), .C(n_566), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_373), .B(n_374), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_373), .B(n_515), .Y(n_558) );
INVx1_ASAP7_75t_L g442 ( .A(n_374), .Y(n_442) );
AND2x4_ASAP7_75t_L g508 ( .A(n_374), .B(n_509), .Y(n_508) );
INVx3_ASAP7_75t_L g529 ( .A(n_375), .Y(n_529) );
OR2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
AND2x4_ASAP7_75t_L g421 ( .A(n_376), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g403 ( .A(n_377), .Y(n_403) );
NOR4xp25_ASAP7_75t_L g378 ( .A(n_379), .B(n_383), .C(n_384), .D(n_386), .Y(n_378) );
NAND2x1_ASAP7_75t_L g419 ( .A(n_379), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_380), .A2(n_455), .B1(n_502), .B2(n_503), .Y(n_501) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
OAI322xp33_ASAP7_75t_L g540 ( .A1(n_383), .A2(n_541), .A3(n_543), .B1(n_549), .B2(n_552), .C1(n_553), .C2(n_557), .Y(n_540) );
AND2x2_ASAP7_75t_L g500 ( .A(n_384), .B(n_468), .Y(n_500) );
BUFx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g483 ( .A(n_385), .B(n_439), .Y(n_483) );
INVx1_ASAP7_75t_L g506 ( .A(n_385), .Y(n_506) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2x1_ASAP7_75t_L g455 ( .A(n_387), .B(n_432), .Y(n_455) );
AOI211xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B(n_393), .C(n_404), .Y(n_388) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_L g464 ( .A(n_391), .Y(n_464) );
NOR2x1_ASAP7_75t_L g564 ( .A(n_391), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g450 ( .A(n_392), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_SL g393 ( .A1(n_394), .A2(n_396), .B(n_399), .C(n_402), .Y(n_393) );
INVxp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
AND2x2_ASAP7_75t_L g556 ( .A(n_397), .B(n_527), .Y(n_556) );
INVx2_ASAP7_75t_L g431 ( .A(n_398), .Y(n_431) );
OR2x6_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx2_ASAP7_75t_L g476 ( .A(n_401), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_401), .B(n_488), .Y(n_487) );
NAND2xp33_ASAP7_75t_SL g538 ( .A(n_402), .B(n_539), .Y(n_538) );
INVx2_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
OAI32xp33_ASAP7_75t_L g404 ( .A1(n_403), .A2(n_405), .A3(n_409), .B1(n_411), .B2(n_414), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_403), .B(n_506), .Y(n_552) );
OR2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx2_ASAP7_75t_L g515 ( .A(n_407), .Y(n_515) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g486 ( .A(n_413), .B(n_458), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_434), .C(n_452), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_423), .B2(n_426), .Y(n_417) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
O2A1O1Ixp5_ASAP7_75t_L g463 ( .A1(n_422), .A2(n_464), .B(n_465), .C(n_469), .Y(n_463) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_422), .Y(n_521) );
INVx1_ASAP7_75t_L g565 ( .A(n_422), .Y(n_565) );
INVxp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_430), .Y(n_427) );
INVx1_ASAP7_75t_L g532 ( .A(n_428), .Y(n_532) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g537 ( .A(n_429), .B(n_494), .Y(n_537) );
INVx1_ASAP7_75t_L g444 ( .A(n_430), .Y(n_444) );
NOR2x1p5_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g495 ( .A(n_433), .Y(n_495) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_440), .B1(n_443), .B2(n_446), .C(n_451), .Y(n_434) );
INVx1_ASAP7_75t_L g490 ( .A(n_435), .Y(n_490) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g525 ( .A(n_438), .B(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_440), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_450), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g517 ( .A(n_449), .B(n_483), .Y(n_517) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_455), .B1(n_456), .B2(n_459), .C(n_463), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
AND2x4_ASAP7_75t_L g536 ( .A(n_460), .B(n_537), .Y(n_536) );
INVx2_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g535 ( .A(n_461), .B(n_510), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx3_ASAP7_75t_R g539 ( .A(n_468), .Y(n_539) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NOR4xp25_ASAP7_75t_L g472 ( .A(n_473), .B(n_485), .C(n_489), .D(n_504), .Y(n_472) );
OAI21xp33_ASAP7_75t_SL g473 ( .A1(n_474), .A2(n_477), .B(n_479), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AOI21xp33_ASAP7_75t_SL g485 ( .A1(n_477), .A2(n_486), .B(n_487), .Y(n_485) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g566 ( .A1(n_481), .A2(n_517), .B(n_567), .Y(n_566) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI221xp5_ASAP7_75t_SL g489 ( .A1(n_490), .A2(n_491), .B1(n_497), .B2(n_499), .C(n_501), .Y(n_489) );
OAI221xp5_ASAP7_75t_L g504 ( .A1(n_491), .A2(n_505), .B1(n_507), .B2(n_511), .C(n_513), .Y(n_504) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_496), .Y(n_492) );
INVx1_ASAP7_75t_L g531 ( .A(n_493), .Y(n_531) );
AND2x4_ASAP7_75t_L g550 ( .A(n_493), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g547 ( .A(n_494), .Y(n_547) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVxp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND4xp25_ASAP7_75t_L g528 ( .A(n_506), .B(n_529), .C(n_530), .D(n_532), .Y(n_528) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVxp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_517), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
NOR3xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_540), .C(n_559), .Y(n_518) );
NAND4xp25_ASAP7_75t_L g519 ( .A(n_520), .B(n_522), .C(n_528), .D(n_533), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_527), .Y(n_548) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_SL g543 ( .A(n_544), .B(n_548), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_568), .Y(n_571) );
BUFx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx12f_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_574), .Y(n_579) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
INVx3_ASAP7_75t_L g950 ( .A(n_581), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_581), .B(n_956), .Y(n_955) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_944), .B(n_951), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_936), .B1(n_942), .B2(n_943), .Y(n_583) );
INVx2_ASAP7_75t_L g943 ( .A(n_584), .Y(n_943) );
AO21x2_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_588), .B(n_589), .Y(n_584) );
AOI31xp33_ASAP7_75t_L g589 ( .A1(n_585), .A2(n_590), .A3(n_824), .B(n_899), .Y(n_589) );
INVxp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
BUFx6f_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
NOR2x1_ASAP7_75t_L g590 ( .A(n_591), .B(n_771), .Y(n_590) );
NAND3xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_741), .C(n_761), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_635), .B1(n_695), .B2(n_704), .C(n_719), .Y(n_592) );
INVxp67_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_625), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_613), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g794 ( .A(n_597), .Y(n_794) );
AND2x2_ASAP7_75t_L g848 ( .A(n_597), .B(n_840), .Y(n_848) );
AND2x2_ASAP7_75t_L g929 ( .A(n_597), .B(n_627), .Y(n_929) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_598), .B(n_706), .Y(n_737) );
AND2x2_ASAP7_75t_L g871 ( .A(n_598), .B(n_627), .Y(n_871) );
INVx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g718 ( .A(n_599), .B(n_614), .Y(n_718) );
AND2x2_ASAP7_75t_L g722 ( .A(n_599), .B(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g750 ( .A(n_599), .B(n_627), .Y(n_750) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_599), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_599), .B(n_614), .Y(n_805) );
AND2x4_ASAP7_75t_L g599 ( .A(n_600), .B(n_603), .Y(n_599) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_608), .B(n_612), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B(n_607), .Y(n_604) );
OAI21xp5_ASAP7_75t_L g673 ( .A1(n_607), .A2(n_674), .B(n_677), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_611), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_611), .A2(n_710), .B(n_711), .Y(n_709) );
OR2x2_ASAP7_75t_L g770 ( .A(n_613), .B(n_725), .Y(n_770) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g723 ( .A(n_614), .Y(n_723) );
INVx1_ASAP7_75t_L g735 ( .A(n_614), .Y(n_735) );
INVx1_ASAP7_75t_L g760 ( .A(n_614), .Y(n_760) );
AND2x2_ASAP7_75t_L g818 ( .A(n_614), .B(n_707), .Y(n_818) );
OAI21xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_620), .B(n_623), .Y(n_615) );
AND2x4_ASAP7_75t_L g640 ( .A(n_623), .B(n_641), .Y(n_640) );
AOI21xp33_ASAP7_75t_L g693 ( .A1(n_623), .A2(n_692), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g779 ( .A(n_625), .Y(n_779) );
OR2x2_ASAP7_75t_L g808 ( .A(n_625), .B(n_770), .Y(n_808) );
OR2x2_ASAP7_75t_L g827 ( .A(n_625), .B(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g789 ( .A(n_626), .Y(n_789) );
AND2x2_ASAP7_75t_L g836 ( .A(n_626), .B(n_727), .Y(n_836) );
HB1xp67_ASAP7_75t_L g906 ( .A(n_626), .Y(n_906) );
BUFx3_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g705 ( .A(n_627), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g724 ( .A(n_627), .B(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g792 ( .A(n_627), .B(n_723), .Y(n_792) );
INVx2_ASAP7_75t_SL g840 ( .A(n_627), .Y(n_840) );
AO31x2_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .A3(n_632), .B(n_633), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_631), .B(n_671), .Y(n_670) );
INVxp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_662), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_637), .B(n_776), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_637), .A2(n_811), .B1(n_818), .B2(n_819), .Y(n_817) );
AND2x2_ASAP7_75t_L g902 ( .A(n_637), .B(n_903), .Y(n_902) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_652), .Y(n_637) );
INVx2_ASAP7_75t_L g699 ( .A(n_638), .Y(n_699) );
INVx1_ASAP7_75t_L g754 ( .A(n_638), .Y(n_754) );
OR2x2_ASAP7_75t_L g765 ( .A(n_638), .B(n_681), .Y(n_765) );
AND2x2_ASAP7_75t_L g860 ( .A(n_638), .B(n_653), .Y(n_860) );
NAND2x1p5_ASAP7_75t_L g638 ( .A(n_639), .B(n_647), .Y(n_638) );
NAND2x1_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
AOI21x1_ASAP7_75t_L g647 ( .A1(n_640), .A2(n_648), .B(n_651), .Y(n_647) );
O2A1O1Ixp5_ASAP7_75t_L g708 ( .A1(n_640), .A2(n_709), .B(n_712), .C(n_715), .Y(n_708) );
INVx2_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g731 ( .A(n_652), .Y(n_731) );
INVx1_ASAP7_75t_L g745 ( .A(n_652), .Y(n_745) );
INVx1_ASAP7_75t_L g755 ( .A(n_652), .Y(n_755) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVxp33_ASAP7_75t_L g843 ( .A(n_653), .Y(n_843) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_662), .Y(n_773) );
INVx1_ASAP7_75t_L g872 ( .A(n_662), .Y(n_872) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g859 ( .A(n_664), .B(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g886 ( .A(n_664), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_680), .Y(n_664) );
INVx3_ASAP7_75t_L g703 ( .A(n_665), .Y(n_703) );
AND2x2_ASAP7_75t_L g785 ( .A(n_665), .B(n_731), .Y(n_785) );
AO21x2_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_668), .B(n_672), .Y(n_665) );
AO21x1_ASAP7_75t_SL g728 ( .A1(n_666), .A2(n_668), .B(n_672), .Y(n_728) );
INVxp67_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
OAI21x1_ASAP7_75t_SL g672 ( .A1(n_667), .A2(n_673), .B(n_679), .Y(n_672) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_L g683 ( .A(n_676), .Y(n_683) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g700 ( .A(n_681), .Y(n_700) );
INVx2_ASAP7_75t_L g730 ( .A(n_681), .Y(n_730) );
AND2x2_ASAP7_75t_L g740 ( .A(n_681), .B(n_699), .Y(n_740) );
AND2x2_ASAP7_75t_L g776 ( .A(n_681), .B(n_703), .Y(n_776) );
AND2x2_ASAP7_75t_L g856 ( .A(n_681), .B(n_698), .Y(n_856) );
AO21x2_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_687), .B(n_693), .Y(n_681) );
NOR2xp67_ASAP7_75t_L g684 ( .A(n_683), .B(n_685), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_691), .B(n_692), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_694), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OR2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_701), .Y(n_696) );
OR2x2_ASAP7_75t_L g924 ( .A(n_697), .B(n_745), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .Y(n_697) );
OR2x2_ASAP7_75t_L g802 ( .A(n_698), .B(n_731), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_698), .B(n_702), .Y(n_933) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g809 ( .A(n_701), .Y(n_809) );
BUFx2_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g747 ( .A(n_702), .Y(n_747) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g842 ( .A(n_703), .B(n_843), .Y(n_842) );
AND2x2_ASAP7_75t_L g849 ( .A(n_703), .B(n_730), .Y(n_849) );
OR2x2_ASAP7_75t_L g865 ( .A(n_703), .B(n_730), .Y(n_865) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_717), .Y(n_704) );
AND2x4_ASAP7_75t_L g804 ( .A(n_705), .B(n_805), .Y(n_804) );
AND2x4_ASAP7_75t_L g823 ( .A(n_705), .B(n_722), .Y(n_823) );
INVx2_ASAP7_75t_L g725 ( .A(n_706), .Y(n_725) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g749 ( .A(n_707), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_707), .B(n_760), .Y(n_759) );
BUFx2_ASAP7_75t_SL g781 ( .A(n_707), .Y(n_781) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g837 ( .A(n_717), .Y(n_837) );
BUFx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g780 ( .A(n_718), .B(n_781), .Y(n_780) );
AND2x4_ASAP7_75t_SL g854 ( .A(n_718), .B(n_840), .Y(n_854) );
AND2x2_ASAP7_75t_L g915 ( .A(n_718), .B(n_749), .Y(n_915) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_726), .B1(n_732), .B2(n_738), .Y(n_719) );
INVx3_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AND2x4_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
NAND3xp33_ASAP7_75t_L g894 ( .A(n_725), .B(n_895), .C(n_896), .Y(n_894) );
INVx1_ASAP7_75t_L g928 ( .A(n_725), .Y(n_928) );
OR2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
AND2x2_ASAP7_75t_L g739 ( .A(n_727), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g762 ( .A(n_727), .B(n_763), .Y(n_762) );
AND2x4_ASAP7_75t_SL g821 ( .A(n_727), .B(n_813), .Y(n_821) );
INVx5_ASAP7_75t_L g875 ( .A(n_727), .Y(n_875) );
AND2x4_ASAP7_75t_L g914 ( .A(n_727), .B(n_856), .Y(n_914) );
AND2x2_ASAP7_75t_L g918 ( .A(n_727), .B(n_801), .Y(n_918) );
BUFx6f_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVxp67_ASAP7_75t_L g903 ( .A(n_728), .Y(n_903) );
NOR2x1_ASAP7_75t_L g932 ( .A(n_729), .B(n_933), .Y(n_932) );
OR2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g797 ( .A(n_730), .Y(n_797) );
NAND2xp5_ASAP7_75t_SL g893 ( .A(n_732), .B(n_894), .Y(n_893) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AND2x4_ASAP7_75t_L g905 ( .A(n_733), .B(n_906), .Y(n_905) );
AND2x4_ASAP7_75t_L g733 ( .A(n_734), .B(n_736), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_735), .B(n_840), .Y(n_839) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OR2x2_ASAP7_75t_L g838 ( .A(n_737), .B(n_839), .Y(n_838) );
OR2x2_ASAP7_75t_L g880 ( .A(n_737), .B(n_792), .Y(n_880) );
INVx2_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
AND2x4_ASAP7_75t_L g746 ( .A(n_740), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g757 ( .A(n_740), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_740), .B(n_785), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_748), .B(n_751), .Y(n_741) );
OAI21xp5_ASAP7_75t_L g922 ( .A1(n_742), .A2(n_923), .B(n_925), .Y(n_922) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2x1_ASAP7_75t_SL g743 ( .A(n_744), .B(n_746), .Y(n_743) );
BUFx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_745), .B(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_745), .B(n_849), .Y(n_878) );
INVx2_ASAP7_75t_L g887 ( .A(n_745), .Y(n_887) );
AND2x4_ASAP7_75t_SL g892 ( .A(n_745), .B(n_834), .Y(n_892) );
NOR2x1_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_749), .B(n_789), .Y(n_788) );
AND2x2_ASAP7_75t_L g812 ( .A(n_749), .B(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g819 ( .A(n_749), .Y(n_819) );
OR2x2_ASAP7_75t_L g758 ( .A(n_750), .B(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g813 ( .A(n_750), .Y(n_813) );
INVx1_ASAP7_75t_L g890 ( .A(n_750), .Y(n_890) );
AOI21xp33_ASAP7_75t_SL g751 ( .A1(n_752), .A2(n_756), .B(n_758), .Y(n_751) );
AOI32xp33_ASAP7_75t_L g881 ( .A1(n_752), .A2(n_849), .A3(n_882), .B1(n_883), .B2(n_888), .Y(n_881) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
INVx3_ASAP7_75t_L g811 ( .A(n_754), .Y(n_811) );
OR2x2_ASAP7_75t_L g764 ( .A(n_755), .B(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g852 ( .A(n_755), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_756), .A2(n_817), .B1(n_820), .B2(n_822), .Y(n_816) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NAND2xp33_ASAP7_75t_L g879 ( .A(n_758), .B(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g795 ( .A(n_759), .Y(n_795) );
BUFx2_ASAP7_75t_L g868 ( .A(n_759), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_766), .Y(n_761) );
AOI221xp5_ASAP7_75t_L g825 ( .A1(n_763), .A2(n_797), .B1(n_826), .B2(n_829), .C(n_832), .Y(n_825) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g801 ( .A(n_765), .Y(n_801) );
INVx1_ASAP7_75t_L g834 ( .A(n_765), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_767), .B(n_831), .Y(n_830) );
AND2x2_ASAP7_75t_L g873 ( .A(n_767), .B(n_795), .Y(n_873) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OR2x6_ASAP7_75t_L g919 ( .A(n_770), .B(n_920), .Y(n_919) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_782), .C(n_806), .Y(n_771) );
OAI21xp33_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_774), .B(n_777), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
OAI22xp33_ASAP7_75t_L g907 ( .A1(n_775), .A2(n_808), .B1(n_908), .B2(n_909), .Y(n_907) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
INVx2_ASAP7_75t_L g921 ( .A(n_780), .Y(n_921) );
OR2x2_ASAP7_75t_L g791 ( .A(n_781), .B(n_792), .Y(n_791) );
NOR2x1_ASAP7_75t_SL g831 ( .A(n_781), .B(n_792), .Y(n_831) );
AOI221xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_786), .B1(n_790), .B2(n_796), .C(n_798), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
AND2x2_ASAP7_75t_L g796 ( .A(n_785), .B(n_797), .Y(n_796) );
INVxp67_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
OR2x2_ASAP7_75t_L g935 ( .A(n_788), .B(n_794), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
INVx1_ASAP7_75t_L g896 ( .A(n_794), .Y(n_896) );
AND2x2_ASAP7_75t_L g847 ( .A(n_795), .B(n_848), .Y(n_847) );
AND2x2_ASAP7_75t_L g882 ( .A(n_795), .B(n_871), .Y(n_882) );
AOI21xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_802), .B(n_803), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_799), .A2(n_917), .B1(n_919), .B2(n_921), .Y(n_916) );
BUFx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_800), .B(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g876 ( .A(n_802), .Y(n_876) );
OR2x2_ASAP7_75t_L g908 ( .A(n_802), .B(n_875), .Y(n_908) );
INVx4_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
AOI321xp33_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_809), .A3(n_810), .B1(n_812), .B2(n_814), .C(n_816), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx2_ASAP7_75t_SL g828 ( .A(n_818), .Y(n_828) );
AND2x4_ASAP7_75t_L g870 ( .A(n_818), .B(n_871), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_818), .B(n_890), .Y(n_889) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx4_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
AND5x1_ASAP7_75t_L g824 ( .A(n_825), .B(n_844), .C(n_869), .D(n_881), .E(n_891), .Y(n_824) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
OAI22xp33_ASAP7_75t_L g857 ( .A1(n_827), .A2(n_858), .B1(n_861), .B2(n_866), .Y(n_857) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
OAI32xp33_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_835), .A3(n_837), .B1(n_838), .B2(n_841), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g912 ( .A(n_842), .Y(n_912) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_845), .B(n_857), .Y(n_844) );
OAI32xp33_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_849), .A3(n_850), .B1(n_853), .B2(n_855), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g920 ( .A(n_848), .Y(n_920) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
A2O1A1Ixp33_ASAP7_75t_L g911 ( .A1(n_853), .A2(n_865), .B(n_912), .C(n_913), .Y(n_911) );
INVx2_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVxp33_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_856), .B(n_887), .Y(n_898) );
AND2x2_ASAP7_75t_L g904 ( .A(n_856), .B(n_875), .Y(n_904) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx4_ASAP7_75t_L g863 ( .A(n_860), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_864), .Y(n_861) );
AOI322xp5_ASAP7_75t_L g869 ( .A1(n_862), .A2(n_870), .A3(n_872), .B1(n_873), .B2(n_874), .C1(n_877), .C2(n_879), .Y(n_869) );
INVx6_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVxp67_ASAP7_75t_L g909 ( .A(n_870), .Y(n_909) );
AND2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
INVx1_ASAP7_75t_L g895 ( .A(n_875), .Y(n_895) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g891 ( .A1(n_882), .A2(n_892), .B1(n_893), .B2(n_897), .Y(n_891) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g931 ( .A(n_884), .Y(n_931) );
OR2x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_887), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
OAI31xp33_ASAP7_75t_L g930 ( .A1(n_892), .A2(n_931), .A3(n_932), .B(n_934), .Y(n_930) );
INVx2_ASAP7_75t_SL g897 ( .A(n_898), .Y(n_897) );
AND4x1_ASAP7_75t_L g899 ( .A(n_900), .B(n_910), .C(n_922), .D(n_930), .Y(n_899) );
O2A1O1Ixp33_ASAP7_75t_SL g900 ( .A1(n_901), .A2(n_904), .B(n_905), .C(n_907), .Y(n_900) );
HB1xp67_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
NOR2xp33_ASAP7_75t_SL g910 ( .A(n_911), .B(n_916), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_914), .B(n_915), .Y(n_913) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .Y(n_927) );
INVx2_ASAP7_75t_SL g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g942 ( .A(n_936), .Y(n_942) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g944 ( .A(n_945), .Y(n_944) );
BUFx8_ASAP7_75t_SL g945 ( .A(n_946), .Y(n_945) );
OR2x6_ASAP7_75t_L g946 ( .A(n_947), .B(n_950), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_948), .B(n_949), .Y(n_947) );
NOR2xp33_ASAP7_75t_L g951 ( .A(n_952), .B(n_953), .Y(n_951) );
BUFx3_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
BUFx3_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
NOR2xp33_ASAP7_75t_L g957 ( .A(n_958), .B(n_959), .Y(n_957) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx4_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
endmodule