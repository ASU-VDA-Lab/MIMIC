module fake_jpeg_15257_n_225 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_225);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_29),
.B(n_19),
.Y(n_47)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_24),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_13),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_29),
.B(n_22),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_25),
.B1(n_21),
.B2(n_22),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_45),
.B1(n_13),
.B2(n_27),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_25),
.B1(n_22),
.B2(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_47),
.B(n_15),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_14),
.Y(n_61)
);

INVxp67_ASAP7_75t_SL g62 ( 
.A(n_54),
.Y(n_62)
);

INVxp67_ASAP7_75t_SL g88 ( 
.A(n_62),
.Y(n_88)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_66),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_65),
.A2(n_17),
.B(n_9),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_15),
.B1(n_19),
.B2(n_21),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_69),
.A2(n_74),
.B1(n_75),
.B2(n_80),
.Y(n_92)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_15),
.B1(n_26),
.B2(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_14),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_79),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_81),
.B(n_26),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_17),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_39),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_39),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_83),
.B(n_85),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_42),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_89),
.A2(n_104),
.B1(n_17),
.B2(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_42),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_91),
.B(n_95),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_66),
.B(n_41),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_26),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_41),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_100),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_45),
.B1(n_54),
.B2(n_37),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_106),
.B1(n_107),
.B2(n_43),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_63),
.B(n_77),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_63),
.B(n_44),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_60),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_59),
.A2(n_50),
.B1(n_43),
.B2(n_31),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_60),
.A2(n_37),
.B1(n_43),
.B2(n_50),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_50),
.B1(n_103),
.B2(n_64),
.Y(n_137)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_112),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_113),
.B(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_67),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_120),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_67),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_123),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_101),
.B(n_89),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_131),
.C(n_7),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_78),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_89),
.A2(n_84),
.B1(n_95),
.B2(n_108),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_126),
.B1(n_122),
.B2(n_115),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_57),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_130),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_0),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_129),
.A2(n_133),
.B(n_23),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_80),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_SL g131 ( 
.A(n_104),
.B(n_74),
.C(n_32),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_134),
.B(n_150),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_99),
.B1(n_84),
.B2(n_106),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_136),
.A2(n_137),
.B1(n_121),
.B2(n_113),
.Y(n_173)
);

NAND2xp33_ASAP7_75t_SL g178 ( 
.A(n_140),
.B(n_23),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_102),
.B1(n_94),
.B2(n_87),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_151),
.B1(n_156),
.B2(n_157),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_124),
.B(n_130),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_120),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_107),
.C(n_93),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_154),
.C(n_109),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_132),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_68),
.B1(n_73),
.B2(n_72),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_93),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_153),
.B(n_36),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_115),
.Y(n_154)
);

AOI221xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_109),
.B1(n_118),
.B2(n_126),
.C(n_131),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_112),
.A2(n_70),
.B1(n_88),
.B2(n_32),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_93),
.B1(n_20),
.B2(n_16),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_152),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_160),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_152),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_117),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_135),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_163),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_142),
.Y(n_163)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_125),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_170),
.C(n_171),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_168),
.B(n_176),
.Y(n_188)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_128),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_174),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_129),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_175),
.A2(n_178),
.B1(n_179),
.B2(n_147),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_134),
.A2(n_129),
.B1(n_20),
.B2(n_16),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_176),
.A2(n_158),
.B1(n_20),
.B2(n_141),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_177),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_158),
.A2(n_148),
.B1(n_136),
.B2(n_150),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_141),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_189),
.C(n_24),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_145),
.C(n_138),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_145),
.C(n_138),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_163),
.C(n_164),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_197),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_168),
.C(n_173),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_200),
.C(n_202),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g197 ( 
.A(n_191),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_192),
.A2(n_175),
.B(n_10),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_184),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_14),
.C(n_24),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_186),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_24),
.C(n_34),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_189),
.C(n_180),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_187),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_206),
.C(n_208),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_190),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_207),
.B(n_210),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_198),
.A2(n_194),
.B(n_193),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_211),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_1),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_212),
.A2(n_214),
.B(n_209),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_217),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_213),
.A2(n_6),
.B(n_12),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_1),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_2),
.B(n_3),
.Y(n_222)
);

NAND2xp33_ASAP7_75t_SL g221 ( 
.A(n_220),
.B(n_5),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_221),
.A2(n_222),
.B(n_2),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_4),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_33),
.C(n_36),
.Y(n_225)
);


endmodule