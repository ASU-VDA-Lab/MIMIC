module fake_jpeg_18004_n_348 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx8_ASAP7_75t_SL g23 ( 
.A(n_4),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_6),
.B(n_12),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2x1_ASAP7_75t_SL g41 ( 
.A(n_24),
.B(n_0),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_26),
.B(n_21),
.Y(n_71)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_18),
.Y(n_65)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_20),
.B1(n_24),
.B2(n_16),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_51),
.A2(n_61),
.B1(n_17),
.B2(n_19),
.Y(n_109)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_20),
.B1(n_27),
.B2(n_30),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_65),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_73),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_71),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_72),
.Y(n_79)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g121 ( 
.A(n_75),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_30),
.B1(n_27),
.B2(n_47),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_76),
.A2(n_28),
.B1(n_21),
.B2(n_32),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_68),
.A2(n_30),
.B1(n_16),
.B2(n_17),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_77),
.A2(n_32),
.B(n_31),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_87),
.Y(n_113)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_53),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_91),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_56),
.A2(n_30),
.B1(n_50),
.B2(n_47),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_94),
.A2(n_25),
.B1(n_21),
.B2(n_32),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_37),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_97),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_31),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_55),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_98),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_58),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_100),
.Y(n_128)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_103),
.Y(n_137)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_34),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_106),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_34),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_16),
.B(n_25),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_49),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_49),
.B1(n_44),
.B2(n_28),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_122),
.B1(n_127),
.B2(n_131),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_41),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_129),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_79),
.B1(n_86),
.B2(n_78),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_94),
.B1(n_98),
.B2(n_100),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_41),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_28),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_76),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_81),
.C(n_84),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_129),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_141),
.A2(n_19),
.B1(n_35),
.B2(n_79),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_17),
.B1(n_19),
.B2(n_35),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_111),
.B(n_85),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_149),
.B(n_161),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_144),
.B(n_150),
.Y(n_178)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_147),
.A2(n_121),
.B1(n_117),
.B2(n_104),
.Y(n_187)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_148),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_31),
.B(n_25),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_138),
.Y(n_152)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_102),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_153),
.B(n_155),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_93),
.B1(n_89),
.B2(n_82),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_154),
.A2(n_156),
.B1(n_23),
.B2(n_22),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_84),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_93),
.B1(n_96),
.B2(n_92),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_157),
.A2(n_166),
.B1(n_121),
.B2(n_119),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_125),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_158),
.B(n_159),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_160),
.B(n_167),
.Y(n_208)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_124),
.B(n_87),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_SL g162 ( 
.A1(n_124),
.A2(n_96),
.B(n_79),
.C(n_99),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_139),
.B(n_114),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_170),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_165),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_116),
.A2(n_123),
.B1(n_132),
.B2(n_112),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_116),
.B(n_29),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_0),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_22),
.B(n_29),
.Y(n_206)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_169),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_78),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_135),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_173),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_88),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_174),
.Y(n_209)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_139),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_182),
.A2(n_189),
.B(n_194),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_192),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_142),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_184),
.A2(n_200),
.B1(n_201),
.B2(n_206),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_187),
.A2(n_191),
.B1(n_146),
.B2(n_165),
.Y(n_236)
);

AND2x6_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_128),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g232 ( 
.A1(n_190),
.A2(n_168),
.A3(n_167),
.B1(n_157),
.B2(n_170),
.C1(n_162),
.C2(n_175),
.Y(n_232)
);

AO22x2_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_106),
.B1(n_103),
.B2(n_75),
.Y(n_191)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

AND2x4_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_121),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_151),
.A2(n_101),
.B1(n_115),
.B2(n_118),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_196),
.B1(n_172),
.B2(n_152),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_150),
.A2(n_115),
.B1(n_137),
.B2(n_35),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_145),
.B(n_29),
.C(n_36),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_203),
.C(n_209),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_162),
.A2(n_1),
.B(n_2),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_203),
.B(n_205),
.Y(n_213)
);

OAI22x1_ASAP7_75t_SL g200 ( 
.A1(n_162),
.A2(n_36),
.B1(n_23),
.B2(n_135),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_168),
.A2(n_23),
.B1(n_22),
.B2(n_29),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_162),
.A2(n_1),
.B(n_2),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_182),
.A2(n_143),
.B1(n_173),
.B2(n_147),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_230),
.B1(n_234),
.B2(n_236),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_212),
.B(n_219),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_204),
.B(n_145),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_217),
.C(n_226),
.Y(n_243)
);

A2O1A1O1Ixp25_ASAP7_75t_L g215 ( 
.A1(n_180),
.A2(n_184),
.B(n_194),
.C(n_190),
.D(n_206),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_192),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_166),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_218),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_188),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_222),
.Y(n_258)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_155),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_225),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_224),
.A2(n_228),
.B1(n_237),
.B2(n_29),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_153),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_159),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_191),
.A2(n_194),
.B1(n_199),
.B2(n_205),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_227),
.A2(n_186),
.B1(n_189),
.B2(n_195),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_176),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_198),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_229),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_191),
.A2(n_200),
.B1(n_194),
.B2(n_209),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_225),
.B(n_223),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_226),
.C(n_217),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_191),
.A2(n_158),
.B1(n_144),
.B2(n_174),
.Y(n_234)
);

AOI22x1_ASAP7_75t_L g237 ( 
.A1(n_191),
.A2(n_163),
.B1(n_164),
.B2(n_156),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_189),
.A2(n_171),
.B1(n_163),
.B2(n_22),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_238),
.A2(n_183),
.B(n_198),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_240),
.B(n_235),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_242),
.A2(n_244),
.B1(n_246),
.B2(n_253),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_207),
.B1(n_208),
.B2(n_187),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_247),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_176),
.C(n_202),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g264 ( 
.A(n_250),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_216),
.A2(n_187),
.B1(n_207),
.B2(n_179),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_251),
.A2(n_257),
.B1(n_210),
.B2(n_221),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_224),
.B1(n_231),
.B2(n_233),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_177),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_263),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_187),
.B1(n_179),
.B2(n_196),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_213),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_215),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_236),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_234),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_228),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_260),
.Y(n_269)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_213),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_212),
.Y(n_267)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_267),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_270),
.B(n_275),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_235),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_280),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_218),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_277),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_243),
.B(n_238),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_262),
.B(n_210),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_276),
.B(n_278),
.Y(n_288)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_249),
.A2(n_222),
.B1(n_220),
.B2(n_9),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_279),
.A2(n_260),
.B1(n_263),
.B2(n_259),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_22),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_243),
.B(n_22),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_282),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_240),
.B(n_29),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_283),
.A2(n_284),
.B(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_241),
.Y(n_284)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_285),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_242),
.B(n_253),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_286),
.A2(n_275),
.B(n_281),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_273),
.B1(n_269),
.B2(n_270),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_287),
.A2(n_13),
.B1(n_14),
.B2(n_286),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_247),
.C(n_246),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_291),
.C(n_293),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_266),
.B(n_262),
.CI(n_244),
.CON(n_290),
.SN(n_290)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_290),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_256),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_255),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_294),
.Y(n_303)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_248),
.C(n_29),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_7),
.C(n_8),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_264),
.Y(n_304)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_304),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_308),
.C(n_295),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_297),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_299),
.Y(n_324)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_307),
.Y(n_323)
);

XNOR2x1_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_9),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_10),
.Y(n_311)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_311),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_10),
.C(n_11),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_313),
.B(n_314),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_11),
.C(n_12),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_12),
.C(n_13),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_315),
.B(n_316),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_319),
.A2(n_308),
.B1(n_305),
.B2(n_312),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_293),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_302),
.C(n_292),
.Y(n_332)
);

OR2x2_ASAP7_75t_SL g322 ( 
.A(n_303),
.B(n_290),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_316),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_324),
.B(n_325),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_310),
.B(n_296),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_309),
.A2(n_287),
.B(n_290),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_313),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_328),
.A2(n_329),
.B(n_321),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_330),
.A2(n_332),
.B(n_315),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_311),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_333),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_322),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_317),
.B(n_314),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_334),
.B(n_318),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_337),
.B(n_338),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_323),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_339),
.B(n_340),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_335),
.C(n_320),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_343),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_341),
.C(n_336),
.Y(n_345)
);

OAI311xp33_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_324),
.A3(n_319),
.B1(n_306),
.C1(n_307),
.Y(n_346)
);

AOI21x1_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_294),
.B(n_301),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_347),
.A2(n_298),
.B(n_14),
.Y(n_348)
);


endmodule