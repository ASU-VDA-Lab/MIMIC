module fake_jpeg_31154_n_33 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_33);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_33;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_31;
wire n_25;
wire n_17;
wire n_29;
wire n_32;
wire n_15;

INVx5_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_1),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_18),
.A2(n_12),
.B1(n_10),
.B2(n_6),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_19),
.A2(n_21),
.B1(n_15),
.B2(n_14),
.Y(n_28)
);

CKINVDCx12_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_20),
.B(n_22),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_3),
.C(n_4),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_3),
.C(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_20),
.Y(n_26)
);

NOR3xp33_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_28),
.C(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_30),
.Y(n_31)
);

AOI322xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_25),
.A3(n_30),
.B1(n_28),
.B2(n_24),
.C1(n_17),
.C2(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_32),
.B(n_17),
.Y(n_33)
);


endmodule