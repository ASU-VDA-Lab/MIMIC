module fake_jpeg_31795_n_264 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_33),
.Y(n_52)
);

NAND3xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_14),
.C(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_41),
.Y(n_55)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_43),
.Y(n_59)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_47),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_18),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_19),
.B1(n_27),
.B2(n_24),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_62),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_23),
.B1(n_17),
.B2(n_16),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_57),
.B1(n_16),
.B2(n_45),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_27),
.B1(n_24),
.B2(n_30),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_39),
.B1(n_30),
.B2(n_22),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_23),
.B1(n_17),
.B2(n_16),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_32),
.B(n_22),
.C(n_21),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_61),
.B(n_42),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_24),
.B1(n_27),
.B2(n_16),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_47),
.B1(n_43),
.B2(n_33),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_67),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_62),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_34),
.A3(n_48),
.B1(n_46),
.B2(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_75),
.Y(n_102)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_52),
.B1(n_32),
.B2(n_22),
.Y(n_110)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_60),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_31),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_79),
.Y(n_112)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_26),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_89),
.C(n_29),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_88),
.B1(n_53),
.B2(n_84),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_39),
.B1(n_33),
.B2(n_30),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_52),
.B1(n_35),
.B2(n_41),
.Y(n_93)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_31),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_86),
.B(n_29),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_61),
.B(n_36),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_61),
.C(n_57),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_32),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_90),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_92),
.A2(n_49),
.B(n_16),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_52),
.B(n_74),
.C(n_41),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_109),
.Y(n_123)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_107),
.B(n_11),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_53),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_106),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_84),
.A2(n_63),
.B1(n_49),
.B2(n_47),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_113),
.A2(n_88),
.B1(n_78),
.B2(n_65),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_100),
.B1(n_60),
.B2(n_85),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_84),
.B1(n_67),
.B2(n_70),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_115),
.A2(n_119),
.B1(n_122),
.B2(n_60),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_80),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_133),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_95),
.B1(n_113),
.B2(n_105),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_77),
.B1(n_79),
.B2(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_106),
.B(n_86),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_127),
.C(n_131),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_75),
.B1(n_76),
.B2(n_69),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_89),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_102),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_21),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_90),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_74),
.B(n_52),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_95),
.B(n_52),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_101),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_97),
.B(n_94),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_63),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_105),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_136),
.A2(n_144),
.B(n_145),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_141),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_128),
.C(n_122),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_143),
.C(n_134),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_97),
.C(n_109),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_132),
.A2(n_100),
.B(n_101),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_156),
.Y(n_167)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_100),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_152),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_151),
.A2(n_125),
.B1(n_116),
.B2(n_91),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_98),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_154),
.B(n_114),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_119),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_126),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_103),
.B(n_73),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_121),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_159),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_115),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_160),
.B(n_177),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_151),
.B1(n_156),
.B2(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_171),
.B1(n_178),
.B2(n_174),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_174),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_126),
.B1(n_118),
.B2(n_131),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_169),
.A2(n_91),
.B1(n_60),
.B2(n_54),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_150),
.C(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_153),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_136),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_118),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_118),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_176),
.C(n_178),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_116),
.C(n_58),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_108),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_118),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_147),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_179),
.B(n_25),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_182),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_146),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_191),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_167),
.A2(n_145),
.B(n_148),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_187),
.A2(n_192),
.B(n_45),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_188),
.B(n_162),
.Y(n_207)
);

OAI22x1_ASAP7_75t_L g190 ( 
.A1(n_173),
.A2(n_149),
.B1(n_146),
.B2(n_137),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_197),
.B1(n_169),
.B2(n_181),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_137),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_167),
.A2(n_108),
.B(n_36),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_54),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_196),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_198),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_162),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_206),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_168),
.C(n_175),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_208),
.C(n_180),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_173),
.C(n_108),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_211),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_190),
.A2(n_45),
.B(n_41),
.Y(n_211)
);

AO22x1_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_35),
.B1(n_25),
.B2(n_3),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_213),
.A2(n_189),
.B1(n_196),
.B2(n_35),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_186),
.B1(n_185),
.B2(n_205),
.Y(n_214)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_200),
.B(n_195),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_219),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_184),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_217),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_197),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_192),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_220),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_212),
.B(n_180),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_193),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g227 ( 
.A(n_222),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_232),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_203),
.Y(n_228)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_225),
.A2(n_213),
.B1(n_199),
.B2(n_211),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_220),
.B(n_203),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_221),
.B(n_216),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_24),
.B1(n_17),
.B2(n_23),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_189),
.Y(n_235)
);

OAI21x1_ASAP7_75t_L g237 ( 
.A1(n_235),
.A2(n_201),
.B(n_223),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_230),
.A2(n_213),
.B1(n_217),
.B2(n_210),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_237),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_221),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_241),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_239),
.B(n_240),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_231),
.A2(n_10),
.B(n_14),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_238),
.A2(n_231),
.B(n_226),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_244),
.B(n_9),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_249),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_243),
.B(n_226),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_8),
.C(n_13),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_5),
.C(n_6),
.Y(n_254)
);

AOI322xp5_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_8),
.A3(n_13),
.B1(n_12),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_253),
.B1(n_245),
.B2(n_2),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_252),
.B(n_254),
.Y(n_259)
);

AOI322xp5_ASAP7_75t_L g253 ( 
.A1(n_247),
.A2(n_10),
.A3(n_13),
.B1(n_12),
.B2(n_5),
.C1(n_6),
.C2(n_11),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_257),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_248),
.C(n_25),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

NAND2xp33_ASAP7_75t_SL g261 ( 
.A(n_258),
.B(n_0),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_259),
.B(n_2),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_262),
.A2(n_263),
.B1(n_3),
.B2(n_25),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_260),
.A2(n_0),
.B(n_2),
.Y(n_263)
);


endmodule