module fake_jpeg_29204_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_31),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_2),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_42),
.Y(n_62)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_3),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_3),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_22),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_24),
.B(n_4),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_51),
.Y(n_58)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_29),
.B1(n_26),
.B2(n_20),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_72),
.B1(n_77),
.B2(n_43),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_18),
.B1(n_16),
.B2(n_20),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_55),
.A2(n_45),
.B1(n_51),
.B2(n_21),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_63),
.Y(n_99)
);

OR2x6_ASAP7_75t_SL g65 ( 
.A(n_36),
.B(n_31),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_66),
.B(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_32),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_32),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_37),
.A2(n_28),
.B(n_23),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_43),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_4),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_23),
.B1(n_22),
.B2(n_18),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_16),
.B1(n_5),
.B2(n_7),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_21),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_37),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_106),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_85),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_98),
.Y(n_123)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_40),
.B1(n_53),
.B2(n_35),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_92),
.B1(n_94),
.B2(n_54),
.Y(n_117)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_50),
.B1(n_47),
.B2(n_51),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_51),
.B1(n_45),
.B2(n_41),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_45),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_70),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_102),
.Y(n_124)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_56),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_62),
.B(n_4),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_105),
.B(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_5),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_57),
.B(n_5),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_77),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_106),
.B(n_90),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_110),
.B(n_99),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_126),
.C(n_10),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_122),
.B1(n_100),
.B2(n_97),
.Y(n_134)
);

FAx1_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_64),
.CI(n_73),
.CON(n_118),
.SN(n_118)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_120),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_74),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_85),
.A2(n_74),
.B1(n_64),
.B2(n_78),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_80),
.C(n_9),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_81),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_91),
.Y(n_144)
);

OAI22x1_ASAP7_75t_SL g129 ( 
.A1(n_86),
.A2(n_100),
.B1(n_87),
.B2(n_89),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_131),
.B1(n_104),
.B2(n_56),
.Y(n_142)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_118),
.B(n_120),
.C(n_115),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_149),
.B(n_132),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_134),
.A2(n_144),
.B1(n_111),
.B2(n_121),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_135),
.B(n_136),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_87),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_110),
.B(n_8),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_141),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_118),
.B1(n_127),
.B2(n_114),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_142),
.B1(n_147),
.B2(n_122),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_92),
.B1(n_104),
.B2(n_108),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_140),
.A2(n_145),
.B1(n_142),
.B2(n_117),
.Y(n_152)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_143),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_78),
.B1(n_103),
.B2(n_88),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_128),
.Y(n_146)
);

BUFx4f_ASAP7_75t_SL g151 ( 
.A(n_146),
.Y(n_151)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_112),
.C(n_121),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_98),
.B(n_11),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_152),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_SL g155 ( 
.A1(n_137),
.A2(n_113),
.A3(n_126),
.B1(n_112),
.B2(n_116),
.C1(n_131),
.C2(n_123),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_160),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_159),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_119),
.C(n_128),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_11),
.C(n_12),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_12),
.C(n_144),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_161),
.A2(n_158),
.B(n_154),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_132),
.B1(n_145),
.B2(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_162),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_163),
.A2(n_147),
.B(n_164),
.C(n_160),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_148),
.B1(n_135),
.B2(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_163),
.A2(n_149),
.B1(n_146),
.B2(n_141),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_151),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_157),
.Y(n_172)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_159),
.B(n_152),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_175),
.B(n_161),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_180),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_177),
.B(n_179),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_153),
.C(n_151),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_167),
.B(n_175),
.Y(n_182)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

OA21x2_ASAP7_75t_SL g183 ( 
.A1(n_169),
.A2(n_173),
.B(n_174),
.Y(n_183)
);

BUFx24_ASAP7_75t_SL g189 ( 
.A(n_183),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_181),
.A2(n_171),
.B(n_180),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_179),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_176),
.A2(n_166),
.B1(n_165),
.B2(n_168),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_176),
.Y(n_193)
);

NOR2xp67_ASAP7_75t_SL g190 ( 
.A(n_189),
.B(n_182),
.Y(n_190)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_187),
.A2(n_184),
.B(n_188),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_192),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_194),
.C(n_173),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_177),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_178),
.B(n_166),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_199),
.B(n_197),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_195),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_194),
.B(n_174),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_174),
.Y(n_202)
);


endmodule