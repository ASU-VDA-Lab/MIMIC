module real_aes_1741_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_0), .B(n_148), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_1), .A2(n_156), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_2), .B(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_3), .B(n_148), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_4), .B(n_175), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_5), .B(n_175), .Y(n_509) );
INVx1_ASAP7_75t_L g144 ( .A(n_6), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_7), .B(n_175), .Y(n_538) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_8), .Y(n_112) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_9), .A2(n_463), .B1(n_758), .B2(n_762), .Y(n_757) );
NAND2xp33_ASAP7_75t_L g579 ( .A(n_10), .B(n_173), .Y(n_579) );
AND2x2_ASAP7_75t_L g178 ( .A(n_11), .B(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g189 ( .A(n_12), .B(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g135 ( .A(n_13), .Y(n_135) );
AOI221x1_ASAP7_75t_L g484 ( .A1(n_14), .A2(n_26), .B1(n_148), .B2(n_156), .C(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_15), .B(n_175), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_16), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_17), .B(n_148), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_18), .A2(n_89), .B1(n_466), .B2(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_18), .Y(n_466) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_19), .A2(n_190), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_20), .B(n_133), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_21), .B(n_175), .Y(n_562) );
AO21x1_ASAP7_75t_L g504 ( .A1(n_22), .A2(n_148), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_23), .B(n_148), .Y(n_229) );
INVx1_ASAP7_75t_L g116 ( .A(n_24), .Y(n_116) );
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_25), .A2(n_93), .B1(n_139), .B2(n_148), .Y(n_138) );
NAND2x1_ASAP7_75t_L g496 ( .A(n_27), .B(n_175), .Y(n_496) );
NAND2x1_ASAP7_75t_L g537 ( .A(n_28), .B(n_173), .Y(n_537) );
OR2x2_ASAP7_75t_L g136 ( .A(n_29), .B(n_90), .Y(n_136) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_29), .A2(n_90), .B(n_135), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_30), .B(n_173), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_31), .B(n_175), .Y(n_578) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_32), .A2(n_179), .B(n_240), .Y(n_239) );
INVxp33_ASAP7_75t_L g771 ( .A(n_33), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_34), .B(n_173), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_35), .A2(n_156), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_36), .B(n_175), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_37), .A2(n_156), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g146 ( .A(n_38), .B(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g154 ( .A(n_38), .B(n_144), .Y(n_154) );
INVx1_ASAP7_75t_L g160 ( .A(n_38), .Y(n_160) );
NOR3xp33_ASAP7_75t_L g110 ( .A(n_39), .B(n_111), .C(n_113), .Y(n_110) );
OR2x6_ASAP7_75t_L g454 ( .A(n_39), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_40), .B(n_148), .Y(n_519) );
OAI22xp5_ASAP7_75t_SL g441 ( .A1(n_41), .A2(n_442), .B1(n_443), .B2(n_446), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_41), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_42), .B(n_148), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_43), .B(n_175), .Y(n_214) );
XNOR2xp5_ASAP7_75t_L g464 ( .A(n_44), .B(n_465), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_45), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_46), .B(n_173), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_47), .B(n_148), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_48), .A2(n_156), .B(n_171), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_49), .A2(n_63), .B1(n_444), .B2(n_445), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_49), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_50), .A2(n_156), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_51), .B(n_173), .Y(n_201) );
XNOR2xp5_ASAP7_75t_L g463 ( .A(n_52), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_53), .B(n_173), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_54), .B(n_148), .Y(n_241) );
INVx1_ASAP7_75t_L g142 ( .A(n_55), .Y(n_142) );
INVx1_ASAP7_75t_L g151 ( .A(n_55), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_56), .B(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g209 ( .A(n_57), .B(n_133), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_58), .B(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_59), .B(n_175), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_60), .B(n_173), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_61), .A2(n_156), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_62), .B(n_148), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_63), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_64), .B(n_148), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_65), .B(n_458), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_66), .A2(n_156), .B(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g235 ( .A(n_67), .B(n_134), .Y(n_235) );
AO21x1_ASAP7_75t_L g506 ( .A1(n_68), .A2(n_156), .B(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_69), .B(n_148), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_70), .B(n_173), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_71), .B(n_148), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_72), .B(n_173), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g155 ( .A1(n_73), .A2(n_97), .B1(n_156), .B2(n_158), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_74), .B(n_175), .Y(n_232) );
AND2x2_ASAP7_75t_L g520 ( .A(n_75), .B(n_134), .Y(n_520) );
INVx1_ASAP7_75t_L g147 ( .A(n_76), .Y(n_147) );
INVx1_ASAP7_75t_L g153 ( .A(n_76), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g119 ( .A1(n_77), .A2(n_120), .B1(n_448), .B2(n_449), .Y(n_119) );
INVxp33_ASAP7_75t_L g449 ( .A(n_77), .Y(n_449) );
AND2x2_ASAP7_75t_L g540 ( .A(n_77), .B(n_179), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_78), .B(n_173), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_79), .A2(n_156), .B(n_213), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_80), .A2(n_156), .B(n_199), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_81), .A2(n_156), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g226 ( .A(n_82), .B(n_134), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g132 ( .A(n_83), .B(n_133), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_84), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g456 ( .A(n_84), .Y(n_456) );
AND2x2_ASAP7_75t_L g525 ( .A(n_85), .B(n_179), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_86), .B(n_148), .Y(n_564) );
AND2x2_ASAP7_75t_L g202 ( .A(n_87), .B(n_190), .Y(n_202) );
AND2x2_ASAP7_75t_L g505 ( .A(n_88), .B(n_216), .Y(n_505) );
INVx1_ASAP7_75t_L g467 ( .A(n_89), .Y(n_467) );
AND2x2_ASAP7_75t_L g499 ( .A(n_91), .B(n_179), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_92), .B(n_173), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_94), .B(n_175), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_95), .B(n_173), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_96), .A2(n_156), .B(n_561), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_98), .A2(n_156), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_99), .B(n_175), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_100), .B(n_175), .Y(n_530) );
BUFx2_ASAP7_75t_L g234 ( .A(n_101), .Y(n_234) );
OA22x2_ASAP7_75t_L g117 ( .A1(n_102), .A2(n_118), .B1(n_460), .B2(n_765), .Y(n_117) );
BUFx2_ASAP7_75t_L g769 ( .A(n_102), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_103), .A2(n_156), .B(n_577), .Y(n_576) );
AOI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_117), .B(n_770), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx8_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
BUFx4f_ASAP7_75t_SL g773 ( .A(n_109), .Y(n_773) );
NAND2xp5_ASAP7_75t_SL g109 ( .A(n_110), .B(n_115), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_114), .B(n_453), .Y(n_452) );
AND2x6_ASAP7_75t_SL g472 ( .A(n_114), .B(n_454), .Y(n_472) );
OR2x6_ASAP7_75t_SL g475 ( .A(n_114), .B(n_453), .Y(n_475) );
OR2x2_ASAP7_75t_L g764 ( .A(n_114), .B(n_454), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_116), .B(n_456), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_450), .B(n_457), .Y(n_118) );
INVx2_ASAP7_75t_L g448 ( .A(n_120), .Y(n_448) );
AOI22x1_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_122), .B1(n_441), .B2(n_447), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_121), .A2(n_469), .B1(n_473), .B2(n_476), .Y(n_468) );
INVx4_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_122), .A2(n_477), .B1(n_759), .B2(n_760), .Y(n_758) );
OR2x6_ASAP7_75t_L g122 ( .A(n_123), .B(n_378), .Y(n_122) );
NAND3xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_294), .C(n_331), .Y(n_123) );
NOR3xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_262), .C(n_277), .Y(n_124) );
OAI221xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_206), .B1(n_236), .B2(n_248), .C(n_249), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g127 ( .A(n_128), .B(n_191), .Y(n_127) );
OAI22xp33_ASAP7_75t_SL g322 ( .A1(n_128), .A2(n_286), .B1(n_323), .B2(n_326), .Y(n_322) );
OR2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_163), .Y(n_128) );
OAI21xp33_ASAP7_75t_SL g332 ( .A1(n_129), .A2(n_333), .B(n_339), .Y(n_332) );
OR2x2_ASAP7_75t_L g361 ( .A(n_129), .B(n_193), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_129), .B(n_281), .Y(n_362) );
INVx2_ASAP7_75t_L g393 ( .A(n_129), .Y(n_393) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_130), .B(n_253), .Y(n_374) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OR2x2_ASAP7_75t_L g248 ( .A(n_131), .B(n_166), .Y(n_248) );
BUFx3_ASAP7_75t_L g274 ( .A(n_131), .Y(n_274) );
AND2x2_ASAP7_75t_L g410 ( .A(n_131), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g433 ( .A(n_131), .B(n_194), .Y(n_433) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_137), .Y(n_131) );
AND2x4_ASAP7_75t_L g205 ( .A(n_132), .B(n_137), .Y(n_205) );
AO21x2_ASAP7_75t_L g137 ( .A1(n_133), .A2(n_138), .B(n_155), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_133), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_133), .A2(n_197), .B(n_198), .Y(n_196) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_133), .A2(n_484), .B(n_488), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_133), .A2(n_527), .B(n_528), .Y(n_526) );
OA21x2_ASAP7_75t_L g627 ( .A1(n_133), .A2(n_484), .B(n_488), .Y(n_627) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_SL g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x4_ASAP7_75t_L g216 ( .A(n_135), .B(n_136), .Y(n_216) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_145), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g157 ( .A(n_142), .B(n_144), .Y(n_157) );
AND2x4_ASAP7_75t_L g175 ( .A(n_142), .B(n_152), .Y(n_175) );
HB1xp67_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x6_ASAP7_75t_L g156 ( .A(n_146), .B(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g162 ( .A(n_147), .Y(n_162) );
AND2x6_ASAP7_75t_L g173 ( .A(n_147), .B(n_150), .Y(n_173) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_154), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx5_ASAP7_75t_L g176 ( .A(n_154), .Y(n_176) );
AND2x4_ASAP7_75t_L g158 ( .A(n_157), .B(n_159), .Y(n_158) );
NOR2x1p5_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_164), .B(n_194), .Y(n_353) );
INVx1_ASAP7_75t_L g390 ( .A(n_164), .Y(n_390) );
AND2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_180), .Y(n_164) );
AND2x2_ASAP7_75t_L g204 ( .A(n_165), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g411 ( .A(n_165), .Y(n_411) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g254 ( .A(n_166), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_166), .B(n_180), .Y(n_255) );
AND2x2_ASAP7_75t_L g276 ( .A(n_166), .B(n_195), .Y(n_276) );
AND2x2_ASAP7_75t_L g358 ( .A(n_166), .B(n_181), .Y(n_358) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_169), .B(n_178), .Y(n_166) );
INVx4_ASAP7_75t_L g179 ( .A(n_167), .Y(n_179) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx4f_ASAP7_75t_L g190 ( .A(n_168), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_177), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_174), .B(n_176), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_173), .B(n_234), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_176), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_176), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_176), .A2(n_214), .B(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_176), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_176), .A2(n_232), .B(n_233), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_176), .A2(n_244), .B(n_245), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_176), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_176), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_176), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_176), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_176), .A2(n_530), .B(n_531), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_176), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_176), .A2(n_562), .B(n_563), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_176), .A2(n_578), .B(n_579), .Y(n_577) );
INVx3_ASAP7_75t_L g219 ( .A(n_179), .Y(n_219) );
AND2x4_ASAP7_75t_SL g251 ( .A(n_180), .B(n_195), .Y(n_251) );
INVx1_ASAP7_75t_L g282 ( .A(n_180), .Y(n_282) );
INVx2_ASAP7_75t_L g290 ( .A(n_180), .Y(n_290) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_180), .Y(n_314) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_181), .Y(n_203) );
AOI21x1_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_189), .Y(n_181) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_182), .A2(n_534), .B(n_540), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_188), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_190), .A2(n_229), .B(n_230), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_192), .B(n_204), .Y(n_191) );
AND2x2_ASAP7_75t_L g429 ( .A(n_192), .B(n_292), .Y(n_429) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_203), .Y(n_193) );
NAND2x1p5_ASAP7_75t_L g288 ( .A(n_194), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g340 ( .A(n_194), .B(n_255), .Y(n_340) );
AND2x2_ASAP7_75t_L g357 ( .A(n_194), .B(n_358), .Y(n_357) );
INVx4_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x4_ASAP7_75t_L g281 ( .A(n_195), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g297 ( .A(n_195), .Y(n_297) );
AND2x2_ASAP7_75t_L g341 ( .A(n_195), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g348 ( .A(n_195), .B(n_349), .Y(n_348) );
NOR2x1_ASAP7_75t_L g363 ( .A(n_195), .B(n_254), .Y(n_363) );
BUFx2_ASAP7_75t_L g373 ( .A(n_195), .Y(n_373) );
AND2x2_ASAP7_75t_L g398 ( .A(n_195), .B(n_358), .Y(n_398) );
AND2x2_ASAP7_75t_L g419 ( .A(n_195), .B(n_420), .Y(n_419) );
OR2x6_ASAP7_75t_L g195 ( .A(n_196), .B(n_202), .Y(n_195) );
INVx1_ASAP7_75t_L g350 ( .A(n_203), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_204), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g380 ( .A(n_204), .B(n_251), .Y(n_380) );
INVx3_ASAP7_75t_L g287 ( .A(n_205), .Y(n_287) );
AND2x2_ASAP7_75t_L g420 ( .A(n_205), .B(n_342), .Y(n_420) );
INVx1_ASAP7_75t_SL g206 ( .A(n_207), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_207), .A2(n_250), .B1(n_255), .B2(n_256), .Y(n_249) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_217), .Y(n_207) );
INVx4_ASAP7_75t_L g247 ( .A(n_208), .Y(n_247) );
INVx2_ASAP7_75t_L g284 ( .A(n_208), .Y(n_284) );
NAND2x1_ASAP7_75t_L g310 ( .A(n_208), .B(n_227), .Y(n_310) );
OR2x2_ASAP7_75t_L g325 ( .A(n_208), .B(n_260), .Y(n_325) );
OR2x2_ASAP7_75t_SL g352 ( .A(n_208), .B(n_324), .Y(n_352) );
AND2x2_ASAP7_75t_L g365 ( .A(n_208), .B(n_239), .Y(n_365) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_208), .Y(n_386) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_216), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_216), .A2(n_241), .B(n_242), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_216), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_SL g558 ( .A(n_216), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_216), .A2(n_575), .B(n_576), .Y(n_574) );
INVx2_ASAP7_75t_L g265 ( .A(n_217), .Y(n_265) );
AND2x2_ASAP7_75t_L g397 ( .A(n_217), .B(n_371), .Y(n_397) );
NOR2x1_ASAP7_75t_SL g217 ( .A(n_218), .B(n_227), .Y(n_217) );
AND2x2_ASAP7_75t_L g238 ( .A(n_218), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g414 ( .A(n_218), .B(n_337), .Y(n_414) );
AO21x1_ASAP7_75t_SL g218 ( .A1(n_219), .A2(n_220), .B(n_226), .Y(n_218) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_219), .A2(n_220), .B(n_226), .Y(n_261) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_219), .A2(n_493), .B(n_499), .Y(n_492) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_219), .A2(n_514), .B(n_520), .Y(n_513) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_219), .A2(n_514), .B(n_520), .Y(n_547) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_219), .A2(n_493), .B(n_499), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_225), .Y(n_220) );
OR2x2_ASAP7_75t_L g246 ( .A(n_227), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g257 ( .A(n_227), .B(n_247), .Y(n_257) );
AND2x2_ASAP7_75t_L g303 ( .A(n_227), .B(n_260), .Y(n_303) );
OR2x2_ASAP7_75t_L g324 ( .A(n_227), .B(n_239), .Y(n_324) );
INVx2_ASAP7_75t_SL g330 ( .A(n_227), .Y(n_330) );
AND2x2_ASAP7_75t_L g336 ( .A(n_227), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g346 ( .A(n_227), .B(n_329), .Y(n_346) );
BUFx2_ASAP7_75t_L g368 ( .A(n_227), .Y(n_368) );
OR2x6_ASAP7_75t_L g227 ( .A(n_228), .B(n_235), .Y(n_227) );
INVx2_ASAP7_75t_L g415 ( .A(n_236), .Y(n_415) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_246), .Y(n_236) );
OR2x2_ASAP7_75t_L g440 ( .A(n_237), .B(n_284), .Y(n_440) );
INVx2_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_238), .B(n_247), .Y(n_306) );
AND2x2_ASAP7_75t_L g377 ( .A(n_238), .B(n_257), .Y(n_377) );
INVx1_ASAP7_75t_L g259 ( .A(n_239), .Y(n_259) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_239), .Y(n_268) );
INVx1_ASAP7_75t_L g301 ( .A(n_239), .Y(n_301) );
INVx2_ASAP7_75t_L g337 ( .A(n_239), .Y(n_337) );
NOR2xp67_ASAP7_75t_L g267 ( .A(n_247), .B(n_268), .Y(n_267) );
BUFx2_ASAP7_75t_L g327 ( .A(n_247), .Y(n_327) );
INVx2_ASAP7_75t_SL g403 ( .A(n_248), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_250), .A2(n_305), .B1(n_307), .B2(n_311), .Y(n_304) );
AND2x2_ASAP7_75t_SL g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AND2x2_ASAP7_75t_L g431 ( .A(n_251), .B(n_287), .Y(n_431) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_253), .B(n_297), .Y(n_376) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g342 ( .A(n_254), .B(n_290), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_255), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g285 ( .A(n_256), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_256), .A2(n_400), .B1(n_404), .B2(n_406), .C(n_408), .Y(n_399) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
AND2x2_ASAP7_75t_L g269 ( .A(n_257), .B(n_270), .Y(n_269) );
INVxp67_ASAP7_75t_SL g293 ( .A(n_257), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_257), .B(n_300), .Y(n_355) );
INVx1_ASAP7_75t_SL g351 ( .A(n_258), .Y(n_351) );
AOI221xp5_ASAP7_75t_SL g379 ( .A1(n_258), .A2(n_269), .B1(n_380), .B2(n_381), .C(n_384), .Y(n_379) );
AOI322xp5_ASAP7_75t_L g412 ( .A1(n_258), .A2(n_330), .A3(n_357), .B1(n_413), .B2(n_415), .C1(n_416), .C2(n_419), .Y(n_412) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
BUFx2_ASAP7_75t_L g279 ( .A(n_259), .Y(n_279) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_260), .Y(n_271) );
INVx2_ASAP7_75t_L g329 ( .A(n_260), .Y(n_329) );
AND2x2_ASAP7_75t_L g370 ( .A(n_260), .B(n_371), .Y(n_370) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OA21x2_ASAP7_75t_SL g262 ( .A1(n_263), .A2(n_269), .B(n_272), .Y(n_262) );
AOI211xp5_ASAP7_75t_L g432 ( .A1(n_263), .A2(n_433), .B(n_434), .C(n_438), .Y(n_432) );
INVx1_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
OR2x2_ASAP7_75t_L g321 ( .A(n_265), .B(n_283), .Y(n_321) );
OR2x2_ASAP7_75t_L g405 ( .A(n_265), .B(n_300), .Y(n_405) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g345 ( .A(n_267), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g423 ( .A(n_270), .Y(n_423) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g309 ( .A(n_271), .Y(n_309) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
OR2x2_ASAP7_75t_L g278 ( .A(n_274), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g313 ( .A(n_276), .B(n_314), .Y(n_313) );
OAI322xp33_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_280), .A3(n_283), .B1(n_285), .B2(n_286), .C1(n_291), .C2(n_293), .Y(n_277) );
INVx1_ASAP7_75t_L g319 ( .A(n_278), .Y(n_319) );
OR2x2_ASAP7_75t_L g291 ( .A(n_280), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_280), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g302 ( .A(n_284), .B(n_303), .Y(n_302) );
OAI32xp33_ASAP7_75t_L g347 ( .A1(n_284), .A2(n_348), .A3(n_351), .B1(n_352), .B2(n_353), .Y(n_347) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx2_ASAP7_75t_L g292 ( .A(n_287), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_287), .B(n_350), .Y(n_349) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_287), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g413 ( .A(n_287), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g334 ( .A(n_288), .Y(n_334) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_292), .B(n_358), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_295), .B(n_315), .Y(n_294) );
OAI21xp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_298), .B(n_304), .Y(n_295) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x4_ASAP7_75t_SL g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g364 ( .A(n_303), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_306), .A2(n_326), .B1(n_428), .B2(n_430), .Y(n_427) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g354 ( .A1(n_308), .A2(n_355), .B(n_356), .C(n_359), .Y(n_354) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx3_ASAP7_75t_L g436 ( .A(n_310), .Y(n_436) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g317 ( .A(n_314), .Y(n_317) );
AO21x1_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_318), .B(n_322), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g382 ( .A(n_317), .Y(n_382) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_323), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g338 ( .A(n_325), .Y(n_338) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx1_ASAP7_75t_L g395 ( .A(n_328), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
NOR3xp33_ASAP7_75t_L g331 ( .A(n_332), .B(n_354), .C(n_366), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
OAI21xp5_ASAP7_75t_SL g396 ( .A1(n_335), .A2(n_397), .B(n_398), .Y(n_396) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx1_ASAP7_75t_L g371 ( .A(n_337), .Y(n_371) );
O2A1O1Ixp5_ASAP7_75t_SL g339 ( .A1(n_340), .A2(n_341), .B(n_343), .C(n_347), .Y(n_339) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_349), .Y(n_439) );
INVx2_ASAP7_75t_L g424 ( .A(n_352), .Y(n_424) );
AOI21xp33_ASAP7_75t_L g438 ( .A1(n_353), .A2(n_439), .B(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g418 ( .A(n_358), .Y(n_418) );
OAI31xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .A3(n_363), .B(n_364), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g437 ( .A(n_365), .Y(n_437) );
OAI21xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_372), .B(n_375), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
BUFx2_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g387 ( .A(n_370), .Y(n_387) );
AOI21xp33_ASAP7_75t_SL g434 ( .A1(n_372), .A2(n_435), .B(n_437), .Y(n_434) );
OR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx2_ASAP7_75t_L g402 ( .A(n_373), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_373), .B(n_393), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_373), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g383 ( .A(n_374), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
NAND5xp2_ASAP7_75t_L g378 ( .A(n_379), .B(n_399), .C(n_412), .D(n_421), .E(n_432), .Y(n_378) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_388), .B1(n_391), .B2(n_394), .C(n_396), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_425), .B(n_427), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g447 ( .A(n_441), .Y(n_447) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_L g459 ( .A(n_452), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_457), .B(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_757), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_468), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_463), .Y(n_462) );
CKINVDCx11_ASAP7_75t_R g469 ( .A(n_470), .Y(n_469) );
CKINVDCx6p67_ASAP7_75t_R g759 ( .A(n_470), .Y(n_759) );
INVx3_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_474), .Y(n_761) );
CKINVDCx11_ASAP7_75t_R g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND4xp75_ASAP7_75t_L g477 ( .A(n_478), .B(n_667), .C(n_707), .D(n_736), .Y(n_477) );
NOR2x1_ASAP7_75t_L g478 ( .A(n_479), .B(n_629), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_586), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_521), .B(n_541), .Y(n_480) );
AND2x2_ASAP7_75t_SL g481 ( .A(n_482), .B(n_489), .Y(n_481) );
AND2x4_ASAP7_75t_L g585 ( .A(n_482), .B(n_546), .Y(n_585) );
INVx1_ASAP7_75t_SL g638 ( .A(n_482), .Y(n_638) );
AOI21xp33_ASAP7_75t_L g673 ( .A1(n_482), .A2(n_674), .B(n_677), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_SL g677 ( .A1(n_482), .A2(n_678), .B(n_679), .C(n_680), .Y(n_677) );
NAND2x1_ASAP7_75t_L g718 ( .A(n_482), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_482), .B(n_679), .Y(n_740) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g544 ( .A(n_483), .Y(n_544) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_483), .Y(n_617) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_500), .Y(n_489) );
AND2x2_ASAP7_75t_L g609 ( .A(n_490), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g690 ( .A(n_490), .B(n_546), .Y(n_690) );
INVx1_ASAP7_75t_L g750 ( .A(n_490), .Y(n_750) );
BUFx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g594 ( .A(n_491), .B(n_512), .Y(n_594) );
AND2x2_ASAP7_75t_L g719 ( .A(n_491), .B(n_513), .Y(n_719) );
AND2x2_ASAP7_75t_L g724 ( .A(n_491), .B(n_684), .Y(n_724) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVxp67_ASAP7_75t_L g600 ( .A(n_492), .Y(n_600) );
BUFx3_ASAP7_75t_L g633 ( .A(n_492), .Y(n_633) );
AND2x2_ASAP7_75t_L g679 ( .A(n_492), .B(n_513), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_498), .Y(n_493) );
AND2x2_ASAP7_75t_L g664 ( .A(n_500), .B(n_543), .Y(n_664) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_512), .Y(n_500) );
AND2x4_ASAP7_75t_L g546 ( .A(n_501), .B(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g656 ( .A(n_501), .B(n_640), .Y(n_656) );
AND2x2_ASAP7_75t_SL g699 ( .A(n_501), .B(n_627), .Y(n_699) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx2_ASAP7_75t_L g635 ( .A(n_502), .Y(n_635) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g596 ( .A(n_503), .Y(n_596) );
OAI21x1_ASAP7_75t_SL g503 ( .A1(n_504), .A2(n_506), .B(n_510), .Y(n_503) );
INVx1_ASAP7_75t_L g511 ( .A(n_505), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_512), .B(n_596), .Y(n_599) );
AND2x2_ASAP7_75t_L g684 ( .A(n_512), .B(n_627), .Y(n_684) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g681 ( .A(n_513), .B(n_544), .Y(n_681) );
AND2x2_ASAP7_75t_L g701 ( .A(n_513), .B(n_627), .Y(n_701) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_515), .B(n_519), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_521), .B(n_590), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_521), .A2(n_713), .B1(n_714), .B2(n_715), .C(n_717), .Y(n_712) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OAI332xp33_ASAP7_75t_L g746 ( .A1(n_522), .A2(n_606), .A3(n_613), .B1(n_672), .B2(n_747), .B3(n_748), .C1(n_749), .C2(n_751), .Y(n_746) );
NAND2x1p5_ASAP7_75t_L g522 ( .A(n_523), .B(n_532), .Y(n_522) );
AND2x2_ASAP7_75t_L g552 ( .A(n_523), .B(n_533), .Y(n_552) );
AND2x2_ASAP7_75t_L g569 ( .A(n_523), .B(n_570), .Y(n_569) );
INVx4_ASAP7_75t_L g581 ( .A(n_523), .Y(n_581) );
AND2x2_ASAP7_75t_SL g641 ( .A(n_523), .B(n_582), .Y(n_641) );
INVx5_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NOR2x1_ASAP7_75t_SL g603 ( .A(n_524), .B(n_570), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_524), .B(n_532), .Y(n_607) );
AND2x2_ASAP7_75t_L g614 ( .A(n_524), .B(n_533), .Y(n_614) );
BUFx2_ASAP7_75t_L g649 ( .A(n_524), .Y(n_649) );
AND2x2_ASAP7_75t_L g704 ( .A(n_524), .B(n_573), .Y(n_704) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
OR2x2_ASAP7_75t_L g572 ( .A(n_532), .B(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g582 ( .A(n_532), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g622 ( .A(n_532), .Y(n_622) );
AND2x2_ASAP7_75t_L g692 ( .A(n_532), .B(n_591), .Y(n_692) );
AND2x2_ASAP7_75t_L g705 ( .A(n_532), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_532), .B(n_706), .Y(n_723) );
INVx4_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_533), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_539), .Y(n_534) );
OAI32xp33_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_548), .A3(n_553), .B1(n_567), .B2(n_584), .Y(n_541) );
INVx2_ASAP7_75t_L g650 ( .A(n_542), .Y(n_650) );
OR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
INVx1_ASAP7_75t_L g661 ( .A(n_543), .Y(n_661) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x4_ASAP7_75t_L g595 ( .A(n_544), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g728 ( .A(n_544), .B(n_633), .Y(n_728) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g640 ( .A(n_547), .Y(n_640) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
INVx2_ASAP7_75t_L g628 ( .A(n_550), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_550), .B(n_671), .Y(n_670) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x4_ASAP7_75t_SL g639 ( .A(n_551), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g716 ( .A(n_551), .Y(n_716) );
AND2x2_ASAP7_75t_L g734 ( .A(n_551), .B(n_596), .Y(n_734) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NOR2xp67_ASAP7_75t_SL g678 ( .A(n_554), .B(n_607), .Y(n_678) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_555), .B(n_589), .Y(n_676) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g752 ( .A(n_556), .B(n_622), .Y(n_752) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g583 ( .A(n_557), .Y(n_583) );
INVx2_ASAP7_75t_L g624 ( .A(n_557), .Y(n_624) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B(n_565), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_558), .B(n_566), .Y(n_565) );
AO21x2_ASAP7_75t_L g570 ( .A1(n_558), .A2(n_559), .B(n_565), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_564), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_580), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_568), .B(n_626), .Y(n_711) );
AND2x4_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
AND3x2_ASAP7_75t_L g666 ( .A(n_569), .B(n_613), .C(n_622), .Y(n_666) );
AND2x2_ASAP7_75t_L g590 ( .A(n_570), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_570), .B(n_573), .Y(n_647) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g601 ( .A(n_572), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g591 ( .A(n_573), .Y(n_591) );
INVx1_ASAP7_75t_L g606 ( .A(n_573), .Y(n_606) );
BUFx3_ASAP7_75t_L g613 ( .A(n_573), .Y(n_613) );
AND2x2_ASAP7_75t_L g623 ( .A(n_573), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AND2x4_ASAP7_75t_L g632 ( .A(n_581), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_581), .B(n_591), .Y(n_675) );
AND2x2_ASAP7_75t_L g631 ( .A(n_582), .B(n_606), .Y(n_631) );
INVx2_ASAP7_75t_L g658 ( .A(n_582), .Y(n_658) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
AOI211xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_592), .B(n_597), .C(n_618), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g738 ( .A1(n_587), .A2(n_714), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_590), .B(n_649), .Y(n_648) );
AOI211xp5_ASAP7_75t_SL g668 ( .A1(n_590), .A2(n_669), .B(n_673), .C(n_682), .Y(n_668) );
AND2x2_ASAP7_75t_L g654 ( .A(n_591), .B(n_614), .Y(n_654) );
OR2x2_ASAP7_75t_L g657 ( .A(n_591), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g744 ( .A(n_594), .B(n_699), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_595), .B(n_640), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_595), .A2(n_621), .B1(n_701), .B2(n_704), .C(n_710), .Y(n_709) );
AND2x4_ASAP7_75t_L g626 ( .A(n_596), .B(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g672 ( .A(n_596), .B(n_627), .Y(n_672) );
OAI221xp5_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_601), .B1(n_604), .B2(n_608), .C(n_611), .Y(n_597) );
AND2x2_ASAP7_75t_L g743 ( .A(n_598), .B(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g610 ( .A(n_599), .Y(n_610) );
INVx1_ASAP7_75t_L g696 ( .A(n_600), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_601), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g615 ( .A(n_603), .B(n_606), .Y(n_615) );
AND2x2_ASAP7_75t_L g691 ( .A(n_603), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g616 ( .A(n_610), .B(n_617), .Y(n_616) );
OAI21xp5_ASAP7_75t_SL g611 ( .A1(n_612), .A2(n_615), .B(n_616), .Y(n_611) );
INVx1_ASAP7_75t_L g735 ( .A(n_612), .Y(n_735) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g714 ( .A(n_613), .B(n_641), .Y(n_714) );
AND2x2_ASAP7_75t_SL g687 ( .A(n_614), .B(n_623), .Y(n_687) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B(n_625), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_619), .A2(n_653), .B1(n_656), .B2(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g725 ( .A(n_619), .Y(n_725) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g645 ( .A(n_622), .Y(n_645) );
INVx1_ASAP7_75t_L g706 ( .A(n_624), .Y(n_706) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_626), .B(n_628), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g747 ( .A(n_626), .B(n_696), .Y(n_747) );
AND2x2_ASAP7_75t_L g715 ( .A(n_627), .B(n_716), .Y(n_715) );
OAI211xp5_ASAP7_75t_L g708 ( .A1(n_628), .A2(n_709), .B(n_712), .C(n_720), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_651), .Y(n_629) );
AOI322xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .A3(n_634), .B1(n_636), .B2(n_641), .C1(n_642), .C2(n_650), .Y(n_630) );
CKINVDCx16_ASAP7_75t_R g748 ( .A(n_632), .Y(n_748) );
AND2x2_ASAP7_75t_L g698 ( .A(n_633), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g732 ( .A(n_633), .Y(n_732) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NOR2xp33_ASAP7_75t_SL g683 ( .A(n_635), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_SL g689 ( .A(n_635), .B(n_681), .Y(n_689) );
AND2x2_ASAP7_75t_L g713 ( .A(n_635), .B(n_679), .Y(n_713) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g685 ( .A(n_639), .Y(n_685) );
NAND2xp33_ASAP7_75t_SL g642 ( .A(n_643), .B(n_648), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI221xp5_ASAP7_75t_SL g688 ( .A1(n_644), .A2(n_689), .B1(n_690), .B2(n_691), .C(n_693), .Y(n_688) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVxp67_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g755 ( .A(n_647), .Y(n_755) );
AOI211xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B(n_655), .C(n_659), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g730 ( .A(n_654), .Y(n_730) );
INVx1_ASAP7_75t_L g662 ( .A(n_656), .Y(n_662) );
OR2x2_ASAP7_75t_L g749 ( .A(n_656), .B(n_750), .Y(n_749) );
INVx2_ASAP7_75t_SL g745 ( .A(n_657), .Y(n_745) );
AOI21xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B(n_665), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_661), .B(n_679), .Y(n_756) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_688), .Y(n_667) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_671), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
OR2x2_ASAP7_75t_L g722 ( .A(n_675), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI21xp33_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_685), .B(n_686), .Y(n_682) );
INVx2_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
AOI31xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_697), .A3(n_700), .B(n_702), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_699), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
AND2x4_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_724), .B1(n_725), .B2(n_726), .C(n_729), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B1(n_733), .B2(n_735), .Y(n_729) );
CKINVDCx16_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
NOR3xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_746), .C(n_753), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g737 ( .A(n_738), .B(n_741), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_745), .Y(n_741) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_756), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
BUFx4f_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
BUFx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_768), .Y(n_767) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_773), .Y(n_772) );
endmodule