module fake_jpeg_11763_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g49 ( 
.A(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_59),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_1),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_41),
.B1(n_48),
.B2(n_39),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_63),
.Y(n_65)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_54),
.B(n_43),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_63),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_74),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_40),
.B1(n_53),
.B2(n_38),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_48),
.B1(n_4),
.B2(n_5),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_77),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_82),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_38),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_83),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_3),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_85),
.Y(n_107)
);

NOR2x1_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_6),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_11),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_91),
.C(n_18),
.Y(n_101)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_12),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_66),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_97),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_84),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_101),
.Y(n_109)
);

AOI21x1_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_16),
.B(n_17),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_108),
.B(n_30),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_20),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_115),
.C(n_117),
.Y(n_120)
);

AOI22x1_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_21),
.B1(n_23),
.B2(n_26),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_104),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_116),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_28),
.C(n_29),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_112),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_113),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_123),
.Y(n_125)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_109),
.C(n_121),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_109),
.B(n_120),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_125),
.C(n_107),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_104),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_105),
.C(n_106),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_98),
.Y(n_130)
);


endmodule