module fake_jpeg_20296_n_286 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_286);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_286;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_48)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_22),
.B1(n_17),
.B2(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_18),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_23),
.B1(n_27),
.B2(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_34),
.A2(n_30),
.B1(n_17),
.B2(n_22),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_39),
.B1(n_37),
.B2(n_27),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_30),
.B1(n_17),
.B2(n_22),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_23),
.B1(n_29),
.B2(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_26),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_56),
.B(n_18),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_24),
.B1(n_16),
.B2(n_20),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_31),
.B1(n_1),
.B2(n_2),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_57),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_60),
.B(n_94),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_56),
.A2(n_26),
.B(n_25),
.C(n_29),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_61),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_44),
.B1(n_42),
.B2(n_41),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_62),
.A2(n_92),
.B1(n_101),
.B2(n_18),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_41),
.B1(n_36),
.B2(n_40),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_121)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_45),
.B1(n_35),
.B2(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx11_ASAP7_75t_SL g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_86),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_16),
.B1(n_20),
.B2(n_23),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_98),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_76),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_39),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_77),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_25),
.B1(n_35),
.B2(n_24),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_15),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_58),
.A2(n_31),
.B1(n_15),
.B2(n_24),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_81),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_15),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_31),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_88),
.Y(n_124)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_93),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_51),
.A2(n_24),
.B1(n_31),
.B2(n_18),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_31),
.Y(n_93)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_18),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_99),
.A2(n_100),
.B1(n_37),
.B2(n_39),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_54),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_48),
.A2(n_18),
.B1(n_32),
.B2(n_28),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_122),
.B1(n_101),
.B2(n_64),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_14),
.C(n_28),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_123),
.C(n_133),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_14),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_111),
.A2(n_88),
.B(n_73),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_81),
.A2(n_32),
.B1(n_28),
.B2(n_14),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_68),
.B(n_14),
.C(n_32),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_67),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_95),
.B1(n_71),
.B2(n_96),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_14),
.C(n_10),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_134),
.A2(n_159),
.B1(n_119),
.B2(n_115),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_104),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_139),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_128),
.B(n_60),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_136),
.B(n_154),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_98),
.B1(n_77),
.B2(n_62),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_137),
.A2(n_145),
.B1(n_148),
.B2(n_152),
.Y(n_186)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_104),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_77),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_141),
.A2(n_111),
.B(n_125),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_143),
.A2(n_106),
.B1(n_121),
.B2(n_127),
.Y(n_163)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_103),
.A2(n_79),
.B1(n_82),
.B2(n_72),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_70),
.B1(n_83),
.B2(n_97),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_61),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_145),
.Y(n_183)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_151),
.Y(n_165)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_120),
.A2(n_85),
.B1(n_89),
.B2(n_90),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_158),
.Y(n_167)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_156),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_131),
.A2(n_99),
.B1(n_91),
.B2(n_87),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_124),
.B(n_115),
.Y(n_182)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_173),
.B1(n_174),
.B2(n_122),
.Y(n_196)
);

AND2x6_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_131),
.Y(n_164)
);

XNOR2x1_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_133),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_170),
.B(n_172),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_120),
.C(n_123),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_148),
.C(n_159),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_142),
.B(n_125),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_152),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_126),
.B(n_116),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_121),
.B1(n_105),
.B2(n_110),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_137),
.A2(n_118),
.B1(n_129),
.B2(n_111),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_149),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_175),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_141),
.A2(n_153),
.B(n_139),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_176),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_138),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_185),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_183),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_155),
.A2(n_119),
.B1(n_118),
.B2(n_132),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_184),
.A2(n_151),
.B1(n_150),
.B2(n_129),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_144),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_186),
.A2(n_135),
.B1(n_154),
.B2(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_193),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_186),
.A2(n_173),
.B1(n_183),
.B2(n_163),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_205),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_158),
.C(n_156),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_201),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_199),
.B1(n_200),
.B2(n_209),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_172),
.B(n_182),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_157),
.B1(n_65),
.B2(n_132),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_147),
.B1(n_76),
.B2(n_140),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_147),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_0),
.C(n_1),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_203),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_0),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_0),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_207),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_0),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_178),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_185),
.B1(n_181),
.B2(n_170),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_221),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_214),
.B(n_1),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_167),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

NAND3xp33_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_180),
.C(n_179),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_217),
.B(n_2),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_191),
.A2(n_165),
.B(n_162),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_227),
.B(n_178),
.Y(n_243)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_180),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_191),
.A2(n_165),
.B(n_162),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_229),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_160),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_192),
.B1(n_196),
.B2(n_203),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_230),
.A2(n_238),
.B1(n_226),
.B2(n_222),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_194),
.C(n_193),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_234),
.C(n_236),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_221),
.B1(n_213),
.B2(n_216),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_237),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_200),
.B1(n_199),
.B2(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_190),
.C(n_201),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_205),
.C(n_179),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_160),
.C(n_202),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_171),
.B1(n_178),
.B2(n_204),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_171),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_239),
.B(n_3),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_215),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_225),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_3),
.B(n_4),
.Y(n_253)
);

NOR3xp33_ASAP7_75t_SL g254 ( 
.A(n_245),
.B(n_246),
.C(n_3),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_229),
.B1(n_224),
.B2(n_211),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_249),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_220),
.B1(n_222),
.B2(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

INVxp33_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_253),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_256),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_230),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_243),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_231),
.C(n_238),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_260),
.C(n_261),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_234),
.C(n_237),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_236),
.C(n_240),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_267),
.A2(n_253),
.B1(n_248),
.B2(n_257),
.Y(n_271)
);

OAI21xp33_ASAP7_75t_L g268 ( 
.A1(n_265),
.A2(n_251),
.B(n_244),
.Y(n_268)
);

AOI21x1_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_262),
.B(n_266),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_262),
.A2(n_249),
.B(n_247),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_271),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_274),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_250),
.C(n_245),
.Y(n_273)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_6),
.C(n_8),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_263),
.A2(n_254),
.B1(n_7),
.B2(n_8),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_272),
.Y(n_279)
);

OA21x2_ASAP7_75t_SL g281 ( 
.A1(n_278),
.A2(n_6),
.B(n_8),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_280),
.C(n_281),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_270),
.B1(n_268),
.B2(n_9),
.Y(n_280)
);

AOI21x1_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_275),
.B(n_9),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_283),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_9),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_9),
.Y(n_286)
);


endmodule