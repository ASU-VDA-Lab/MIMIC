module fake_aes_4193_n_32 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_32);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
OAI22xp5_ASAP7_75t_SL g12 ( .A1(n_2), .A2(n_3), .B1(n_4), .B2(n_0), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
XNOR2xp5_ASAP7_75t_L g16 ( .A(n_12), .B(n_1), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_14), .B(n_1), .Y(n_17) );
OR2x6_ASAP7_75t_L g18 ( .A(n_11), .B(n_2), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_17), .B(n_13), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_18), .B(n_11), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
NOR2xp33_ASAP7_75t_R g22 ( .A(n_19), .B(n_16), .Y(n_22) );
INVxp67_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
INVxp67_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
NAND2xp5_ASAP7_75t_SL g25 ( .A(n_23), .B(n_20), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_24), .B(n_22), .Y(n_26) );
AO22x2_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_15), .B1(n_13), .B2(n_18), .Y(n_27) );
OAI22xp5_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_3), .B1(n_5), .B2(n_6), .Y(n_28) );
CKINVDCx5p33_ASAP7_75t_R g29 ( .A(n_28), .Y(n_29) );
NAND2xp5_ASAP7_75t_L g30 ( .A(n_27), .B(n_6), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_30), .B(n_10), .Y(n_31) );
OAI22xp5_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_29), .B1(n_7), .B2(n_8), .Y(n_32) );
endmodule