module fake_jpeg_8222_n_335 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_37),
.B(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_20),
.B(n_7),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_6),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_24),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_17),
.Y(n_51)
);

HAxp5_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_78),
.CON(n_85),
.SN(n_85)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_54),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_56),
.B(n_63),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_26),
.B(n_33),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_57),
.A2(n_73),
.B(n_33),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_59),
.A2(n_67),
.B1(n_76),
.B2(n_33),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_68),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_71),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_26),
.B1(n_17),
.B2(n_24),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_34),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_44),
.B(n_17),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_77),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_24),
.B1(n_30),
.B2(n_35),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_27),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_29),
.B1(n_35),
.B2(n_34),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_83),
.A2(n_92),
.B1(n_94),
.B2(n_99),
.Y(n_126)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_86),
.B(n_98),
.Y(n_132)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_91),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_82),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_90),
.A2(n_100),
.B1(n_105),
.B2(n_106),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_52),
.A2(n_36),
.B1(n_21),
.B2(n_19),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_95),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_19),
.B1(n_21),
.B2(n_36),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_96),
.Y(n_150)
);

BUFx8_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_56),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_36),
.B1(n_21),
.B2(n_19),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_103),
.B(n_23),
.CI(n_31),
.CON(n_144),
.SN(n_144)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_58),
.A2(n_36),
.B1(n_21),
.B2(n_32),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_78),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_51),
.B(n_85),
.Y(n_127)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_32),
.B1(n_31),
.B2(n_23),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_75),
.B1(n_78),
.B2(n_70),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_71),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_61),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_122),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_123),
.B(n_139),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_87),
.B1(n_101),
.B2(n_89),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_73),
.C(n_51),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_146),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_135),
.A2(n_147),
.B1(n_148),
.B2(n_84),
.Y(n_156)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_50),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_48),
.Y(n_162)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_101),
.B(n_6),
.Y(n_174)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_85),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_50),
.B1(n_48),
.B2(n_81),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_50),
.B1(n_48),
.B2(n_81),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_112),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_115),
.Y(n_160)
);

AO22x1_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_144),
.B1(n_135),
.B2(n_148),
.Y(n_154)
);

AO22x1_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_171),
.B1(n_177),
.B2(n_168),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_136),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_155),
.B(n_158),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_171),
.B1(n_186),
.B2(n_121),
.Y(n_190)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_160),
.B(n_161),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_13),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_169),
.Y(n_189)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_177),
.C(n_32),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_125),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_124),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_180),
.Y(n_206)
);

OA22x2_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_144),
.B1(n_140),
.B2(n_110),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_87),
.B1(n_95),
.B2(n_96),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_173),
.A2(n_183),
.B1(n_138),
.B2(n_118),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_185),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_0),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_179),
.B(n_184),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_31),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_139),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_124),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_150),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_181),
.B(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_187),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_130),
.A2(n_122),
.B1(n_102),
.B2(n_100),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_145),
.A2(n_60),
.B1(n_98),
.B2(n_106),
.Y(n_184)
);

INVx13_ASAP7_75t_SL g185 ( 
.A(n_131),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_153),
.A2(n_88),
.B1(n_60),
.B2(n_90),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_131),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_153),
.B1(n_88),
.B2(n_134),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_188),
.A2(n_190),
.B1(n_194),
.B2(n_212),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_192),
.B(n_198),
.Y(n_225)
);

AND2x6_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_137),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_193),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_137),
.B1(n_134),
.B2(n_86),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_203),
.B1(n_214),
.B2(n_216),
.Y(n_221)
);

CKINVDCx12_ASAP7_75t_R g197 ( 
.A(n_179),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_183),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_205),
.Y(n_220)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_10),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_179),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_10),
.C(n_14),
.Y(n_240)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_167),
.B(n_28),
.Y(n_211)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_154),
.A2(n_138),
.B1(n_28),
.B2(n_23),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_165),
.A2(n_28),
.B1(n_39),
.B2(n_107),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_186),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_215),
.B(n_161),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_171),
.A2(n_28),
.B1(n_39),
.B2(n_97),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_171),
.A2(n_97),
.B1(n_1),
.B2(n_2),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_217),
.A2(n_178),
.B1(n_176),
.B2(n_158),
.Y(n_232)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_173),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_203),
.Y(n_230)
);

OAI21x1_ASAP7_75t_R g222 ( 
.A1(n_209),
.A2(n_166),
.B(n_182),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_222),
.A2(n_230),
.B(n_233),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_223),
.B(n_239),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_164),
.C(n_169),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_229),
.C(n_231),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_175),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_163),
.C(n_175),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_232),
.A2(n_15),
.B1(n_6),
.B2(n_4),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_204),
.A2(n_184),
.B(n_160),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_157),
.C(n_1),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_242),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_216),
.B(n_210),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_238),
.B(n_191),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_157),
.Y(n_237)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_0),
.B(n_2),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_191),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_210),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_241),
.B(n_244),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_201),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_246),
.Y(n_250)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_196),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_247),
.B(n_260),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_226),
.A2(n_219),
.B1(n_190),
.B2(n_195),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_251),
.A2(n_255),
.B1(n_263),
.B2(n_236),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_236),
.A2(n_213),
.B1(n_217),
.B2(n_195),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_235),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_212),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_221),
.C(n_234),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_224),
.A2(n_194),
.B1(n_213),
.B2(n_188),
.Y(n_255)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_192),
.Y(n_257)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_257),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_245),
.B(n_205),
.Y(n_260)
);

NOR3xp33_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_211),
.C(n_202),
.Y(n_262)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_226),
.A2(n_202),
.B1(n_214),
.B2(n_218),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_220),
.B(n_11),
.Y(n_264)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_237),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_268),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_266),
.Y(n_270)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_225),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_229),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_273),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_233),
.B(n_227),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_276),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_275),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_221),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_249),
.A2(n_227),
.B(n_230),
.Y(n_276)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_242),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_256),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_222),
.B1(n_243),
.B2(n_232),
.Y(n_280)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_222),
.C(n_243),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_253),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_264),
.Y(n_289)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_258),
.Y(n_290)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_296),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_259),
.Y(n_294)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_250),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_295),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_250),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_298),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_251),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_273),
.C(n_279),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_270),
.A2(n_265),
.B1(n_261),
.B2(n_267),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_300),
.B(n_261),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_307),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g305 ( 
.A(n_299),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_307),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_SL g306 ( 
.A1(n_296),
.A2(n_278),
.A3(n_271),
.B1(n_252),
.B2(n_274),
.C1(n_275),
.C2(n_280),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_306),
.B(n_291),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_281),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_287),
.A2(n_284),
.B(n_276),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_311),
.A2(n_297),
.B(n_277),
.Y(n_313)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_312),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_313),
.A2(n_314),
.B(n_320),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_301),
.Y(n_322)
);

NOR2x1_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_293),
.Y(n_318)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_318),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_302),
.B(n_263),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_319),
.Y(n_323)
);

OAI321xp33_ASAP7_75t_L g320 ( 
.A1(n_311),
.A2(n_238),
.A3(n_288),
.B1(n_4),
.B2(n_5),
.C(n_12),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_325),
.C(n_288),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_304),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_318),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_309),
.B(n_303),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_327),
.A2(n_329),
.B(n_325),
.C(n_323),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_321),
.A2(n_317),
.B(n_316),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_328),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_330),
.A2(n_324),
.B(n_310),
.Y(n_332)
);

AOI322xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_331),
.A3(n_310),
.B1(n_5),
.B2(n_13),
.C1(n_14),
.C2(n_3),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_13),
.B(n_2),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_3),
.Y(n_335)
);


endmodule