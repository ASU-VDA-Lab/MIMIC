module fake_jpeg_18194_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_10),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_38),
.Y(n_56)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_32),
.B1(n_33),
.B2(n_24),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_46),
.A2(n_60),
.B1(n_61),
.B2(n_65),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_47),
.B(n_58),
.Y(n_102)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_50),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_30),
.Y(n_81)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_23),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_32),
.B1(n_33),
.B2(n_24),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_32),
.B1(n_33),
.B2(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_67),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_33),
.B1(n_32),
.B2(n_24),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_68),
.B1(n_20),
.B2(n_18),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_32),
.B1(n_19),
.B2(n_27),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_29),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_29),
.C(n_17),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_35),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_23),
.B1(n_17),
.B2(n_31),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_16),
.B(n_34),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_48),
.C(n_69),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_73),
.Y(n_111)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_35),
.B(n_34),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_31),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_99),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_22),
.B1(n_30),
.B2(n_19),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_76),
.A2(n_79),
.B1(n_90),
.B2(n_100),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_80),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_81),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_21),
.B1(n_30),
.B2(n_19),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_31),
.B1(n_18),
.B2(n_20),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_27),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_83),
.Y(n_130)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_85),
.Y(n_120)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_20),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_28),
.Y(n_125)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_88),
.A2(n_103),
.B1(n_108),
.B2(n_51),
.Y(n_131)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_94),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_66),
.Y(n_94)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_97),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_11),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

CKINVDCx12_ASAP7_75t_R g118 ( 
.A(n_98),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_66),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_27),
.B1(n_22),
.B2(n_21),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_48),
.A2(n_22),
.B1(n_21),
.B2(n_17),
.Y(n_103)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_18),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_110),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_63),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_1),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_125),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_71),
.A2(n_50),
.B1(n_55),
.B2(n_52),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_124),
.B1(n_127),
.B2(n_135),
.Y(n_143)
);

AOI22x1_ASAP7_75t_SL g117 ( 
.A1(n_86),
.A2(n_55),
.B1(n_59),
.B2(n_57),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_98),
.B1(n_107),
.B2(n_94),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_78),
.A2(n_55),
.B1(n_57),
.B2(n_59),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_74),
.A2(n_28),
.B1(n_51),
.B2(n_3),
.Y(n_127)
);

NAND2xp33_ASAP7_75t_SL g129 ( 
.A(n_80),
.B(n_28),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_72),
.B(n_99),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_131),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_89),
.A2(n_51),
.B1(n_14),
.B2(n_13),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_93),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_106),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_14),
.C(n_13),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_140),
.C(n_70),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_13),
.C(n_12),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_141),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_142),
.A2(n_156),
.B1(n_165),
.B2(n_129),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_75),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_134),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_147),
.B(n_164),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_119),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_151),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_SL g202 ( 
.A(n_150),
.B(n_167),
.C(n_101),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_153),
.A2(n_158),
.B(n_95),
.Y(n_196)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_104),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_155),
.B(n_171),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_117),
.A2(n_80),
.B1(n_104),
.B2(n_90),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_159),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_87),
.B(n_83),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_110),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_168),
.Y(n_181)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_77),
.C(n_87),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_114),
.C(n_125),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_109),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_117),
.A2(n_80),
.B1(n_83),
.B2(n_96),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_132),
.A2(n_88),
.B1(n_82),
.B2(n_109),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_166),
.A2(n_95),
.B1(n_82),
.B2(n_91),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_122),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_85),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_136),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_130),
.B(n_111),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_111),
.B(n_12),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_172),
.B(n_137),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_195),
.C(n_150),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_143),
.A2(n_128),
.B1(n_116),
.B2(n_121),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_178),
.A2(n_192),
.B1(n_144),
.B2(n_152),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_132),
.B(n_118),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_140),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_180),
.B(n_196),
.Y(n_215)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_187),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_185),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_121),
.Y(n_185)
);

AND2x6_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_118),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_188),
.A2(n_189),
.B1(n_203),
.B2(n_145),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_124),
.B1(n_112),
.B2(n_127),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_153),
.A2(n_112),
.B1(n_123),
.B2(n_133),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_84),
.Y(n_194)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_194),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_123),
.C(n_105),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_108),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_201),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_151),
.B(n_101),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_157),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_212),
.B1(n_214),
.B2(n_225),
.Y(n_232)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_219),
.C(n_220),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_184),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_210),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_143),
.B1(n_155),
.B2(n_172),
.Y(n_212)
);

XNOR2x2_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_158),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_213),
.B(n_11),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_176),
.A2(n_170),
.B1(n_169),
.B2(n_154),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_189),
.B1(n_188),
.B2(n_193),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_217),
.A2(n_229),
.B1(n_197),
.B2(n_190),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_148),
.C(n_146),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_162),
.C(n_159),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_221),
.A2(n_149),
.B1(n_2),
.B2(n_3),
.Y(n_249)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_224),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_181),
.A2(n_147),
.B1(n_141),
.B2(n_95),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_186),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_193),
.A2(n_181),
.B1(n_177),
.B2(n_201),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_149),
.C(n_12),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_180),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_218),
.Y(n_255)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_196),
.B(n_179),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_235),
.A2(n_223),
.B(n_2),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_177),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_242),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_175),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_243),
.Y(n_256)
);

OAI22x1_ASAP7_75t_SL g239 ( 
.A1(n_217),
.A2(n_173),
.B1(n_182),
.B2(n_202),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_239),
.A2(n_207),
.B1(n_228),
.B2(n_211),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_175),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_205),
.B(n_11),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_250),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_248),
.A2(n_213),
.B1(n_230),
.B2(n_221),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_249),
.Y(n_254)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_220),
.C(n_209),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_260),
.C(n_263),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_261),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_232),
.B1(n_233),
.B2(n_239),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_268),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_219),
.C(n_221),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_218),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_204),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_262),
.B(n_266),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_229),
.C(n_223),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_264),
.A2(n_234),
.B(n_251),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_226),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_267),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_240),
.B(n_1),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_2),
.C(n_4),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_241),
.C(n_244),
.Y(n_283)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_235),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_282),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_245),
.B(n_248),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_275),
.A2(n_250),
.B(n_244),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_238),
.Y(n_276)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_278),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_256),
.A2(n_233),
.B1(n_254),
.B2(n_247),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_283),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_241),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_252),
.C(n_263),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_293),
.C(n_271),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_283),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_294),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_269),
.Y(n_288)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_274),
.A2(n_273),
.B(n_277),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_289),
.A2(n_295),
.B1(n_4),
.B2(n_6),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_257),
.C(n_259),
.Y(n_293)
);

OAI31xp33_ASAP7_75t_L g295 ( 
.A1(n_270),
.A2(n_257),
.A3(n_5),
.B(n_6),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_290),
.A2(n_281),
.B1(n_272),
.B2(n_282),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_299),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_297),
.B(n_298),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_291),
.B(n_271),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_4),
.C(n_5),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_295),
.A3(n_302),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_7),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_6),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_303),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_300),
.A2(n_287),
.B(n_289),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_305),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_299),
.A2(n_293),
.B1(n_292),
.B2(n_286),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_308),
.B(n_309),
.C(n_297),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_311),
.B(n_307),
.Y(n_313)
);

NAND4xp25_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_301),
.C(n_296),
.D(n_292),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_313),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_6),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_314),
.A3(n_310),
.B1(n_9),
.B2(n_10),
.C1(n_8),
.C2(n_7),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_8),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_10),
.Y(n_318)
);


endmodule