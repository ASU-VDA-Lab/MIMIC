module fake_jpeg_12967_n_441 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_441);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_441;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_48),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_7),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_49),
.B(n_54),
.Y(n_103)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_26),
.B(n_7),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_26),
.B(n_7),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_57),
.B(n_58),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_59),
.B(n_63),
.Y(n_132)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_23),
.B(n_7),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_66),
.B(n_69),
.Y(n_137)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_22),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_67),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

INVx2_ASAP7_75t_R g77 ( 
.A(n_17),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_77),
.B(n_88),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_19),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_80),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_79),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_6),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx6_ASAP7_75t_SL g85 ( 
.A(n_21),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_91),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_23),
.B(n_6),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_87),
.B(n_14),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_19),
.A2(n_6),
.B1(n_2),
.B2(n_3),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_90),
.A2(n_27),
.B1(n_30),
.B2(n_34),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_19),
.B(n_8),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_8),
.Y(n_112)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_95),
.B(n_122),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_47),
.A2(n_42),
.B1(n_46),
.B2(n_16),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_97),
.A2(n_37),
.B1(n_76),
.B2(n_65),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_31),
.B1(n_39),
.B2(n_42),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_98),
.A2(n_70),
.B1(n_64),
.B2(n_82),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_92),
.A2(n_42),
.B1(n_39),
.B2(n_40),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_99),
.A2(n_72),
.B1(n_86),
.B2(n_84),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_40),
.B1(n_38),
.B2(n_34),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_104),
.A2(n_139),
.B1(n_35),
.B2(n_16),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_77),
.B(n_21),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_105),
.B(n_21),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_123),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_50),
.B(n_38),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_51),
.A2(n_39),
.B1(n_17),
.B2(n_46),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_48),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_131),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_60),
.B(n_27),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_61),
.B(n_30),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_142),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_67),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_8),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_73),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_148),
.B(n_154),
.Y(n_209)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_132),
.B(n_83),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_150),
.B(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_153),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_32),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_157),
.Y(n_193)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_156),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_118),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_158),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_159),
.A2(n_169),
.B1(n_175),
.B2(n_183),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_118),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_171),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_113),
.B(n_55),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_163),
.A2(n_189),
.B1(n_127),
.B2(n_140),
.Y(n_222)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_165),
.A2(n_172),
.B1(n_180),
.B2(n_115),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_167),
.Y(n_192)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_105),
.B(n_75),
.C(n_74),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_179),
.C(n_138),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_L g169 ( 
.A1(n_97),
.A2(n_93),
.B1(n_89),
.B2(n_94),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_105),
.B(n_46),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_170),
.B(n_181),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_129),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_70),
.B1(n_35),
.B2(n_16),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_176),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_139),
.A2(n_68),
.B1(n_81),
.B2(n_79),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_184),
.Y(n_213)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_71),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_117),
.A2(n_35),
.B1(n_37),
.B2(n_52),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_134),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_103),
.A2(n_37),
.B(n_0),
.C(n_3),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_182),
.A2(n_2),
.B(n_4),
.C(n_5),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_96),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_0),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_185),
.B(n_186),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_116),
.B(n_2),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_123),
.A2(n_98),
.B1(n_143),
.B2(n_120),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_187),
.A2(n_115),
.B1(n_107),
.B2(n_127),
.Y(n_191)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_143),
.A2(n_53),
.B1(n_88),
.B2(n_56),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_191),
.A2(n_215),
.B1(n_181),
.B2(n_162),
.Y(n_227)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_163),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_SL g232 ( 
.A1(n_195),
.A2(n_200),
.B(n_223),
.C(n_225),
.Y(n_232)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_148),
.B(n_136),
.CI(n_135),
.CON(n_199),
.SN(n_199)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_199),
.B(n_221),
.Y(n_253)
);

AO22x1_ASAP7_75t_L g200 ( 
.A1(n_154),
.A2(n_100),
.B1(n_130),
.B2(n_107),
.Y(n_200)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_201),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_161),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_152),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

XNOR2x1_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_166),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_175),
.A2(n_147),
.B1(n_119),
.B2(n_101),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_182),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_152),
.B(n_130),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_220),
.B(n_186),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g221 ( 
.A(n_168),
.B(n_136),
.CI(n_100),
.CON(n_221),
.SN(n_221)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_222),
.A2(n_179),
.B1(n_159),
.B2(n_190),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_166),
.A2(n_91),
.B(n_147),
.C(n_101),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_157),
.A2(n_140),
.B1(n_114),
.B2(n_109),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_183),
.B(n_179),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_160),
.A2(n_114),
.B1(n_109),
.B2(n_102),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_226),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_227),
.A2(n_234),
.B1(n_252),
.B2(n_223),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_229),
.B(n_240),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_206),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_247),
.Y(n_259)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_211),
.A2(n_150),
.B1(n_161),
.B2(n_151),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_235),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_236),
.A2(n_239),
.B1(n_241),
.B2(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_246),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_222),
.B1(n_201),
.B2(n_211),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_171),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_209),
.A2(n_166),
.B1(n_151),
.B2(n_170),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_242),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_249),
.C(n_212),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_201),
.A2(n_167),
.B1(n_164),
.B2(n_153),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_245),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_185),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_193),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_194),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_251),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_202),
.B(n_179),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_250),
.B(n_254),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_194),
.B(n_182),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_215),
.A2(n_173),
.B1(n_177),
.B2(n_102),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_173),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_277),
.C(n_281),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_253),
.A2(n_233),
.B(n_238),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_260),
.A2(n_200),
.B(n_232),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_261),
.B(n_266),
.Y(n_295)
);

HAxp5_ASAP7_75t_SL g264 ( 
.A(n_247),
.B(n_221),
.CON(n_264),
.SN(n_264)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_267),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_213),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_240),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_221),
.B1(n_199),
.B2(n_192),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_269),
.A2(n_283),
.B1(n_253),
.B2(n_245),
.Y(n_292)
);

AOI22x1_ASAP7_75t_L g271 ( 
.A1(n_227),
.A2(n_199),
.B1(n_195),
.B2(n_191),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_271),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_244),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_236),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_202),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_246),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_239),
.A2(n_224),
.B1(n_195),
.B2(n_192),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_276),
.A2(n_226),
.B1(n_242),
.B2(n_232),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_192),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_241),
.B(n_217),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_251),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_210),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_231),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_252),
.A2(n_195),
.B1(n_200),
.B2(n_210),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_259),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_290),
.Y(n_311)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_256),
.Y(n_287)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_287),
.Y(n_337)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_256),
.Y(n_288)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_291),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_292),
.A2(n_308),
.B1(n_285),
.B2(n_279),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_258),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_229),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_294),
.B(n_296),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_237),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_298),
.A2(n_300),
.B1(n_310),
.B2(n_283),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_276),
.A2(n_255),
.B1(n_232),
.B2(n_235),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_274),
.B(n_254),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_302),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_250),
.Y(n_302)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_303),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_305),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_259),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_184),
.C(n_232),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_277),
.C(n_281),
.Y(n_312)
);

A2O1A1O1Ixp25_ASAP7_75t_L g307 ( 
.A1(n_262),
.A2(n_232),
.B(n_228),
.C(n_216),
.D(n_219),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_309),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_261),
.A2(n_255),
.B1(n_228),
.B2(n_196),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g309 ( 
.A1(n_263),
.A2(n_265),
.A3(n_274),
.B1(n_262),
.B2(n_260),
.C1(n_269),
.C2(n_258),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_265),
.A2(n_196),
.B1(n_218),
.B2(n_216),
.Y(n_310)
);

MAJx2_ASAP7_75t_L g354 ( 
.A(n_312),
.B(n_309),
.C(n_291),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_277),
.C(n_278),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_316),
.C(n_324),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_315),
.A2(n_327),
.B1(n_303),
.B2(n_310),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_278),
.C(n_263),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_317),
.B(n_271),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_275),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_322),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_295),
.Y(n_320)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_320),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_280),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_295),
.Y(n_323)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_323),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_280),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_285),
.A2(n_279),
.B1(n_272),
.B2(n_271),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_272),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_334),
.C(n_319),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_329),
.A2(n_308),
.B1(n_305),
.B2(n_307),
.Y(n_342)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_286),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_297),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_299),
.B(n_266),
.Y(n_334)
);

OAI22x1_ASAP7_75t_L g335 ( 
.A1(n_298),
.A2(n_271),
.B1(n_273),
.B2(n_282),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_335),
.Y(n_356)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_299),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_338),
.B(n_343),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_284),
.Y(n_340)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_340),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_341),
.A2(n_335),
.B1(n_327),
.B2(n_315),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_342),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_324),
.B(n_290),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_345),
.B(n_318),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_326),
.A2(n_307),
.B1(n_296),
.B2(n_302),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_348),
.A2(n_357),
.B1(n_346),
.B2(n_347),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_301),
.C(n_304),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_350),
.B(n_322),
.C(n_317),
.Y(n_366)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_328),
.Y(n_351)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_351),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_352),
.Y(n_370)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_311),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_358),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_354),
.B(n_359),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_313),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_331),
.A2(n_288),
.B1(n_287),
.B2(n_196),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_333),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_332),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_321),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_360),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_350),
.A2(n_330),
.B(n_312),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_361),
.B(n_366),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_373),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_339),
.B(n_337),
.C(n_325),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_371),
.B(n_374),
.C(n_378),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_338),
.C(n_344),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_375),
.B(n_178),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_357),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_376),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_343),
.B(n_203),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_377),
.B(n_345),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_219),
.C(n_198),
.Y(n_378)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_379),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_380),
.B(n_386),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_363),
.B(n_348),
.Y(n_382)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_382),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_354),
.C(n_355),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_388),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_377),
.B(n_342),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_367),
.A2(n_356),
.B1(n_349),
.B2(n_218),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_387),
.A2(n_383),
.B1(n_367),
.B2(n_391),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_365),
.B(n_356),
.C(n_198),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_364),
.Y(n_389)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_389),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_368),
.A2(n_155),
.B(n_188),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_391),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_370),
.B(n_218),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_375),
.Y(n_409)
);

INVx11_ASAP7_75t_L g395 ( 
.A(n_371),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_395),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_393),
.B(n_378),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_394),
.C(n_203),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_362),
.Y(n_400)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_400),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_381),
.B(n_365),
.C(n_366),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_401),
.A2(n_403),
.B(n_407),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_SL g419 ( 
.A(n_402),
.B(n_409),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_373),
.C(n_372),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_392),
.B(n_369),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_404),
.B(n_382),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_395),
.B(n_384),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_408),
.B(n_388),
.C(n_386),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_412),
.B(n_415),
.Y(n_422)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_413),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_401),
.A2(n_387),
.B(n_390),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_414),
.A2(n_417),
.B(n_420),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_396),
.B(n_380),
.C(n_393),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_418),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_403),
.A2(n_197),
.B(n_158),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_176),
.C(n_174),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_405),
.B(n_398),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_410),
.A2(n_406),
.B(n_397),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_423),
.A2(n_419),
.B(n_5),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_412),
.Y(n_424)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_424),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_396),
.C(n_409),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_425),
.B(n_4),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_415),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_427),
.A2(n_9),
.B1(n_11),
.B2(n_14),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_428),
.A2(n_419),
.B1(n_156),
.B2(n_9),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_429),
.B(n_9),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_430),
.A2(n_431),
.B(n_432),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_433),
.A2(n_422),
.B(n_421),
.Y(n_434)
);

OAI21x1_ASAP7_75t_SL g437 ( 
.A1(n_434),
.A2(n_436),
.B(n_424),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_437),
.B(n_438),
.C(n_11),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_435),
.A2(n_426),
.B(n_11),
.Y(n_438)
);

AO21x2_ASAP7_75t_L g440 ( 
.A1(n_439),
.A2(n_11),
.B(n_15),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_440),
.A2(n_15),
.B(n_182),
.Y(n_441)
);


endmodule