module fake_aes_7559_n_1068 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1068);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1068;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_968;
wire n_1042;
wire n_1060;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1011;
wire n_1025;
wire n_880;
wire n_630;
wire n_511;
wire n_1002;
wire n_467;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1063;
wire n_767;
wire n_828;
wire n_1014;
wire n_293;
wire n_506;
wire n_533;
wire n_490;
wire n_393;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_875;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_716;
wire n_653;
wire n_899;
wire n_806;
wire n_881;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_721;
wire n_438;
wire n_656;
wire n_640;
wire n_908;
wire n_955;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_912;
wire n_620;
wire n_841;
wire n_947;
wire n_924;
wire n_1043;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_992;
INVx1_ASAP7_75t_L g278 ( .A(n_110), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_69), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_102), .Y(n_280) );
CKINVDCx16_ASAP7_75t_R g281 ( .A(n_21), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_62), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_234), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_70), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_206), .Y(n_285) );
CKINVDCx16_ASAP7_75t_R g286 ( .A(n_14), .Y(n_286) );
INVxp67_ASAP7_75t_L g287 ( .A(n_237), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_72), .Y(n_288) );
INVxp67_ASAP7_75t_SL g289 ( .A(n_225), .Y(n_289) );
BUFx10_ASAP7_75t_L g290 ( .A(n_245), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_177), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_114), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_164), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_129), .B(n_8), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_131), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_266), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_73), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_276), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_128), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_238), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_263), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_187), .Y(n_302) );
CKINVDCx16_ASAP7_75t_R g303 ( .A(n_16), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_40), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_2), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_145), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_47), .Y(n_307) );
BUFx3_ASAP7_75t_L g308 ( .A(n_106), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_82), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_149), .Y(n_310) );
BUFx10_ASAP7_75t_L g311 ( .A(n_84), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_173), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_116), .B(n_33), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_25), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_182), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_242), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_105), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_27), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_44), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_134), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_179), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_162), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_271), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_256), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_217), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_58), .Y(n_326) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_133), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_197), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_201), .Y(n_329) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_188), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_207), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_75), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_49), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_153), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_147), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_180), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_121), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_198), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_252), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_208), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_250), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_146), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_118), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_5), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_235), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_178), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_261), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_89), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_190), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_8), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_60), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_37), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_144), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_189), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_66), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_199), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_113), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_186), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_73), .Y(n_359) );
CKINVDCx20_ASAP7_75t_R g360 ( .A(n_171), .Y(n_360) );
CKINVDCx14_ASAP7_75t_R g361 ( .A(n_130), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_45), .B(n_36), .Y(n_362) );
NOR2xp67_ASAP7_75t_L g363 ( .A(n_9), .B(n_230), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_170), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_247), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_120), .Y(n_366) );
BUFx3_ASAP7_75t_L g367 ( .A(n_59), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_6), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_165), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_226), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_90), .Y(n_371) );
INVxp33_ASAP7_75t_L g372 ( .A(n_243), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_72), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_185), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_202), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_233), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_181), .Y(n_377) );
INVx1_ASAP7_75t_SL g378 ( .A(n_107), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_126), .Y(n_379) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_232), .Y(n_380) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_91), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_135), .B(n_141), .Y(n_382) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_174), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_191), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_172), .B(n_137), .Y(n_385) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_169), .Y(n_386) );
CKINVDCx14_ASAP7_75t_R g387 ( .A(n_50), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_55), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_151), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g390 ( .A(n_93), .Y(n_390) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_251), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_117), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_209), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_267), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_262), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_167), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_88), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_223), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_86), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_38), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_213), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_102), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_132), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_54), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_11), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_29), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_290), .Y(n_407) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_349), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_312), .Y(n_409) );
OAI22xp5_ASAP7_75t_SL g410 ( .A1(n_318), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_312), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_322), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_282), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_387), .A2(n_286), .B1(n_303), .B2(n_281), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_322), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_372), .B(n_0), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_282), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_291), .B(n_3), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_387), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_368), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_288), .Y(n_421) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_349), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_284), .B(n_4), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_284), .B(n_7), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_324), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_304), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_326), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_324), .Y(n_428) );
AOI22x1_ASAP7_75t_SL g429 ( .A1(n_344), .A2(n_11), .B1(n_9), .B2(n_10), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_354), .Y(n_430) );
BUFx8_ASAP7_75t_L g431 ( .A(n_323), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_326), .Y(n_432) );
AND2x6_ASAP7_75t_L g433 ( .A(n_301), .B(n_115), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_354), .Y(n_434) );
INVx3_ASAP7_75t_L g435 ( .A(n_290), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_370), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_333), .Y(n_437) );
NOR2x1_ASAP7_75t_L g438 ( .A(n_308), .B(n_314), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_308), .B(n_12), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_321), .B(n_13), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_408), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_426), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_409), .Y(n_443) );
OR2x6_ASAP7_75t_L g444 ( .A(n_410), .B(n_358), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_407), .B(n_372), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_409), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_416), .A2(n_360), .B1(n_379), .B2(n_327), .Y(n_447) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_423), .B(n_285), .C(n_283), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_407), .B(n_287), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_411), .Y(n_450) );
BUFx4f_ASAP7_75t_L g451 ( .A(n_433), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_407), .B(n_361), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_435), .B(n_369), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_408), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_423), .A2(n_279), .B1(n_280), .B2(n_278), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_408), .Y(n_456) );
BUFx3_ASAP7_75t_L g457 ( .A(n_433), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_435), .B(n_370), .Y(n_458) );
BUFx8_ASAP7_75t_SL g459 ( .A(n_419), .Y(n_459) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_422), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_412), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_412), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_435), .B(n_361), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_415), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_422), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_415), .Y(n_466) );
INVx3_ASAP7_75t_L g467 ( .A(n_423), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_423), .A2(n_297), .B1(n_305), .B2(n_292), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_425), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_420), .B(n_424), .Y(n_470) );
INVx4_ASAP7_75t_L g471 ( .A(n_433), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_424), .A2(n_309), .B1(n_317), .B2(n_307), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_438), .B(n_425), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_431), .B(n_306), .Y(n_474) );
BUFx2_ASAP7_75t_L g475 ( .A(n_424), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_428), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_442), .B(n_414), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_443), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_445), .B(n_440), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_449), .B(n_418), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_453), .B(n_439), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_470), .B(n_413), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_452), .B(n_438), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_446), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_452), .B(n_401), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_442), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_463), .B(n_403), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_451), .A2(n_430), .B(n_428), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_450), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_463), .B(n_433), .Y(n_490) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_457), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g492 ( .A(n_474), .B(n_319), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_470), .B(n_433), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_470), .B(n_433), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_455), .A2(n_472), .B1(n_468), .B2(n_475), .Y(n_495) );
NOR2xp33_ASAP7_75t_SL g496 ( .A(n_471), .B(n_327), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_458), .B(n_433), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g498 ( .A(n_455), .B(n_399), .C(n_352), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_447), .B(n_352), .Y(n_499) );
INVx5_ASAP7_75t_L g500 ( .A(n_467), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_467), .B(n_437), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_467), .B(n_437), .Y(n_502) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_467), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_451), .B(n_293), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_448), .B(n_417), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_451), .B(n_299), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_448), .B(n_417), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_461), .B(n_421), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_462), .A2(n_434), .B1(n_430), .B2(n_436), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_464), .B(n_432), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_473), .B(n_427), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_473), .B(n_432), .Y(n_512) );
NAND2xp33_ASAP7_75t_L g513 ( .A(n_451), .B(n_382), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_447), .B(n_311), .Y(n_514) );
INVx2_ASAP7_75t_SL g515 ( .A(n_464), .Y(n_515) );
INVx8_ASAP7_75t_L g516 ( .A(n_459), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_457), .B(n_466), .Y(n_517) );
AND2x6_ASAP7_75t_L g518 ( .A(n_469), .B(n_301), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_476), .B(n_300), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_476), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_441), .A2(n_296), .B(n_295), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_444), .B(n_298), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_444), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_444), .B(n_316), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_441), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_441), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_444), .B(n_302), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_454), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_465), .B(n_311), .Y(n_529) );
INVx4_ASAP7_75t_L g530 ( .A(n_460), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_460), .B(n_328), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_465), .Y(n_532) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_460), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_486), .B(n_477), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_490), .A2(n_330), .B(n_289), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_479), .B(n_399), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_482), .B(n_400), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_482), .B(n_404), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_497), .A2(n_380), .B(n_310), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_524), .B(n_429), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_480), .B(n_406), .Y(n_541) );
INVx4_ASAP7_75t_L g542 ( .A(n_500), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_515), .A2(n_388), .B1(n_390), .B2(n_348), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_500), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_496), .B(n_331), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_501), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g547 ( .A1(n_481), .A2(n_362), .B(n_367), .C(n_314), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_491), .B(n_339), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_493), .A2(n_320), .B(n_315), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_502), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_485), .B(n_341), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_494), .A2(n_329), .B(n_325), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_SL g553 ( .A1(n_480), .A2(n_294), .B(n_313), .C(n_385), .Y(n_553) );
AO32x1_ASAP7_75t_L g554 ( .A1(n_530), .A2(n_334), .A3(n_337), .B1(n_336), .B2(n_335), .Y(n_554) );
BUFx3_ASAP7_75t_L g555 ( .A(n_516), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_503), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_513), .A2(n_340), .B(n_338), .Y(n_557) );
NOR2xp33_ASAP7_75t_SL g558 ( .A(n_523), .B(n_311), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_522), .A2(n_402), .B1(n_367), .B2(n_332), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_487), .B(n_342), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_503), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_516), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_499), .B(n_378), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_514), .B(n_381), .Y(n_564) );
NOR2xp67_ASAP7_75t_SL g565 ( .A(n_498), .B(n_500), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_512), .B(n_397), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_488), .A2(n_345), .B(n_343), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_511), .B(n_350), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_522), .B(n_351), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_527), .A2(n_402), .B1(n_355), .B2(n_359), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_517), .A2(n_347), .B(n_346), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_483), .A2(n_356), .B(n_353), .Y(n_572) );
BUFx3_ASAP7_75t_L g573 ( .A(n_516), .Y(n_573) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_478), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_492), .B(n_371), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_529), .B(n_373), .Y(n_576) );
OR2x6_ASAP7_75t_L g577 ( .A(n_505), .B(n_507), .Y(n_577) );
INVx3_ASAP7_75t_L g578 ( .A(n_484), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_519), .A2(n_365), .B(n_364), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_504), .A2(n_374), .B(n_366), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_506), .A2(n_376), .B(n_375), .Y(n_581) );
A2O1A1Ixp33_ASAP7_75t_L g582 ( .A1(n_489), .A2(n_405), .B(n_313), .C(n_294), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_520), .B(n_357), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_509), .A2(n_384), .B1(n_389), .B2(n_377), .Y(n_584) );
A2O1A1Ixp33_ASAP7_75t_L g585 ( .A1(n_521), .A2(n_363), .B(n_394), .C(n_392), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_508), .B(n_15), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_510), .Y(n_587) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_518), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_509), .A2(n_396), .B1(n_398), .B2(n_395), .Y(n_589) );
AO21x1_ASAP7_75t_L g590 ( .A1(n_530), .A2(n_385), .B(n_456), .Y(n_590) );
BUFx4f_ASAP7_75t_L g591 ( .A(n_533), .Y(n_591) );
O2A1O1Ixp33_ASAP7_75t_L g592 ( .A1(n_531), .A2(n_18), .B(n_16), .C(n_17), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_L g593 ( .A1(n_532), .A2(n_383), .B(n_386), .C(n_349), .Y(n_593) );
A2O1A1Ixp33_ASAP7_75t_L g594 ( .A1(n_525), .A2(n_528), .B(n_526), .C(n_383), .Y(n_594) );
A2O1A1Ixp33_ASAP7_75t_L g595 ( .A1(n_533), .A2(n_383), .B(n_386), .C(n_349), .Y(n_595) );
CKINVDCx16_ASAP7_75t_R g596 ( .A(n_533), .Y(n_596) );
AOI22x1_ASAP7_75t_L g597 ( .A1(n_488), .A2(n_422), .B1(n_386), .B2(n_391), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_501), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_500), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_501), .Y(n_600) );
O2A1O1Ixp33_ASAP7_75t_L g601 ( .A1(n_495), .A2(n_21), .B(n_19), .C(n_20), .Y(n_601) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_486), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_495), .A2(n_393), .B1(n_391), .B2(n_422), .Y(n_603) );
NAND3xp33_ASAP7_75t_L g604 ( .A(n_481), .B(n_393), .C(n_391), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_486), .A2(n_22), .B1(n_19), .B2(n_20), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_479), .B(n_22), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_495), .A2(n_26), .B1(n_23), .B2(n_24), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_479), .B(n_24), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_501), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_495), .A2(n_29), .B1(n_26), .B2(n_28), .Y(n_610) );
OAI21xp5_ASAP7_75t_L g611 ( .A1(n_493), .A2(n_122), .B(n_119), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_490), .A2(n_124), .B(n_123), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_495), .A2(n_32), .B1(n_30), .B2(n_31), .Y(n_613) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_491), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_486), .B(n_34), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_501), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g617 ( .A1(n_495), .A2(n_36), .B(n_34), .C(n_35), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_522), .A2(n_40), .B1(n_37), .B2(n_39), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_486), .B(n_39), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_501), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_501), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_486), .B(n_41), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_602), .Y(n_623) );
OAI21xp5_ASAP7_75t_L g624 ( .A1(n_549), .A2(n_127), .B(n_125), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_587), .Y(n_625) );
AO31x2_ASAP7_75t_L g626 ( .A1(n_590), .A2(n_43), .A3(n_41), .B(n_42), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_578), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_534), .B(n_43), .Y(n_628) );
AO31x2_ASAP7_75t_L g629 ( .A1(n_603), .A2(n_46), .A3(n_44), .B(n_45), .Y(n_629) );
INVx4_ASAP7_75t_L g630 ( .A(n_596), .Y(n_630) );
AO31x2_ASAP7_75t_L g631 ( .A1(n_547), .A2(n_48), .A3(n_46), .B(n_47), .Y(n_631) );
INVx3_ASAP7_75t_L g632 ( .A(n_542), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_L g633 ( .A1(n_601), .A2(n_53), .B(n_51), .C(n_52), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_556), .Y(n_634) );
AO31x2_ASAP7_75t_L g635 ( .A1(n_585), .A2(n_59), .A3(n_56), .B(n_57), .Y(n_635) );
BUFx2_ASAP7_75t_L g636 ( .A(n_543), .Y(n_636) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_553), .A2(n_63), .B(n_57), .C(n_61), .Y(n_637) );
OAI21xp5_ASAP7_75t_L g638 ( .A1(n_552), .A2(n_138), .B(n_136), .Y(n_638) );
A2O1A1Ixp33_ASAP7_75t_L g639 ( .A1(n_617), .A2(n_64), .B(n_65), .C(n_66), .Y(n_639) );
AO31x2_ASAP7_75t_L g640 ( .A1(n_594), .A2(n_67), .A3(n_68), .B(n_69), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_539), .A2(n_140), .B(n_139), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_558), .B(n_67), .C(n_70), .Y(n_642) );
INVx5_ASAP7_75t_L g643 ( .A(n_588), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_606), .A2(n_143), .B(n_142), .Y(n_644) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_591), .Y(n_645) );
INVx3_ASAP7_75t_L g646 ( .A(n_542), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_608), .A2(n_150), .B(n_148), .Y(n_647) );
A2O1A1Ixp33_ASAP7_75t_L g648 ( .A1(n_557), .A2(n_71), .B(n_74), .C(n_75), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_546), .A2(n_76), .B1(n_77), .B2(n_78), .Y(n_649) );
AO31x2_ASAP7_75t_L g650 ( .A1(n_582), .A2(n_76), .A3(n_77), .B(n_79), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_536), .B(n_80), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_561), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_564), .B(n_81), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_586), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_535), .A2(n_154), .B(n_152), .Y(n_655) );
NAND3xp33_ASAP7_75t_L g656 ( .A(n_558), .B(n_82), .C(n_83), .Y(n_656) );
OAI21x1_ASAP7_75t_L g657 ( .A1(n_597), .A2(n_156), .B(n_155), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_562), .Y(n_658) );
BUFx12f_ASAP7_75t_L g659 ( .A(n_555), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_550), .A2(n_83), .B1(n_85), .B2(n_86), .Y(n_660) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_567), .A2(n_158), .B(n_157), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_598), .B(n_85), .Y(n_662) );
OAI21x1_ASAP7_75t_L g663 ( .A1(n_612), .A2(n_160), .B(n_159), .Y(n_663) );
AO21x1_ASAP7_75t_L g664 ( .A1(n_607), .A2(n_163), .B(n_161), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_600), .A2(n_168), .B(n_166), .Y(n_665) );
CKINVDCx6p67_ASAP7_75t_R g666 ( .A(n_573), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_579), .A2(n_87), .B(n_88), .C(n_89), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_609), .B(n_87), .Y(n_668) );
AO21x1_ASAP7_75t_L g669 ( .A1(n_619), .A2(n_176), .B(n_175), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_540), .A2(n_91), .B1(n_92), .B2(n_93), .Y(n_670) );
AO21x1_ASAP7_75t_L g671 ( .A1(n_592), .A2(n_184), .B(n_183), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_583), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_574), .Y(n_673) );
OR2x2_ASAP7_75t_L g674 ( .A(n_563), .B(n_94), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_616), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_620), .B(n_95), .Y(n_676) );
OAI21x1_ASAP7_75t_L g677 ( .A1(n_604), .A2(n_224), .B(n_275), .Y(n_677) );
INVx3_ASAP7_75t_L g678 ( .A(n_591), .Y(n_678) );
OAI21xp5_ASAP7_75t_L g679 ( .A1(n_621), .A2(n_222), .B(n_274), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g680 ( .A1(n_571), .A2(n_221), .B(n_273), .Y(n_680) );
AO31x2_ASAP7_75t_L g681 ( .A1(n_593), .A2(n_95), .A3(n_96), .B(n_97), .Y(n_681) );
AO31x2_ASAP7_75t_L g682 ( .A1(n_595), .A2(n_98), .A3(n_99), .B(n_100), .Y(n_682) );
OAI21x1_ASAP7_75t_L g683 ( .A1(n_580), .A2(n_228), .B(n_272), .Y(n_683) );
OAI21x1_ASAP7_75t_L g684 ( .A1(n_581), .A2(n_227), .B(n_270), .Y(n_684) );
AO31x2_ASAP7_75t_L g685 ( .A1(n_584), .A2(n_101), .A3(n_103), .B(n_104), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_577), .A2(n_220), .B(n_269), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_569), .A2(n_103), .B1(n_104), .B2(n_105), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_577), .A2(n_231), .B(n_268), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_577), .A2(n_229), .B(n_265), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_541), .B(n_106), .Y(n_690) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_614), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_622), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_537), .B(n_108), .Y(n_693) );
AO32x2_ASAP7_75t_L g694 ( .A1(n_589), .A2(n_109), .A3(n_110), .B1(n_111), .B2(n_112), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_551), .A2(n_236), .B(n_264), .Y(n_695) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_574), .Y(n_696) );
O2A1O1Ixp33_ASAP7_75t_SL g697 ( .A1(n_545), .A2(n_219), .B(n_260), .C(n_259), .Y(n_697) );
AOI21xp33_ASAP7_75t_L g698 ( .A1(n_538), .A2(n_109), .B(n_111), .Y(n_698) );
OAI21xp5_ASAP7_75t_L g699 ( .A1(n_572), .A2(n_192), .B(n_193), .Y(n_699) );
OA21x2_ASAP7_75t_L g700 ( .A1(n_568), .A2(n_575), .B(n_618), .Y(n_700) );
OAI22x1_ASAP7_75t_L g701 ( .A1(n_605), .A2(n_194), .B1(n_195), .B2(n_196), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_560), .A2(n_200), .B(n_203), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g703 ( .A1(n_566), .A2(n_204), .B(n_205), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_576), .A2(n_210), .B(n_211), .Y(n_704) );
AO21x1_ASAP7_75t_L g705 ( .A1(n_615), .A2(n_212), .B(n_214), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_570), .B(n_215), .Y(n_706) );
OR2x6_ASAP7_75t_L g707 ( .A(n_544), .B(n_216), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_559), .B(n_218), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_599), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_565), .Y(n_710) );
A2O1A1Ixp33_ASAP7_75t_L g711 ( .A1(n_548), .A2(n_239), .B(n_240), .C(n_241), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_554), .Y(n_712) );
OAI21xp5_ASAP7_75t_L g713 ( .A1(n_549), .A2(n_244), .B(n_246), .Y(n_713) );
INVx3_ASAP7_75t_L g714 ( .A(n_596), .Y(n_714) );
OAI21xp5_ASAP7_75t_L g715 ( .A1(n_549), .A2(n_248), .B(n_249), .Y(n_715) );
INVx2_ASAP7_75t_SL g716 ( .A(n_602), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_602), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_601), .A2(n_253), .B(n_254), .C(n_255), .Y(n_718) );
O2A1O1Ixp33_ASAP7_75t_L g719 ( .A1(n_553), .A2(n_257), .B(n_258), .C(n_277), .Y(n_719) );
AOI221x1_ASAP7_75t_L g720 ( .A1(n_603), .A2(n_607), .B1(n_613), .B2(n_610), .C(n_604), .Y(n_720) );
INVx1_ASAP7_75t_SL g721 ( .A(n_602), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_602), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_578), .Y(n_723) );
AO21x1_ASAP7_75t_L g724 ( .A1(n_611), .A2(n_603), .B(n_601), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_625), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_636), .B(n_721), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_675), .Y(n_727) );
OR2x6_ASAP7_75t_L g728 ( .A(n_707), .B(n_630), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_675), .Y(n_729) );
AO31x2_ASAP7_75t_L g730 ( .A1(n_712), .A2(n_724), .A3(n_671), .B(n_705), .Y(n_730) );
INVx3_ASAP7_75t_L g731 ( .A(n_645), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_717), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_634), .Y(n_733) );
AO31x2_ASAP7_75t_L g734 ( .A1(n_664), .A2(n_720), .A3(n_718), .B(n_669), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_722), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_652), .Y(n_736) );
OR2x2_ASAP7_75t_L g737 ( .A(n_623), .B(n_716), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_672), .B(n_654), .Y(n_738) );
OR2x2_ASAP7_75t_L g739 ( .A(n_674), .B(n_714), .Y(n_739) );
OAI21xp5_ASAP7_75t_L g740 ( .A1(n_662), .A2(n_676), .B(n_668), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g741 ( .A1(n_633), .A2(n_639), .B(n_693), .Y(n_741) );
INVx3_ASAP7_75t_L g742 ( .A(n_645), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_653), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_649), .Y(n_744) );
OAI21x1_ASAP7_75t_SL g745 ( .A1(n_680), .A2(n_699), .B(n_661), .Y(n_745) );
INVx3_ASAP7_75t_L g746 ( .A(n_645), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_709), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_700), .B(n_628), .Y(n_748) );
OA21x2_ASAP7_75t_L g749 ( .A1(n_657), .A2(n_677), .B(n_715), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_660), .Y(n_750) );
OA21x2_ASAP7_75t_L g751 ( .A1(n_624), .A2(n_638), .B(n_713), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_700), .B(n_690), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_709), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_650), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_685), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_626), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_692), .B(n_651), .Y(n_757) );
OR2x6_ASAP7_75t_L g758 ( .A(n_707), .B(n_678), .Y(n_758) );
AO31x2_ASAP7_75t_L g759 ( .A1(n_701), .A2(n_710), .A3(n_648), .B(n_688), .Y(n_759) );
AO31x2_ASAP7_75t_L g760 ( .A1(n_686), .A2(n_689), .A3(n_667), .B(n_647), .Y(n_760) );
A2O1A1Ixp33_ASAP7_75t_L g761 ( .A1(n_698), .A2(n_706), .B(n_642), .C(n_656), .Y(n_761) );
OA21x2_ASAP7_75t_L g762 ( .A1(n_663), .A2(n_683), .B(n_684), .Y(n_762) );
BUFx8_ASAP7_75t_L g763 ( .A(n_694), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_627), .B(n_723), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_685), .Y(n_765) );
NAND2x1p5_ASAP7_75t_L g766 ( .A(n_678), .B(n_643), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_708), .B(n_632), .Y(n_767) );
BUFx2_ASAP7_75t_L g768 ( .A(n_666), .Y(n_768) );
AO21x2_ASAP7_75t_L g769 ( .A1(n_644), .A2(n_704), .B(n_665), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_687), .Y(n_770) );
A2O1A1Ixp33_ASAP7_75t_L g771 ( .A1(n_670), .A2(n_655), .B(n_641), .C(n_695), .Y(n_771) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_646), .Y(n_772) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_696), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_631), .B(n_635), .Y(n_774) );
BUFx3_ASAP7_75t_L g775 ( .A(n_691), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_694), .Y(n_776) );
AO21x2_ASAP7_75t_L g777 ( .A1(n_711), .A2(n_697), .B(n_702), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_694), .B(n_635), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_631), .Y(n_779) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_673), .Y(n_780) );
BUFx2_ASAP7_75t_L g781 ( .A(n_629), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_640), .B(n_629), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_681), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_682), .Y(n_784) );
BUFx8_ASAP7_75t_L g785 ( .A(n_659), .Y(n_785) );
OR2x2_ASAP7_75t_L g786 ( .A(n_721), .B(n_486), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_675), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_675), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_675), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_625), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_625), .B(n_675), .Y(n_791) );
BUFx2_ASAP7_75t_L g792 ( .A(n_630), .Y(n_792) );
AO31x2_ASAP7_75t_L g793 ( .A1(n_712), .A2(n_590), .A3(n_724), .B(n_671), .Y(n_793) );
OAI21x1_ASAP7_75t_SL g794 ( .A1(n_679), .A2(n_664), .B(n_703), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_625), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_625), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_658), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_625), .Y(n_798) );
BUFx12f_ASAP7_75t_L g799 ( .A(n_659), .Y(n_799) );
AO31x2_ASAP7_75t_L g800 ( .A1(n_712), .A2(n_590), .A3(n_724), .B(n_671), .Y(n_800) );
INVx4_ASAP7_75t_SL g801 ( .A(n_659), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_625), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_625), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_625), .B(n_675), .Y(n_804) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_721), .Y(n_805) );
OR2x6_ASAP7_75t_L g806 ( .A(n_707), .B(n_516), .Y(n_806) );
NAND3xp33_ASAP7_75t_L g807 ( .A(n_637), .B(n_719), .C(n_720), .Y(n_807) );
INVx2_ASAP7_75t_L g808 ( .A(n_675), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_791), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_727), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_729), .Y(n_811) );
BUFx6f_ASAP7_75t_L g812 ( .A(n_775), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_787), .Y(n_813) );
INVx3_ASAP7_75t_L g814 ( .A(n_758), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_732), .Y(n_815) );
INVx5_ASAP7_75t_L g816 ( .A(n_728), .Y(n_816) );
AND2x2_ASAP7_75t_L g817 ( .A(n_747), .B(n_788), .Y(n_817) );
OR2x2_ASAP7_75t_L g818 ( .A(n_804), .B(n_786), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_789), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_808), .Y(n_820) );
OR2x2_ASAP7_75t_L g821 ( .A(n_748), .B(n_753), .Y(n_821) );
BUFx2_ASAP7_75t_L g822 ( .A(n_728), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_725), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_735), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_790), .B(n_795), .Y(n_825) );
HB1xp67_ASAP7_75t_SL g826 ( .A(n_785), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_796), .B(n_798), .Y(n_827) );
AO21x2_ASAP7_75t_L g828 ( .A1(n_782), .A2(n_745), .B(n_794), .Y(n_828) );
AND2x2_ASAP7_75t_L g829 ( .A(n_802), .B(n_803), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_738), .B(n_726), .Y(n_830) );
INVx3_ASAP7_75t_L g831 ( .A(n_766), .Y(n_831) );
AND2x2_ASAP7_75t_L g832 ( .A(n_733), .B(n_736), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_755), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_765), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_784), .Y(n_835) );
AO21x2_ASAP7_75t_L g836 ( .A1(n_752), .A2(n_807), .B(n_754), .Y(n_836) );
AND2x2_ASAP7_75t_L g837 ( .A(n_778), .B(n_743), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_737), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_739), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_805), .Y(n_840) );
BUFx2_ASAP7_75t_L g841 ( .A(n_763), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_779), .Y(n_842) );
AND2x2_ASAP7_75t_L g843 ( .A(n_770), .B(n_744), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_776), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_750), .B(n_741), .Y(n_845) );
AND2x2_ASAP7_75t_L g846 ( .A(n_741), .B(n_781), .Y(n_846) );
AND2x2_ASAP7_75t_L g847 ( .A(n_756), .B(n_772), .Y(n_847) );
INVx1_ASAP7_75t_SL g848 ( .A(n_797), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_757), .B(n_774), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_757), .B(n_764), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_764), .B(n_740), .Y(n_851) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_792), .Y(n_852) );
AND2x2_ASAP7_75t_L g853 ( .A(n_740), .B(n_783), .Y(n_853) );
BUFx3_ASAP7_75t_L g854 ( .A(n_768), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_773), .B(n_780), .Y(n_855) );
INVx2_ASAP7_75t_L g856 ( .A(n_793), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_800), .Y(n_857) );
BUFx2_ASAP7_75t_L g858 ( .A(n_806), .Y(n_858) );
NAND2x1p5_ASAP7_75t_L g859 ( .A(n_731), .B(n_746), .Y(n_859) );
OAI21xp5_ASAP7_75t_L g860 ( .A1(n_761), .A2(n_771), .B(n_767), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_759), .B(n_746), .Y(n_861) );
INVx2_ASAP7_75t_L g862 ( .A(n_762), .Y(n_862) );
OR2x6_ASAP7_75t_L g863 ( .A(n_742), .B(n_751), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_742), .B(n_759), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_730), .B(n_734), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_730), .Y(n_866) );
INVx3_ASAP7_75t_L g867 ( .A(n_760), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_730), .B(n_734), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_850), .B(n_801), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_837), .B(n_734), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_837), .B(n_760), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_850), .B(n_760), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_845), .B(n_749), .Y(n_873) );
AND2x4_ASAP7_75t_L g874 ( .A(n_861), .B(n_769), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_845), .B(n_777), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_849), .B(n_777), .Y(n_876) );
AND2x2_ASAP7_75t_L g877 ( .A(n_849), .B(n_799), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_815), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_824), .Y(n_879) );
BUFx2_ASAP7_75t_L g880 ( .A(n_852), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_818), .B(n_830), .Y(n_881) );
AND2x4_ASAP7_75t_L g882 ( .A(n_861), .B(n_841), .Y(n_882) );
INVx5_ASAP7_75t_L g883 ( .A(n_816), .Y(n_883) );
AND2x4_ASAP7_75t_L g884 ( .A(n_841), .B(n_853), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_846), .B(n_843), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_825), .B(n_827), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_829), .B(n_851), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_829), .B(n_839), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_851), .B(n_823), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_821), .B(n_810), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_838), .B(n_832), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_810), .B(n_811), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_811), .B(n_813), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_817), .Y(n_894) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_855), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_817), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_813), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_819), .B(n_820), .Y(n_898) );
AND2x4_ASAP7_75t_L g899 ( .A(n_833), .B(n_834), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_844), .B(n_833), .Y(n_900) );
BUFx3_ASAP7_75t_L g901 ( .A(n_854), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_840), .Y(n_902) );
AND2x4_ASAP7_75t_L g903 ( .A(n_834), .B(n_835), .Y(n_903) );
AND2x4_ASAP7_75t_L g904 ( .A(n_835), .B(n_842), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_844), .B(n_809), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_847), .B(n_842), .Y(n_906) );
BUFx3_ASAP7_75t_L g907 ( .A(n_831), .Y(n_907) );
INVx2_ASAP7_75t_L g908 ( .A(n_862), .Y(n_908) );
AND2x2_ASAP7_75t_SL g909 ( .A(n_822), .B(n_858), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_847), .B(n_865), .Y(n_910) );
AND2x4_ASAP7_75t_L g911 ( .A(n_816), .B(n_863), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_865), .B(n_868), .Y(n_912) );
AND2x4_ASAP7_75t_L g913 ( .A(n_863), .B(n_814), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_908), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_900), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_912), .B(n_868), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_912), .B(n_828), .Y(n_917) );
INVx5_ASAP7_75t_L g918 ( .A(n_883), .Y(n_918) );
INVxp67_ASAP7_75t_SL g919 ( .A(n_880), .Y(n_919) );
HB1xp67_ASAP7_75t_L g920 ( .A(n_895), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_900), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_885), .B(n_828), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_885), .B(n_828), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_899), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_910), .B(n_857), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_899), .Y(n_926) );
NOR2xp33_ASAP7_75t_L g927 ( .A(n_869), .B(n_848), .Y(n_927) );
AND2x4_ASAP7_75t_L g928 ( .A(n_874), .B(n_863), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_871), .B(n_887), .Y(n_929) );
INVx4_ASAP7_75t_L g930 ( .A(n_883), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_903), .Y(n_931) );
NAND2xp5_ASAP7_75t_SL g932 ( .A(n_883), .B(n_812), .Y(n_932) );
AND2x2_ASAP7_75t_L g933 ( .A(n_871), .B(n_866), .Y(n_933) );
OR2x2_ASAP7_75t_L g934 ( .A(n_872), .B(n_864), .Y(n_934) );
INVx1_ASAP7_75t_SL g935 ( .A(n_901), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_906), .B(n_836), .Y(n_936) );
HB1xp67_ASAP7_75t_L g937 ( .A(n_901), .Y(n_937) );
OR2x2_ASAP7_75t_L g938 ( .A(n_886), .B(n_836), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_904), .Y(n_939) );
HB1xp67_ASAP7_75t_L g940 ( .A(n_892), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_870), .B(n_876), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_905), .Y(n_942) );
HB1xp67_ASAP7_75t_L g943 ( .A(n_892), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_905), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_870), .B(n_867), .Y(n_945) );
HB1xp67_ASAP7_75t_L g946 ( .A(n_893), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_876), .B(n_867), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_897), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_893), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_889), .B(n_856), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_898), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_898), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_929), .B(n_875), .Y(n_953) );
HB1xp67_ASAP7_75t_L g954 ( .A(n_920), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_948), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_948), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_929), .B(n_873), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_941), .B(n_873), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_949), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_942), .B(n_944), .Y(n_960) );
INVx3_ASAP7_75t_L g961 ( .A(n_930), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_949), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_941), .B(n_874), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_951), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_951), .Y(n_965) );
AND2x4_ASAP7_75t_SL g966 ( .A(n_930), .B(n_911), .Y(n_966) );
AND2x2_ASAP7_75t_L g967 ( .A(n_917), .B(n_874), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_942), .B(n_902), .Y(n_968) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_937), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_952), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_952), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_944), .B(n_894), .Y(n_972) );
INVx4_ASAP7_75t_L g973 ( .A(n_918), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_915), .Y(n_974) );
HB1xp67_ASAP7_75t_L g975 ( .A(n_935), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_915), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_921), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_921), .B(n_896), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_917), .B(n_882), .Y(n_979) );
OR2x2_ASAP7_75t_L g980 ( .A(n_940), .B(n_884), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_916), .B(n_913), .Y(n_981) );
INVx2_ASAP7_75t_L g982 ( .A(n_914), .Y(n_982) );
INVx3_ASAP7_75t_L g983 ( .A(n_930), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_922), .B(n_913), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_922), .B(n_913), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_923), .B(n_890), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_950), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_943), .B(n_878), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_936), .Y(n_989) );
AOI21xp5_ASAP7_75t_L g990 ( .A1(n_932), .A2(n_860), .B(n_909), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_923), .B(n_890), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_946), .B(n_879), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_953), .B(n_925), .Y(n_993) );
HB1xp67_ASAP7_75t_L g994 ( .A(n_969), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_960), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_957), .B(n_945), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_955), .Y(n_997) );
HB1xp67_ASAP7_75t_L g998 ( .A(n_954), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_953), .B(n_925), .Y(n_999) );
AOI22x1_ASAP7_75t_L g1000 ( .A1(n_973), .A2(n_919), .B1(n_826), .B2(n_877), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_956), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_986), .B(n_933), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_974), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_974), .Y(n_1004) );
OR2x2_ASAP7_75t_L g1005 ( .A(n_989), .B(n_934), .Y(n_1005) );
HB1xp67_ASAP7_75t_L g1006 ( .A(n_975), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_986), .B(n_933), .Y(n_1007) );
INVx2_ASAP7_75t_L g1008 ( .A(n_982), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_957), .B(n_945), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_956), .Y(n_1010) );
INVxp67_ASAP7_75t_SL g1011 ( .A(n_961), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_958), .B(n_947), .Y(n_1012) );
HB1xp67_ASAP7_75t_L g1013 ( .A(n_980), .Y(n_1013) );
INVx2_ASAP7_75t_L g1014 ( .A(n_982), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_976), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_958), .B(n_947), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_977), .Y(n_1017) );
INVxp67_ASAP7_75t_L g1018 ( .A(n_988), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_959), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1005), .Y(n_1020) );
OAI21xp5_ASAP7_75t_L g1021 ( .A1(n_1000), .A2(n_990), .B(n_973), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_995), .B(n_989), .Y(n_1022) );
OAI221xp5_ASAP7_75t_L g1023 ( .A1(n_1018), .A2(n_992), .B1(n_968), .B2(n_927), .C(n_983), .Y(n_1023) );
INVxp67_ASAP7_75t_L g1024 ( .A(n_998), .Y(n_1024) );
AND2x4_ASAP7_75t_L g1025 ( .A(n_1011), .B(n_966), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_994), .B(n_959), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_1012), .B(n_963), .Y(n_1027) );
INVxp67_ASAP7_75t_L g1028 ( .A(n_1006), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1015), .Y(n_1029) );
INVx1_ASAP7_75t_SL g1030 ( .A(n_1013), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1015), .Y(n_1031) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_993), .B(n_962), .Y(n_1032) );
AOI221xp5_ASAP7_75t_L g1033 ( .A1(n_1023), .A2(n_1009), .B1(n_996), .B2(n_1016), .C(n_1012), .Y(n_1033) );
AOI322xp5_ASAP7_75t_L g1034 ( .A1(n_1030), .A2(n_999), .A3(n_1002), .B1(n_1007), .B2(n_1009), .C1(n_996), .C2(n_1016), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_1027), .B(n_981), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1026), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_1028), .B(n_964), .Y(n_1037) );
AOI221xp5_ASAP7_75t_L g1038 ( .A1(n_1024), .A2(n_1003), .B1(n_1017), .B2(n_1004), .C(n_1019), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_1028), .B(n_964), .Y(n_1039) );
AOI221xp5_ASAP7_75t_L g1040 ( .A1(n_1020), .A2(n_1019), .B1(n_965), .B2(n_971), .C(n_970), .Y(n_1040) );
OAI321xp33_ASAP7_75t_L g1041 ( .A1(n_1022), .A2(n_938), .A3(n_939), .B1(n_931), .B2(n_924), .C(n_926), .Y(n_1041) );
AOI22xp5_ASAP7_75t_L g1042 ( .A1(n_1025), .A2(n_979), .B1(n_967), .B2(n_985), .Y(n_1042) );
AOI221xp5_ASAP7_75t_SL g1043 ( .A1(n_1032), .A2(n_979), .B1(n_984), .B2(n_985), .C(n_987), .Y(n_1043) );
AOI21xp5_ASAP7_75t_L g1044 ( .A1(n_1029), .A2(n_1031), .B(n_978), .Y(n_1044) );
AOI21xp5_ASAP7_75t_L g1045 ( .A1(n_1021), .A2(n_972), .B(n_970), .Y(n_1045) );
AOI221xp5_ASAP7_75t_L g1046 ( .A1(n_1023), .A2(n_965), .B1(n_971), .B2(n_987), .C(n_1010), .Y(n_1046) );
AOI221xp5_ASAP7_75t_L g1047 ( .A1(n_1033), .A2(n_1046), .B1(n_1045), .B2(n_1043), .C(n_1041), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_1034), .B(n_1036), .Y(n_1048) );
NAND4xp25_ASAP7_75t_L g1049 ( .A(n_1042), .B(n_1038), .C(n_1040), .D(n_907), .Y(n_1049) );
NOR2xp33_ASAP7_75t_L g1050 ( .A(n_1039), .B(n_1037), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_1050), .B(n_1035), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1048), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_1047), .B(n_1044), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1049), .Y(n_1054) );
AND2x4_ASAP7_75t_L g1055 ( .A(n_1054), .B(n_984), .Y(n_1055) );
INVx2_ASAP7_75t_L g1056 ( .A(n_1053), .Y(n_1056) );
AND2x4_ASAP7_75t_L g1057 ( .A(n_1051), .B(n_991), .Y(n_1057) );
NOR4xp25_ASAP7_75t_L g1058 ( .A(n_1052), .B(n_1001), .C(n_997), .D(n_891), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1056), .Y(n_1059) );
HB1xp67_ASAP7_75t_L g1060 ( .A(n_1055), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1057), .Y(n_1061) );
AOI211x1_ASAP7_75t_L g1062 ( .A1(n_1059), .A2(n_1058), .B(n_881), .C(n_888), .Y(n_1062) );
BUFx3_ASAP7_75t_L g1063 ( .A(n_1061), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_1063), .B(n_1060), .Y(n_1064) );
OR2x6_ASAP7_75t_L g1065 ( .A(n_1064), .B(n_1062), .Y(n_1065) );
XNOR2x1_ASAP7_75t_L g1066 ( .A(n_1065), .B(n_859), .Y(n_1066) );
HB1xp67_ASAP7_75t_L g1067 ( .A(n_1066), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_1067), .A2(n_928), .B1(n_1014), .B2(n_1008), .Y(n_1068) );
endmodule