module real_aes_6467_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_728;
wire n_735;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g724 ( .A(n_0), .Y(n_724) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_1), .A2(n_132), .B(n_136), .C(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g185 ( .A(n_2), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_3), .A2(n_127), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_4), .B(n_149), .Y(n_466) );
AOI21xp33_ASAP7_75t_L g153 ( .A1(n_5), .A2(n_127), .B(n_154), .Y(n_153) );
AND2x6_ASAP7_75t_L g132 ( .A(n_6), .B(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_7), .A2(n_235), .B(n_236), .Y(n_234) );
INVx1_ASAP7_75t_L g522 ( .A(n_8), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_9), .B(n_40), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_10), .B(n_158), .Y(n_501) );
INVx1_ASAP7_75t_L g160 ( .A(n_11), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_12), .B(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g125 ( .A(n_13), .Y(n_125) );
INVx1_ASAP7_75t_L g241 ( .A(n_14), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_15), .A2(n_144), .B(n_242), .C(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_16), .B(n_149), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_17), .B(n_141), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_18), .B(n_127), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_19), .B(n_550), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_20), .A2(n_168), .B(n_227), .C(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_21), .B(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_22), .B(n_158), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_23), .A2(n_239), .B(n_240), .C(n_242), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_24), .B(n_158), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g446 ( .A(n_25), .Y(n_446) );
INVx1_ASAP7_75t_L g472 ( .A(n_26), .Y(n_472) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_27), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_28), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_29), .B(n_158), .Y(n_187) );
INVx1_ASAP7_75t_L g547 ( .A(n_30), .Y(n_547) );
INVx1_ASAP7_75t_L g174 ( .A(n_31), .Y(n_174) );
OAI22xp5_ASAP7_75t_SL g754 ( .A1(n_32), .A2(n_91), .B1(n_755), .B2(n_756), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_32), .Y(n_756) );
INVx2_ASAP7_75t_L g130 ( .A(n_33), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_34), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_35), .A2(n_145), .B(n_227), .C(n_464), .Y(n_463) );
INVxp67_ASAP7_75t_L g548 ( .A(n_36), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_37), .A2(n_132), .B(n_136), .C(n_199), .Y(n_198) );
CKINVDCx14_ASAP7_75t_R g462 ( .A(n_38), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_39), .A2(n_136), .B(n_471), .C(n_476), .Y(n_470) );
INVx1_ASAP7_75t_L g172 ( .A(n_41), .Y(n_172) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_42), .A2(n_49), .B1(n_751), .B2(n_752), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_42), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_43), .A2(n_63), .B1(n_719), .B2(n_720), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_43), .Y(n_720) );
OAI22xp5_ASAP7_75t_SL g716 ( .A1(n_44), .A2(n_717), .B1(n_718), .B2(n_721), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_44), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_45), .A2(n_157), .B(n_203), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_46), .B(n_158), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_47), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_48), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_49), .Y(n_751) );
INVx1_ASAP7_75t_L g487 ( .A(n_50), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_51), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_52), .B(n_127), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_53), .A2(n_136), .B1(n_168), .B2(n_170), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g207 ( .A(n_54), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_55), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g156 ( .A1(n_56), .A2(n_145), .B(n_157), .C(n_159), .Y(n_156) );
CKINVDCx14_ASAP7_75t_R g519 ( .A(n_57), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g217 ( .A(n_58), .Y(n_217) );
INVx1_ASAP7_75t_L g155 ( .A(n_59), .Y(n_155) );
INVx1_ASAP7_75t_L g133 ( .A(n_60), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_61), .Y(n_729) );
INVx1_ASAP7_75t_L g124 ( .A(n_62), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_63), .Y(n_719) );
INVx1_ASAP7_75t_SL g465 ( .A(n_64), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_65), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_66), .B(n_149), .Y(n_491) );
INVx1_ASAP7_75t_L g449 ( .A(n_67), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_68), .Y(n_760) );
A2O1A1Ixp33_ASAP7_75t_SL g140 ( .A1(n_69), .A2(n_141), .B(n_142), .C(n_145), .Y(n_140) );
INVxp67_ASAP7_75t_L g143 ( .A(n_70), .Y(n_143) );
INVx1_ASAP7_75t_L g735 ( .A(n_71), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_72), .A2(n_127), .B(n_518), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_73), .A2(n_715), .B1(n_716), .B2(n_722), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_73), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_74), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_75), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_76), .A2(n_127), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g210 ( .A(n_77), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_78), .A2(n_235), .B(n_543), .Y(n_542) );
CKINVDCx16_ASAP7_75t_R g469 ( .A(n_79), .Y(n_469) );
INVx1_ASAP7_75t_L g507 ( .A(n_80), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_81), .A2(n_132), .B(n_136), .C(n_212), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_82), .A2(n_127), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g510 ( .A(n_83), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_84), .B(n_186), .Y(n_200) );
INVx2_ASAP7_75t_L g122 ( .A(n_85), .Y(n_122) );
INVx1_ASAP7_75t_L g500 ( .A(n_86), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_87), .B(n_141), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_88), .A2(n_132), .B(n_136), .C(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g109 ( .A(n_89), .Y(n_109) );
OR2x2_ASAP7_75t_L g739 ( .A(n_89), .B(n_728), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_90), .A2(n_136), .B(n_448), .C(n_452), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g103 ( .A1(n_91), .A2(n_104), .B1(n_730), .B2(n_740), .C(n_744), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_91), .B(n_162), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_91), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_92), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_93), .A2(n_132), .B(n_136), .C(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_94), .Y(n_231) );
INVx1_ASAP7_75t_L g139 ( .A(n_95), .Y(n_139) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_96), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_97), .B(n_186), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_98), .B(n_120), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_99), .B(n_120), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_100), .A2(n_127), .B(n_134), .Y(n_126) );
INVx2_ASAP7_75t_L g490 ( .A(n_101), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_102), .B(n_735), .Y(n_734) );
OAI22xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_723), .B1(n_726), .B2(n_729), .Y(n_104) );
XOR2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_714), .Y(n_105) );
OAI22xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_110), .B1(n_436), .B2(n_437), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g436 ( .A(n_109), .Y(n_436) );
NOR2x2_ASAP7_75t_L g727 ( .A(n_109), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx3_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND4x1_ASAP7_75t_L g112 ( .A(n_113), .B(n_354), .C(n_401), .D(n_421), .Y(n_112) );
NOR3xp33_ASAP7_75t_SL g113 ( .A(n_114), .B(n_284), .C(n_309), .Y(n_113) );
OAI211xp5_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_192), .B(n_244), .C(n_274), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_163), .Y(n_116) );
INVx3_ASAP7_75t_SL g326 ( .A(n_117), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_117), .B(n_257), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_117), .B(n_179), .Y(n_407) );
AND2x2_ASAP7_75t_L g430 ( .A(n_117), .B(n_296), .Y(n_430) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_151), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g248 ( .A(n_119), .B(n_152), .Y(n_248) );
INVx3_ASAP7_75t_L g261 ( .A(n_119), .Y(n_261) );
AND2x2_ASAP7_75t_L g266 ( .A(n_119), .B(n_151), .Y(n_266) );
OR2x2_ASAP7_75t_L g317 ( .A(n_119), .B(n_258), .Y(n_317) );
BUFx2_ASAP7_75t_L g337 ( .A(n_119), .Y(n_337) );
AND2x2_ASAP7_75t_L g347 ( .A(n_119), .B(n_258), .Y(n_347) );
AND2x2_ASAP7_75t_L g353 ( .A(n_119), .B(n_164), .Y(n_353) );
OA21x2_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_126), .B(n_148), .Y(n_119) );
INVx4_ASAP7_75t_L g150 ( .A(n_120), .Y(n_150) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_120), .Y(n_459) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g165 ( .A(n_121), .Y(n_165) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
AND2x2_ASAP7_75t_SL g162 ( .A(n_122), .B(n_123), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
BUFx2_ASAP7_75t_L g235 ( .A(n_127), .Y(n_235) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_132), .Y(n_127) );
NAND2x1p5_ASAP7_75t_L g176 ( .A(n_128), .B(n_132), .Y(n_176) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
INVx1_ASAP7_75t_L g475 ( .A(n_129), .Y(n_475) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g137 ( .A(n_130), .Y(n_137) );
INVx1_ASAP7_75t_L g169 ( .A(n_130), .Y(n_169) );
INVx1_ASAP7_75t_L g138 ( .A(n_131), .Y(n_138) );
INVx1_ASAP7_75t_L g141 ( .A(n_131), .Y(n_141) );
INVx3_ASAP7_75t_L g144 ( .A(n_131), .Y(n_144) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_131), .Y(n_158) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_131), .Y(n_171) );
INVx4_ASAP7_75t_SL g147 ( .A(n_132), .Y(n_147) );
BUFx3_ASAP7_75t_L g476 ( .A(n_132), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_139), .B(n_140), .C(n_147), .Y(n_134) );
O2A1O1Ixp33_ASAP7_75t_L g154 ( .A1(n_135), .A2(n_147), .B(n_155), .C(n_156), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_135), .A2(n_147), .B(n_237), .C(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_135), .A2(n_147), .B(n_462), .C(n_463), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_SL g486 ( .A1(n_135), .A2(n_147), .B(n_487), .C(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_SL g506 ( .A1(n_135), .A2(n_147), .B(n_507), .C(n_508), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_SL g518 ( .A1(n_135), .A2(n_147), .B(n_519), .C(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_SL g543 ( .A1(n_135), .A2(n_147), .B(n_544), .C(n_545), .Y(n_543) );
INVx5_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_137), .Y(n_146) );
BUFx3_ASAP7_75t_L g204 ( .A(n_137), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_144), .B(n_160), .Y(n_159) );
INVx5_ASAP7_75t_L g186 ( .A(n_144), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_144), .B(n_522), .Y(n_521) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_146), .Y(n_228) );
OAI22xp33_ASAP7_75t_L g166 ( .A1(n_147), .A2(n_167), .B1(n_175), .B2(n_176), .Y(n_166) );
INVx1_ASAP7_75t_L g452 ( .A(n_147), .Y(n_452) );
OA21x2_ASAP7_75t_L g152 ( .A1(n_149), .A2(n_153), .B(n_161), .Y(n_152) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_SL g206 ( .A(n_150), .B(n_207), .Y(n_206) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_150), .A2(n_445), .B(n_453), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_150), .B(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_150), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_SL g151 ( .A(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_152), .B(n_258), .Y(n_272) );
INVx2_ASAP7_75t_L g282 ( .A(n_152), .Y(n_282) );
AND2x2_ASAP7_75t_L g295 ( .A(n_152), .B(n_261), .Y(n_295) );
OR2x2_ASAP7_75t_L g306 ( .A(n_152), .B(n_258), .Y(n_306) );
AND2x2_ASAP7_75t_SL g352 ( .A(n_152), .B(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g364 ( .A(n_152), .Y(n_364) );
AND2x2_ASAP7_75t_L g410 ( .A(n_152), .B(n_164), .Y(n_410) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx4_ASAP7_75t_L g227 ( .A(n_158), .Y(n_227) );
INVx1_ASAP7_75t_L g191 ( .A(n_162), .Y(n_191) );
INVx2_ASAP7_75t_L g221 ( .A(n_162), .Y(n_221) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_162), .A2(n_234), .B(n_243), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_162), .A2(n_176), .B(n_469), .C(n_470), .Y(n_468) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_162), .A2(n_517), .B(n_523), .Y(n_516) );
INVx3_ASAP7_75t_SL g283 ( .A(n_163), .Y(n_283) );
OR2x2_ASAP7_75t_L g336 ( .A(n_163), .B(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_179), .Y(n_163) );
INVx3_ASAP7_75t_L g258 ( .A(n_164), .Y(n_258) );
AND2x2_ASAP7_75t_L g325 ( .A(n_164), .B(n_180), .Y(n_325) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_164), .Y(n_393) );
AOI33xp33_ASAP7_75t_L g397 ( .A1(n_164), .A2(n_326), .A3(n_333), .B1(n_342), .B2(n_398), .B3(n_399), .Y(n_397) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_177), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_165), .B(n_178), .Y(n_177) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_165), .A2(n_181), .B(n_189), .Y(n_180) );
INVx2_ASAP7_75t_L g205 ( .A(n_165), .Y(n_205) );
INVx2_ASAP7_75t_L g188 ( .A(n_168), .Y(n_188) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OAI22xp5_ASAP7_75t_SL g170 ( .A1(n_171), .A2(n_172), .B1(n_173), .B2(n_174), .Y(n_170) );
INVx2_ASAP7_75t_L g173 ( .A(n_171), .Y(n_173) );
INVx4_ASAP7_75t_L g239 ( .A(n_171), .Y(n_239) );
INVx2_ASAP7_75t_L g450 ( .A(n_173), .Y(n_450) );
OAI21xp5_ASAP7_75t_L g181 ( .A1(n_176), .A2(n_182), .B(n_183), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_176), .A2(n_210), .B(n_211), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_176), .A2(n_446), .B(n_447), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_176), .A2(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g246 ( .A(n_179), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_179), .B(n_261), .Y(n_260) );
NOR3xp33_ASAP7_75t_L g320 ( .A(n_179), .B(n_321), .C(n_323), .Y(n_320) );
AND2x2_ASAP7_75t_L g346 ( .A(n_179), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_179), .B(n_353), .Y(n_356) );
AND2x2_ASAP7_75t_L g409 ( .A(n_179), .B(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx3_ASAP7_75t_L g265 ( .A(n_180), .Y(n_265) );
OR2x2_ASAP7_75t_L g359 ( .A(n_180), .B(n_258), .Y(n_359) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .C(n_188), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_186), .A2(n_472), .B(n_473), .C(n_474), .Y(n_471) );
OAI22xp33_ASAP7_75t_L g546 ( .A1(n_186), .A2(n_239), .B1(n_547), .B2(n_548), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_191), .B(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_191), .B(n_231), .Y(n_230) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_191), .A2(n_496), .B(n_502), .Y(n_495) );
OR2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_218), .Y(n_192) );
AOI32xp33_ASAP7_75t_L g310 ( .A1(n_193), .A2(n_311), .A3(n_313), .B1(n_315), .B2(n_318), .Y(n_310) );
NOR2xp67_ASAP7_75t_L g383 ( .A(n_193), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g413 ( .A(n_193), .Y(n_413) );
INVx4_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g345 ( .A(n_194), .B(n_329), .Y(n_345) );
AND2x2_ASAP7_75t_L g365 ( .A(n_194), .B(n_291), .Y(n_365) );
AND2x2_ASAP7_75t_L g433 ( .A(n_194), .B(n_351), .Y(n_433) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_208), .Y(n_194) );
INVx3_ASAP7_75t_L g254 ( .A(n_195), .Y(n_254) );
AND2x2_ASAP7_75t_L g268 ( .A(n_195), .B(n_252), .Y(n_268) );
OR2x2_ASAP7_75t_L g273 ( .A(n_195), .B(n_251), .Y(n_273) );
INVx1_ASAP7_75t_L g280 ( .A(n_195), .Y(n_280) );
AND2x2_ASAP7_75t_L g288 ( .A(n_195), .B(n_262), .Y(n_288) );
AND2x2_ASAP7_75t_L g290 ( .A(n_195), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_195), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g343 ( .A(n_195), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_195), .B(n_428), .Y(n_427) );
OR2x6_ASAP7_75t_L g195 ( .A(n_196), .B(n_206), .Y(n_195) );
AOI21xp5_ASAP7_75t_SL g196 ( .A1(n_197), .A2(n_198), .B(n_205), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_202), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_202), .A2(n_213), .B(n_214), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g448 ( .A1(n_202), .A2(n_449), .B(n_450), .C(n_451), .Y(n_448) );
O2A1O1Ixp5_ASAP7_75t_L g499 ( .A1(n_202), .A2(n_450), .B(n_500), .C(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g242 ( .A(n_204), .Y(n_242) );
INVx1_ASAP7_75t_L g215 ( .A(n_205), .Y(n_215) );
INVx2_ASAP7_75t_L g252 ( .A(n_208), .Y(n_252) );
AND2x2_ASAP7_75t_L g298 ( .A(n_208), .B(n_219), .Y(n_298) );
AND2x2_ASAP7_75t_L g308 ( .A(n_208), .B(n_233), .Y(n_308) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_215), .B(n_216), .Y(n_208) );
INVx1_ASAP7_75t_L g541 ( .A(n_215), .Y(n_541) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_215), .A2(n_558), .B(n_559), .Y(n_557) );
INVx2_ASAP7_75t_L g428 ( .A(n_218), .Y(n_428) );
OR2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_232), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_219), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g269 ( .A(n_219), .Y(n_269) );
AND2x2_ASAP7_75t_L g313 ( .A(n_219), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g329 ( .A(n_219), .B(n_292), .Y(n_329) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g277 ( .A(n_220), .Y(n_277) );
AND2x2_ASAP7_75t_L g291 ( .A(n_220), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g342 ( .A(n_220), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_220), .B(n_252), .Y(n_374) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_230), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_221), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g550 ( .A(n_221), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_229), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_228), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_227), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g253 ( .A(n_232), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g314 ( .A(n_232), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_232), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g351 ( .A(n_232), .Y(n_351) );
INVx1_ASAP7_75t_L g384 ( .A(n_232), .Y(n_384) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g262 ( .A(n_233), .B(n_252), .Y(n_262) );
INVx1_ASAP7_75t_L g292 ( .A(n_233), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_239), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_239), .B(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_239), .B(n_510), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_249), .B1(n_255), .B2(n_262), .C(n_263), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_246), .B(n_266), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_246), .B(n_329), .Y(n_406) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_248), .B(n_296), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_248), .B(n_257), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_248), .B(n_271), .Y(n_400) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_253), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g322 ( .A(n_252), .Y(n_322) );
AND2x2_ASAP7_75t_L g297 ( .A(n_253), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g375 ( .A(n_253), .Y(n_375) );
AND2x2_ASAP7_75t_L g307 ( .A(n_254), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_254), .B(n_277), .Y(n_323) );
AND2x2_ASAP7_75t_L g387 ( .A(n_254), .B(n_313), .Y(n_387) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
BUFx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g296 ( .A(n_258), .B(n_265), .Y(n_296) );
AND2x2_ASAP7_75t_L g392 ( .A(n_259), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_261), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_262), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_262), .B(n_269), .Y(n_357) );
AND2x2_ASAP7_75t_L g377 ( .A(n_262), .B(n_277), .Y(n_377) );
AND2x2_ASAP7_75t_L g398 ( .A(n_262), .B(n_342), .Y(n_398) );
OAI32xp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_267), .A3(n_269), .B1(n_270), .B2(n_273), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_SL g271 ( .A(n_265), .Y(n_271) );
NAND2x1_ASAP7_75t_L g312 ( .A(n_265), .B(n_295), .Y(n_312) );
OR2x2_ASAP7_75t_L g316 ( .A(n_265), .B(n_317), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_265), .B(n_364), .Y(n_417) );
INVx1_ASAP7_75t_L g285 ( .A(n_266), .Y(n_285) );
OAI221xp5_ASAP7_75t_SL g403 ( .A1(n_267), .A2(n_358), .B1(n_404), .B2(n_407), .C(n_408), .Y(n_403) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g275 ( .A(n_268), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g318 ( .A(n_268), .B(n_291), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_268), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g396 ( .A(n_268), .B(n_329), .Y(n_396) );
INVxp67_ASAP7_75t_L g332 ( .A(n_269), .Y(n_332) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
AND2x2_ASAP7_75t_L g402 ( .A(n_271), .B(n_389), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_271), .B(n_352), .Y(n_425) );
INVx1_ASAP7_75t_L g300 ( .A(n_273), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_273), .B(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g418 ( .A(n_273), .B(n_419), .Y(n_418) );
OAI21xp5_ASAP7_75t_SL g274 ( .A1(n_275), .A2(n_278), .B(n_281), .Y(n_274) );
AND2x2_ASAP7_75t_L g287 ( .A(n_276), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g371 ( .A(n_280), .B(n_291), .Y(n_371) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g389 ( .A(n_282), .B(n_347), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_282), .B(n_346), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_283), .B(n_295), .Y(n_369) );
OAI211xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_286), .B(n_289), .C(n_299), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g319 ( .A1(n_285), .A2(n_320), .B1(n_324), .B2(n_327), .C(n_330), .Y(n_319) );
AOI31xp33_ASAP7_75t_L g414 ( .A1(n_285), .A2(n_415), .A3(n_416), .B(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_293), .B1(n_295), .B2(n_297), .Y(n_289) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g415 ( .A(n_295), .Y(n_415) );
INVx1_ASAP7_75t_L g378 ( .A(n_296), .Y(n_378) );
O2A1O1Ixp33_ASAP7_75t_L g421 ( .A1(n_298), .A2(n_422), .B(n_424), .C(n_426), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B1(n_303), .B2(n_307), .Y(n_299) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_304), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI221xp5_ASAP7_75t_SL g394 ( .A1(n_306), .A2(n_340), .B1(n_359), .B2(n_395), .C(n_397), .Y(n_394) );
INVx1_ASAP7_75t_L g390 ( .A(n_307), .Y(n_390) );
INVx1_ASAP7_75t_L g344 ( .A(n_308), .Y(n_344) );
NAND3xp33_ASAP7_75t_SL g309 ( .A(n_310), .B(n_319), .C(n_334), .Y(n_309) );
OAI21xp33_ASAP7_75t_L g360 ( .A1(n_311), .A2(n_361), .B(n_365), .Y(n_360) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_313), .B(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g420 ( .A(n_314), .Y(n_420) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g358 ( .A(n_321), .B(n_341), .Y(n_358) );
INVx1_ASAP7_75t_L g333 ( .A(n_322), .Y(n_333) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g331 ( .A(n_325), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_325), .B(n_363), .Y(n_362) );
NOR4xp25_ASAP7_75t_L g330 ( .A(n_326), .B(n_331), .C(n_332), .D(n_333), .Y(n_330) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI222xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_339), .B1(n_345), .B2(n_346), .C1(n_348), .C2(n_352), .Y(n_334) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx1_ASAP7_75t_L g432 ( .A(n_336), .Y(n_432) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_344), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_348), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI21xp5_ASAP7_75t_SL g408 ( .A1(n_353), .A2(n_409), .B(n_411), .Y(n_408) );
NOR4xp25_ASAP7_75t_L g354 ( .A(n_355), .B(n_366), .C(n_379), .D(n_394), .Y(n_354) );
OAI221xp5_ASAP7_75t_SL g355 ( .A1(n_356), .A2(n_357), .B1(n_358), .B2(n_359), .C(n_360), .Y(n_355) );
INVx1_ASAP7_75t_L g435 ( .A(n_356), .Y(n_435) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_363), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
OAI222xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_370), .B1(n_372), .B2(n_373), .C1(n_376), .C2(n_378), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AOI211xp5_ASAP7_75t_L g401 ( .A1(n_371), .A2(n_402), .B(n_403), .C(n_414), .Y(n_401) );
OR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
OAI222xp33_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_385), .B1(n_386), .B2(n_388), .C1(n_390), .C2(n_391), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_396), .A2(n_399), .B1(n_432), .B2(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI211xp5_ASAP7_75t_SL g426 ( .A1(n_427), .A2(n_429), .B(n_431), .C(n_434), .Y(n_426) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
XNOR2xp5_ASAP7_75t_L g749 ( .A(n_437), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_SL g437 ( .A(n_438), .B(n_669), .Y(n_437) );
NOR4xp25_ASAP7_75t_L g438 ( .A(n_439), .B(n_606), .C(n_640), .D(n_656), .Y(n_438) );
NAND4xp25_ASAP7_75t_SL g439 ( .A(n_440), .B(n_536), .C(n_570), .D(n_586), .Y(n_439) );
AOI222xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_479), .B1(n_512), .B2(n_524), .C1(n_529), .C2(n_535), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AOI31xp33_ASAP7_75t_L g702 ( .A1(n_442), .A2(n_703), .A3(n_704), .B(n_706), .Y(n_702) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_455), .Y(n_442) );
AND2x2_ASAP7_75t_L g677 ( .A(n_443), .B(n_457), .Y(n_677) );
BUFx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_SL g528 ( .A(n_444), .Y(n_528) );
AND2x2_ASAP7_75t_L g535 ( .A(n_444), .B(n_467), .Y(n_535) );
AND2x2_ASAP7_75t_L g591 ( .A(n_444), .B(n_458), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_455), .B(n_621), .Y(n_620) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_456), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_456), .B(n_539), .Y(n_581) );
AND2x2_ASAP7_75t_L g674 ( .A(n_456), .B(n_614), .Y(n_674) );
OAI321xp33_ASAP7_75t_L g708 ( .A1(n_456), .A2(n_528), .A3(n_681), .B1(n_709), .B2(n_711), .C(n_712), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g712 ( .A(n_456), .B(n_515), .C(n_621), .D(n_713), .Y(n_712) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_467), .Y(n_456) );
AND2x2_ASAP7_75t_L g576 ( .A(n_457), .B(n_526), .Y(n_576) );
AND2x2_ASAP7_75t_L g595 ( .A(n_457), .B(n_528), .Y(n_595) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g527 ( .A(n_458), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g551 ( .A(n_458), .B(n_467), .Y(n_551) );
AND2x2_ASAP7_75t_L g637 ( .A(n_458), .B(n_526), .Y(n_637) );
OA21x2_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B(n_466), .Y(n_458) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_459), .A2(n_485), .B(n_491), .Y(n_484) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_459), .A2(n_505), .B(n_511), .Y(n_504) );
INVx3_ASAP7_75t_SL g526 ( .A(n_467), .Y(n_526) );
AND2x2_ASAP7_75t_L g569 ( .A(n_467), .B(n_556), .Y(n_569) );
OR2x2_ASAP7_75t_L g602 ( .A(n_467), .B(n_528), .Y(n_602) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_467), .Y(n_609) );
AND2x2_ASAP7_75t_L g638 ( .A(n_467), .B(n_527), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_467), .B(n_611), .Y(n_653) );
AND2x2_ASAP7_75t_L g685 ( .A(n_467), .B(n_677), .Y(n_685) );
AND2x2_ASAP7_75t_L g694 ( .A(n_467), .B(n_540), .Y(n_694) );
OR2x6_ASAP7_75t_L g467 ( .A(n_468), .B(n_477), .Y(n_467) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_475), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_492), .Y(n_480) );
INVx1_ASAP7_75t_SL g662 ( .A(n_481), .Y(n_662) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g531 ( .A(n_482), .B(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g514 ( .A(n_483), .B(n_494), .Y(n_514) );
AND2x2_ASAP7_75t_L g598 ( .A(n_483), .B(n_516), .Y(n_598) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g568 ( .A(n_484), .B(n_504), .Y(n_568) );
OR2x2_ASAP7_75t_L g579 ( .A(n_484), .B(n_516), .Y(n_579) );
AND2x2_ASAP7_75t_L g605 ( .A(n_484), .B(n_516), .Y(n_605) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_484), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_492), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_492), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_SL g492 ( .A(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g578 ( .A(n_493), .B(n_579), .Y(n_578) );
AOI322xp5_ASAP7_75t_L g664 ( .A1(n_493), .A2(n_568), .A3(n_574), .B1(n_605), .B2(n_655), .C1(n_665), .C2(n_667), .Y(n_664) );
OR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_504), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_494), .B(n_515), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_494), .B(n_516), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_494), .B(n_532), .Y(n_585) );
AND2x2_ASAP7_75t_L g639 ( .A(n_494), .B(n_605), .Y(n_639) );
INVx1_ASAP7_75t_L g643 ( .A(n_494), .Y(n_643) );
AND2x2_ASAP7_75t_L g655 ( .A(n_494), .B(n_504), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_494), .B(n_531), .Y(n_687) );
INVx4_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g552 ( .A(n_495), .B(n_504), .Y(n_552) );
BUFx3_ASAP7_75t_L g566 ( .A(n_495), .Y(n_566) );
AND3x2_ASAP7_75t_L g648 ( .A(n_495), .B(n_628), .C(n_649), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_504), .B(n_514), .C(n_515), .Y(n_513) );
INVx1_ASAP7_75t_SL g532 ( .A(n_504), .Y(n_532) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_504), .Y(n_633) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g627 ( .A(n_514), .B(n_628), .Y(n_627) );
INVxp67_ASAP7_75t_L g634 ( .A(n_514), .Y(n_634) );
AND2x2_ASAP7_75t_L g672 ( .A(n_515), .B(n_650), .Y(n_672) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx3_ASAP7_75t_L g553 ( .A(n_516), .Y(n_553) );
AND2x2_ASAP7_75t_L g628 ( .A(n_516), .B(n_532), .Y(n_628) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
OR2x2_ASAP7_75t_L g572 ( .A(n_526), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g691 ( .A(n_526), .B(n_591), .Y(n_691) );
AND2x2_ASAP7_75t_L g705 ( .A(n_526), .B(n_528), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_527), .B(n_540), .Y(n_646) );
AND2x2_ASAP7_75t_L g693 ( .A(n_527), .B(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g556 ( .A(n_528), .B(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g573 ( .A(n_528), .B(n_540), .Y(n_573) );
INVx1_ASAP7_75t_L g583 ( .A(n_528), .Y(n_583) );
AND2x2_ASAP7_75t_L g614 ( .A(n_528), .B(n_540), .Y(n_614) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g656 ( .A1(n_530), .A2(n_657), .B1(n_661), .B2(n_663), .C(n_664), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_531), .B(n_533), .Y(n_530) );
AND2x2_ASAP7_75t_L g560 ( .A(n_531), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_534), .B(n_567), .Y(n_710) );
AOI322xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_552), .A3(n_553), .B1(n_554), .B2(n_560), .C1(n_562), .C2(n_569), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_551), .Y(n_538) );
NAND2x1p5_ASAP7_75t_L g590 ( .A(n_539), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_539), .B(n_601), .Y(n_600) );
O2A1O1Ixp33_ASAP7_75t_L g624 ( .A1(n_539), .A2(n_551), .B(n_625), .C(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_539), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_539), .B(n_595), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_539), .B(n_677), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_539), .B(n_705), .Y(n_704) );
BUFx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_540), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_540), .B(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g666 ( .A(n_540), .B(n_553), .Y(n_666) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B(n_549), .Y(n_540) );
INVx1_ASAP7_75t_L g558 ( .A(n_542), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_549), .Y(n_559) );
INVx1_ASAP7_75t_L g641 ( .A(n_551), .Y(n_641) );
OAI31xp33_ASAP7_75t_L g651 ( .A1(n_551), .A2(n_576), .A3(n_652), .B(n_654), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_551), .B(n_557), .Y(n_703) );
INVx1_ASAP7_75t_SL g564 ( .A(n_552), .Y(n_564) );
AND2x2_ASAP7_75t_L g597 ( .A(n_552), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g678 ( .A(n_552), .B(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g563 ( .A(n_553), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g588 ( .A(n_553), .Y(n_588) );
AND2x2_ASAP7_75t_L g615 ( .A(n_553), .B(n_568), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_553), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g707 ( .A(n_553), .B(n_655), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_555), .B(n_625), .Y(n_698) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g594 ( .A(n_557), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_SL g612 ( .A(n_557), .Y(n_612) );
NAND2xp33_ASAP7_75t_SL g562 ( .A(n_563), .B(n_565), .Y(n_562) );
OAI211xp5_ASAP7_75t_SL g606 ( .A1(n_564), .A2(n_607), .B(n_613), .C(n_629), .Y(n_606) );
OR2x2_ASAP7_75t_L g681 ( .A(n_564), .B(n_662), .Y(n_681) );
OR2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
CKINVDCx16_ASAP7_75t_R g618 ( .A(n_566), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_566), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g587 ( .A(n_568), .B(n_588), .Y(n_587) );
O2A1O1Ixp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_574), .B(n_577), .C(n_580), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_SL g621 ( .A(n_573), .Y(n_621) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_576), .B(n_614), .Y(n_619) );
INVx1_ASAP7_75t_L g625 ( .A(n_576), .Y(n_625) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g584 ( .A(n_579), .B(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g617 ( .A(n_579), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g679 ( .A(n_579), .Y(n_679) );
AOI21xp33_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_582), .B(n_584), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_582), .A2(n_593), .B(n_596), .Y(n_592) );
AOI211xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_589), .B(n_592), .C(n_599), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_587), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_590), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_SL g603 ( .A(n_591), .Y(n_603) );
OAI21xp5_ASAP7_75t_L g658 ( .A1(n_593), .A2(n_659), .B(n_660), .Y(n_658) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_598), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_SL g623 ( .A(n_598), .Y(n_623) );
AOI21xp33_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_603), .B(n_604), .Y(n_599) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g654 ( .A(n_605), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_611), .B(n_637), .Y(n_663) );
AND2x2_ASAP7_75t_L g676 ( .A(n_611), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g690 ( .A(n_611), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g700 ( .A(n_611), .B(n_638), .Y(n_700) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AOI211xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B(n_616), .C(n_624), .Y(n_613) );
INVx1_ASAP7_75t_L g660 ( .A(n_614), .Y(n_660) );
OAI22xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_619), .B1(n_620), .B2(n_622), .Y(n_616) );
OR2x2_ASAP7_75t_L g622 ( .A(n_618), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_618), .B(n_679), .Y(n_701) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g695 ( .A(n_628), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_635), .B1(n_638), .B2(n_639), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g713 ( .A(n_633), .Y(n_713) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g659 ( .A(n_637), .Y(n_659) );
OAI211xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_642), .B(n_644), .C(n_651), .Y(n_640) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_659), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NOR5xp2_ASAP7_75t_L g669 ( .A(n_670), .B(n_688), .C(n_696), .D(n_702), .E(n_708), .Y(n_669) );
OAI211xp5_ASAP7_75t_SL g670 ( .A1(n_671), .A2(n_673), .B(n_675), .C(n_682), .Y(n_670) );
INVxp67_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_678), .B(n_680), .Y(n_675) );
OAI21xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_685), .B(n_686), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_685), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI21xp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_692), .B(n_695), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g711 ( .A(n_691), .Y(n_711) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_699), .B(n_701), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g728 ( .A(n_723), .Y(n_728) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVx3_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
BUFx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NAND2xp33_ASAP7_75t_L g732 ( .A(n_733), .B(n_737), .Y(n_732) );
NOR2xp33_ASAP7_75t_SL g733 ( .A(n_734), .B(n_736), .Y(n_733) );
INVx1_ASAP7_75t_SL g743 ( .A(n_734), .Y(n_743) );
OA21x2_ASAP7_75t_L g741 ( .A1(n_736), .A2(n_742), .B(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g766 ( .A(n_736), .Y(n_766) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
BUFx2_ASAP7_75t_L g742 ( .A(n_739), .Y(n_742) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_739), .Y(n_746) );
INVx2_ASAP7_75t_L g762 ( .A(n_739), .Y(n_762) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g764 ( .A(n_743), .B(n_765), .Y(n_764) );
O2A1O1Ixp33_ASAP7_75t_SL g744 ( .A1(n_745), .A2(n_747), .B(n_758), .C(n_763), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
INVxp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI22xp5_ASAP7_75t_SL g748 ( .A1(n_749), .A2(n_753), .B1(n_754), .B2(n_757), .Y(n_748) );
INVx1_ASAP7_75t_L g757 ( .A(n_749), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
CKINVDCx14_ASAP7_75t_R g758 ( .A(n_759), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
CKINVDCx6p67_ASAP7_75t_R g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
endmodule