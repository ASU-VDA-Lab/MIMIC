module fake_aes_1716_n_15 (n_1, n_2, n_0, n_15);
input n_1;
input n_2;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_8;
wire n_10;
wire n_7;
INVx1_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
O2A1O1Ixp33_ASAP7_75t_SL g5 ( .A1(n_3), .A2(n_0), .B(n_1), .C(n_2), .Y(n_5) );
AOI21xp5_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_6) );
BUFx2_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
AND2x4_ASAP7_75t_L g8 ( .A(n_6), .B(n_3), .Y(n_8) );
INVx1_ASAP7_75t_SL g9 ( .A(n_8), .Y(n_9) );
OAI21xp33_ASAP7_75t_SL g10 ( .A1(n_9), .A2(n_7), .B(n_8), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
OAI211xp5_ASAP7_75t_SL g12 ( .A1(n_10), .A2(n_7), .B(n_8), .C(n_2), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_11), .B(n_8), .Y(n_13) );
AOI22x1_ASAP7_75t_L g14 ( .A1(n_12), .A2(n_11), .B1(n_0), .B2(n_1), .Y(n_14) );
AO21x2_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_13), .B(n_1), .Y(n_15) );
endmodule