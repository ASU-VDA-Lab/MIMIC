module fake_ariane_1846_n_646 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_122, n_52, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_646);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_122;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_646;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_133;
wire n_610;
wire n_205;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_139;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_143;
wire n_566;
wire n_578;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_166;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_588;
wire n_638;
wire n_136;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_616;
wire n_617;
wire n_630;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_601;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_641;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_613;
wire n_475;
wire n_135;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_544;
wire n_216;
wire n_540;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_509;
wire n_583;
wire n_306;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_292;
wire n_156;
wire n_174;
wire n_275;
wire n_132;
wire n_147;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_155;
wire n_573;
wire n_531;

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_29),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_46),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_55),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_101),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_20),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_42),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_47),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_120),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_103),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_36),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_118),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_12),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

NOR2xp67_ASAP7_75t_L g147 ( 
.A(n_73),
.B(n_8),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_82),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_53),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_99),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_31),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_8),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_33),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_131),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_76),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_115),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_94),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_10),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_123),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_17),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_59),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_9),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_0),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_28),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_125),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_74),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_54),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_129),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_11),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_89),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_92),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_127),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_14),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_5),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_106),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_77),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_100),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_108),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_27),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_25),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_93),
.Y(n_187)
);

NOR2xp67_ASAP7_75t_L g188 ( 
.A(n_22),
.B(n_7),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_111),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_105),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_L g192 ( 
.A(n_35),
.B(n_83),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_4),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_15),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_124),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_97),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_117),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_34),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_24),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_19),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_3),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_0),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_144),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_139),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_143),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_153),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_149),
.B(n_1),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_174),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_158),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

AND2x6_ASAP7_75t_L g221 ( 
.A(n_142),
.B(n_13),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_2),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_142),
.A2(n_69),
.B(n_128),
.Y(n_226)
);

OA21x2_ASAP7_75t_L g227 ( 
.A1(n_167),
.A2(n_4),
.B(n_5),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_169),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_132),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_150),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_145),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_145),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g236 ( 
.A(n_133),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_183),
.B(n_6),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_184),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_170),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_200),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_138),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_134),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_146),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_135),
.Y(n_247)
);

AND2x4_ASAP7_75t_L g248 ( 
.A(n_147),
.B(n_6),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_232),
.Y(n_249)
);

AND3x2_ASAP7_75t_L g250 ( 
.A(n_203),
.B(n_195),
.C(n_173),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_210),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_239),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_220),
.Y(n_259)
);

NOR2x1p5_ASAP7_75t_L g260 ( 
.A(n_217),
.B(n_136),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_230),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_R g262 ( 
.A(n_230),
.B(n_198),
.Y(n_262)
);

NAND2xp33_ASAP7_75t_R g263 ( 
.A(n_217),
.B(n_137),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_236),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_236),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_224),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_R g268 ( 
.A(n_247),
.B(n_197),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_209),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_209),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_245),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_245),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_202),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_202),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_211),
.B(n_177),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_246),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_231),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_R g279 ( 
.A(n_223),
.B(n_196),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_231),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_246),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_242),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_240),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_242),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_206),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_206),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_238),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_240),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_244),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_243),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_243),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_211),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_207),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_207),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_205),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_233),
.B(n_181),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_248),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_214),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_214),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_215),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_252),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_215),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_271),
.B(n_218),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_255),
.Y(n_306)
);

NOR2x1p5_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_248),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_278),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_290),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_218),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_253),
.B(n_233),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_277),
.B(n_237),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_273),
.B(n_225),
.Y(n_313)
);

NAND3xp33_ASAP7_75t_L g314 ( 
.A(n_287),
.B(n_212),
.C(n_227),
.Y(n_314)
);

INVx8_ASAP7_75t_L g315 ( 
.A(n_266),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_280),
.B(n_222),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_254),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_253),
.B(n_225),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_288),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_276),
.B(n_244),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_276),
.B(n_228),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_257),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_298),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_264),
.Y(n_325)
);

BUFx8_ASAP7_75t_L g326 ( 
.A(n_275),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_283),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_299),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_300),
.Y(n_329)
);

NAND3xp33_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_212),
.C(n_227),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_249),
.B(n_241),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_274),
.B(n_241),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_282),
.B(n_286),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_281),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_228),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_269),
.B(n_234),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_295),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_251),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_251),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_268),
.B(n_229),
.Y(n_341)
);

NAND2xp33_ASAP7_75t_L g342 ( 
.A(n_260),
.B(n_221),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_270),
.B(n_234),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_297),
.B(n_229),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_284),
.B(n_204),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_279),
.B(n_188),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_250),
.B(n_205),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_250),
.B(n_205),
.Y(n_348)
);

NOR3xp33_ASAP7_75t_L g349 ( 
.A(n_258),
.B(n_226),
.C(n_140),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_251),
.B(n_256),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_262),
.B(n_141),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_256),
.B(n_208),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_259),
.B(n_148),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_263),
.B(n_151),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_292),
.Y(n_355)
);

NOR3xp33_ASAP7_75t_L g356 ( 
.A(n_261),
.B(n_176),
.C(n_155),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_267),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_259),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_276),
.B(n_208),
.Y(n_359)
);

AOI221xp5_ASAP7_75t_L g360 ( 
.A1(n_292),
.A2(n_178),
.B1(n_156),
.B2(n_159),
.C(n_160),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_271),
.B(n_152),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_L g362 ( 
.A(n_271),
.B(n_221),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_271),
.B(n_162),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_289),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_293),
.B(n_221),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_275),
.A2(n_227),
.B1(n_221),
.B2(n_192),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_271),
.B(n_163),
.Y(n_367)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_319),
.Y(n_368)
);

OR2x6_ASAP7_75t_SL g369 ( 
.A(n_355),
.B(n_166),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_309),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_333),
.B(n_171),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_305),
.B(n_180),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_324),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_331),
.B(n_185),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_321),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_334),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_310),
.B(n_186),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_319),
.B(n_187),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_314),
.A2(n_221),
.B1(n_189),
.B2(n_213),
.Y(n_379)
);

NOR3xp33_ASAP7_75t_SL g380 ( 
.A(n_360),
.B(n_7),
.C(n_9),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_315),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_358),
.B(n_208),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_328),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_329),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_361),
.B(n_16),
.Y(n_385)
);

INVxp33_ASAP7_75t_L g386 ( 
.A(n_353),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_328),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_313),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_332),
.B(n_208),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_339),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_326),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_344),
.A2(n_219),
.B1(n_213),
.B2(n_23),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_323),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g396 ( 
.A(n_341),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_363),
.B(n_18),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_367),
.B(n_21),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_307),
.B(n_26),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_326),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_318),
.B(n_311),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_359),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_R g403 ( 
.A(n_315),
.B(n_30),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_301),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_364),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_340),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_320),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_R g408 ( 
.A(n_338),
.B(n_32),
.Y(n_408)
);

NAND2x1p5_ASAP7_75t_L g409 ( 
.A(n_304),
.B(n_219),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_357),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_325),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_312),
.B(n_219),
.Y(n_412)
);

NOR3xp33_ASAP7_75t_SL g413 ( 
.A(n_346),
.B(n_37),
.C(n_38),
.Y(n_413)
);

NOR3xp33_ASAP7_75t_L g414 ( 
.A(n_356),
.B(n_39),
.C(n_40),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_327),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g416 ( 
.A1(n_314),
.A2(n_219),
.B1(n_213),
.B2(n_44),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_302),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_322),
.Y(n_418)
);

NAND3xp33_ASAP7_75t_SL g419 ( 
.A(n_345),
.B(n_41),
.C(n_43),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_350),
.B(n_45),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_337),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_347),
.Y(n_422)
);

NOR2xp67_ASAP7_75t_L g423 ( 
.A(n_303),
.B(n_48),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_306),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_348),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_303),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_336),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_335),
.B(n_354),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_308),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_352),
.B(n_213),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_317),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_365),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_373),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_384),
.Y(n_434)
);

NOR3xp33_ASAP7_75t_L g435 ( 
.A(n_389),
.B(n_316),
.C(n_351),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_432),
.A2(n_342),
.B(n_431),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_388),
.A2(n_362),
.B(n_365),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_377),
.A2(n_349),
.B(n_330),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_421),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_386),
.B(n_366),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_368),
.B(n_317),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_L g442 ( 
.A(n_368),
.B(n_317),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_381),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_330),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_402),
.A2(n_317),
.B(n_50),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_410),
.A2(n_387),
.B1(n_399),
.B2(n_393),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_370),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_317),
.Y(n_448)
);

A2O1A1Ixp33_ASAP7_75t_L g449 ( 
.A1(n_385),
.A2(n_49),
.B(n_51),
.C(n_52),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_397),
.A2(n_56),
.B(n_57),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_383),
.Y(n_451)
);

O2A1O1Ixp33_ASAP7_75t_L g452 ( 
.A1(n_380),
.A2(n_58),
.B(n_60),
.C(n_61),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_376),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_398),
.A2(n_62),
.B(n_63),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_396),
.B(n_64),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_375),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_395),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_368),
.B(n_65),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_418),
.A2(n_66),
.B(n_67),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_372),
.A2(n_68),
.B(n_70),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_392),
.B(n_71),
.Y(n_461)
);

BUFx2_ASAP7_75t_SL g462 ( 
.A(n_400),
.Y(n_462)
);

AOI22x1_ASAP7_75t_L g463 ( 
.A1(n_383),
.A2(n_72),
.B1(n_75),
.B2(n_79),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_383),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_407),
.B(n_80),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_391),
.Y(n_466)
);

O2A1O1Ixp33_ASAP7_75t_L g467 ( 
.A1(n_378),
.A2(n_81),
.B(n_85),
.C(n_87),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_417),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_424),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_429),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_422),
.B(n_425),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_428),
.A2(n_88),
.B(n_90),
.Y(n_472)
);

NOR3xp33_ASAP7_75t_SL g473 ( 
.A(n_371),
.B(n_91),
.C(n_96),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_404),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_411),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_422),
.B(n_423),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_436),
.A2(n_416),
.B(n_379),
.Y(n_477)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_451),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_440),
.B(n_422),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_453),
.B(n_382),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_433),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_475),
.Y(n_482)
);

NAND2x1p5_ASAP7_75t_L g483 ( 
.A(n_451),
.B(n_464),
.Y(n_483)
);

AO21x2_ASAP7_75t_L g484 ( 
.A1(n_438),
.A2(n_390),
.B(n_394),
.Y(n_484)
);

OR3x4_ASAP7_75t_SL g485 ( 
.A(n_446),
.B(n_369),
.C(n_403),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_434),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_436),
.A2(n_409),
.B(n_430),
.Y(n_487)
);

NAND2x1p5_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_399),
.Y(n_488)
);

AO21x2_ASAP7_75t_L g489 ( 
.A1(n_437),
.A2(n_412),
.B(n_419),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_474),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_443),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_442),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_444),
.B(n_420),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_443),
.Y(n_494)
);

AO21x2_ASAP7_75t_L g495 ( 
.A1(n_437),
.A2(n_374),
.B(n_420),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_445),
.A2(n_405),
.B(n_401),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_470),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_472),
.A2(n_406),
.B(n_391),
.Y(n_498)
);

BUFx6f_ASAP7_75t_SL g499 ( 
.A(n_439),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_447),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_466),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_466),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_471),
.B(n_415),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_472),
.A2(n_465),
.B(n_448),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_SL g505 ( 
.A1(n_455),
.A2(n_408),
.B1(n_415),
.B2(n_406),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_471),
.B(n_415),
.Y(n_506)
);

CKINVDCx8_ASAP7_75t_R g507 ( 
.A(n_462),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_481),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_494),
.Y(n_509)
);

BUFx8_ASAP7_75t_SL g510 ( 
.A(n_499),
.Y(n_510)
);

AO21x1_ASAP7_75t_L g511 ( 
.A1(n_504),
.A2(n_477),
.B(n_493),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_480),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_479),
.B(n_456),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_507),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_486),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_491),
.Y(n_516)
);

AOI21x1_ASAP7_75t_L g517 ( 
.A1(n_504),
.A2(n_476),
.B(n_450),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_493),
.A2(n_457),
.B1(n_414),
.B2(n_469),
.Y(n_518)
);

OA21x2_ASAP7_75t_L g519 ( 
.A1(n_477),
.A2(n_460),
.B(n_449),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_482),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_479),
.B(n_435),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_503),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_490),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_503),
.B(n_506),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_SL g525 ( 
.A(n_499),
.B(n_473),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_500),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_498),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_492),
.A2(n_505),
.B1(n_488),
.B2(n_506),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_492),
.A2(n_452),
.B1(n_441),
.B2(n_476),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_497),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_483),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_496),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_495),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_478),
.B(n_461),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_512),
.B(n_488),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_508),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_513),
.A2(n_505),
.B1(n_468),
.B2(n_495),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_510),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_522),
.B(n_478),
.Y(n_539)
);

OAI22xp33_ASAP7_75t_L g540 ( 
.A1(n_521),
.A2(n_485),
.B1(n_478),
.B2(n_501),
.Y(n_540)
);

AO31x2_ASAP7_75t_L g541 ( 
.A1(n_511),
.A2(n_454),
.A3(n_459),
.B(n_484),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_509),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_478),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_SL g544 ( 
.A1(n_528),
.A2(n_485),
.B1(n_489),
.B2(n_484),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_516),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_515),
.B(n_502),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_R g547 ( 
.A(n_514),
.B(n_502),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_520),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_523),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_520),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_526),
.Y(n_551)
);

CKINVDCx16_ASAP7_75t_R g552 ( 
.A(n_514),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_513),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_524),
.B(n_501),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_524),
.B(n_530),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_531),
.B(n_502),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_534),
.B(n_502),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_R g558 ( 
.A(n_525),
.B(n_501),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_533),
.Y(n_559)
);

AO32x2_ASAP7_75t_L g560 ( 
.A1(n_529),
.A2(n_489),
.A3(n_487),
.B1(n_413),
.B2(n_467),
.Y(n_560)
);

O2A1O1Ixp33_ASAP7_75t_SL g561 ( 
.A1(n_525),
.A2(n_458),
.B(n_463),
.C(n_483),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_533),
.Y(n_562)
);

CKINVDCx16_ASAP7_75t_R g563 ( 
.A(n_534),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_518),
.A2(n_501),
.B(n_406),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_519),
.A2(n_391),
.B(n_102),
.Y(n_565)
);

NAND4xp25_ASAP7_75t_L g566 ( 
.A(n_545),
.B(n_536),
.C(n_549),
.D(n_544),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_562),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_555),
.B(n_534),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_563),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_551),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_L g571 ( 
.A1(n_552),
.A2(n_519),
.B1(n_517),
.B2(n_510),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_559),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_553),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_550),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_564),
.B(n_518),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_535),
.B(n_519),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_548),
.Y(n_577)
);

OR2x2_ASAP7_75t_SL g578 ( 
.A(n_542),
.B(n_546),
.Y(n_578)
);

AO21x2_ASAP7_75t_L g579 ( 
.A1(n_565),
.A2(n_527),
.B(n_532),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_564),
.B(n_527),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_547),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_554),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_554),
.B(n_532),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_540),
.A2(n_98),
.B1(n_104),
.B2(n_107),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_539),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_557),
.B(n_109),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_556),
.B(n_110),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_539),
.B(n_112),
.Y(n_588)
);

INVxp67_ASAP7_75t_SL g589 ( 
.A(n_583),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_570),
.Y(n_590)
);

INVxp67_ASAP7_75t_SL g591 ( 
.A(n_571),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_582),
.B(n_537),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_574),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_573),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_574),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_568),
.B(n_538),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_569),
.B(n_543),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_569),
.B(n_543),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_575),
.B(n_558),
.Y(n_599)
);

BUFx2_ASAP7_75t_SL g600 ( 
.A(n_581),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_576),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_572),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_572),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_596),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_590),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_601),
.B(n_578),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_603),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_601),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_600),
.B(n_585),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_589),
.B(n_571),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_598),
.B(n_585),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_605),
.Y(n_612)
);

INVxp67_ASAP7_75t_SL g613 ( 
.A(n_608),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_608),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_SL g615 ( 
.A1(n_610),
.A2(n_591),
.B1(n_599),
.B2(n_589),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_606),
.B(n_591),
.Y(n_616)
);

INVx5_ASAP7_75t_L g617 ( 
.A(n_609),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_610),
.A2(n_566),
.B1(n_592),
.B2(n_575),
.Y(n_618)
);

AOI21xp33_ASAP7_75t_SL g619 ( 
.A1(n_616),
.A2(n_597),
.B(n_604),
.Y(n_619)
);

NAND3xp33_ASAP7_75t_L g620 ( 
.A(n_615),
.B(n_584),
.C(n_594),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_612),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_618),
.A2(n_613),
.B(n_614),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_L g623 ( 
.A1(n_617),
.A2(n_584),
.B(n_611),
.Y(n_623)
);

NAND3xp33_ASAP7_75t_SL g624 ( 
.A(n_622),
.B(n_588),
.C(n_586),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_621),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_620),
.A2(n_619),
.B1(n_617),
.B2(n_623),
.Y(n_626)
);

O2A1O1Ixp5_ASAP7_75t_SL g627 ( 
.A1(n_621),
.A2(n_602),
.B(n_577),
.C(n_617),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_621),
.Y(n_628)
);

NAND3xp33_ASAP7_75t_L g629 ( 
.A(n_626),
.B(n_587),
.C(n_561),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_625),
.B(n_607),
.Y(n_630)
);

AOI221xp5_ASAP7_75t_L g631 ( 
.A1(n_624),
.A2(n_603),
.B1(n_595),
.B2(n_593),
.C(n_579),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_630),
.B(n_628),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_629),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_633),
.A2(n_632),
.B(n_631),
.Y(n_634)
);

NOR2xp67_ASAP7_75t_L g635 ( 
.A(n_634),
.B(n_632),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_635),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_636),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_637),
.A2(n_627),
.B1(n_579),
.B2(n_585),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_638),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_639),
.A2(n_585),
.B1(n_580),
.B2(n_567),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_640),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_641),
.B(n_113),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_SL g643 ( 
.A1(n_642),
.A2(n_567),
.B1(n_560),
.B2(n_580),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_SL g644 ( 
.A1(n_642),
.A2(n_560),
.B1(n_580),
.B2(n_541),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_643),
.B(n_644),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_SL g646 ( 
.A1(n_645),
.A2(n_560),
.B1(n_541),
.B2(n_116),
.Y(n_646)
);


endmodule