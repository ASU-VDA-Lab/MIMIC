module fake_jpeg_30132_n_99 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_10),
.B(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_46),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_49),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_50),
.B(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_52),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_42),
.C(n_41),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_53),
.A2(n_5),
.B(n_8),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_61),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_37),
.B1(n_32),
.B2(n_21),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_44),
.B1(n_3),
.B2(n_4),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_1),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_58),
.B(n_1),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_63),
.B(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_65),
.Y(n_78)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_68),
.Y(n_76)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_55),
.Y(n_69)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

AO22x1_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_11),
.B(n_14),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_2),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_74),
.Y(n_79)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_82),
.Y(n_89)
);

AOI211xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_85),
.B(n_22),
.C(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_15),
.Y(n_82)
);

OAI22x1_ASAP7_75t_SL g85 ( 
.A1(n_69),
.A2(n_16),
.B1(n_19),
.B2(n_20),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_83),
.B1(n_84),
.B2(n_76),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_75),
.C(n_23),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_88),
.A2(n_90),
.B1(n_85),
.B2(n_81),
.Y(n_91)
);

AO221x1_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_92),
.B1(n_75),
.B2(n_84),
.C(n_89),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_92),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_79),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_83),
.B(n_26),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_30),
.Y(n_99)
);


endmodule