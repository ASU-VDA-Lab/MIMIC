module fake_jpeg_12488_n_296 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_296);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_45),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_24),
.B(n_18),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_46),
.B(n_52),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_57),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_24),
.B(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_37),
.B1(n_41),
.B2(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_63),
.A2(n_37),
.B1(n_35),
.B2(n_30),
.Y(n_66)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_66),
.A2(n_77),
.B1(n_85),
.B2(n_97),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_19),
.C(n_26),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_62),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_70),
.A2(n_80),
.B1(n_82),
.B2(n_90),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_55),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_22),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_20),
.B1(n_35),
.B2(n_30),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_78),
.B(n_22),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_19),
.B1(n_26),
.B2(n_31),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_26),
.B1(n_38),
.B2(n_31),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_42),
.A2(n_20),
.B1(n_35),
.B2(n_30),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_57),
.B(n_41),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_60),
.A2(n_38),
.B1(n_31),
.B2(n_26),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_64),
.A2(n_20),
.B1(n_36),
.B2(n_39),
.Y(n_97)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_59),
.A2(n_40),
.B1(n_39),
.B2(n_38),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_47),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_119),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_104),
.B(n_107),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_75),
.B1(n_27),
.B2(n_28),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_80),
.B1(n_82),
.B2(n_66),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_28),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_27),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

INVx2_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_111),
.B(n_122),
.Y(n_165)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_113),
.A2(n_76),
.B1(n_99),
.B2(n_62),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_40),
.C(n_17),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_117),
.B(n_133),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_23),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_101),
.B(n_69),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_126),
.Y(n_146)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_67),
.B(n_38),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_136),
.Y(n_143)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_69),
.B(n_50),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_45),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_129),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_71),
.B(n_48),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_79),
.A2(n_48),
.B1(n_43),
.B2(n_50),
.Y(n_131)
);

OAI22x1_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_44),
.B1(n_53),
.B2(n_58),
.Y(n_151)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_45),
.Y(n_135)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_76),
.B(n_31),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_128),
.B1(n_73),
.B2(n_126),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_91),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_125),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_128),
.B(n_87),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_91),
.B(n_84),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_154),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_100),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_113),
.A2(n_87),
.B1(n_73),
.B2(n_96),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_129),
.B1(n_118),
.B2(n_110),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_112),
.B(n_103),
.C(n_136),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_4),
.Y(n_190)
);

AND2x6_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_3),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_3),
.Y(n_172)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_174),
.B1(n_182),
.B2(n_194),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_169),
.A2(n_180),
.B1(n_186),
.B2(n_195),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_138),
.B(n_111),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_170),
.B(n_178),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_175),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_189),
.Y(n_215)
);

AOI22x1_ASAP7_75t_SL g177 ( 
.A1(n_146),
.A2(n_134),
.B1(n_114),
.B2(n_109),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_165),
.B(n_151),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_130),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_158),
.B(n_4),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_179),
.B(n_183),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_139),
.A2(n_143),
.B1(n_154),
.B2(n_165),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_162),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_184),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_105),
.B1(n_132),
.B2(n_120),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_159),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_123),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_115),
.B1(n_89),
.B2(n_96),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_115),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_147),
.B(n_99),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_190),
.A2(n_153),
.B(n_137),
.Y(n_203)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

FAx1_ASAP7_75t_SL g193 ( 
.A(n_160),
.B(n_4),
.CI(n_5),
.CON(n_193),
.SN(n_193)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_193),
.B(n_5),
.CI(n_6),
.CON(n_206),
.SN(n_206)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_152),
.A2(n_89),
.B1(n_116),
.B2(n_133),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_156),
.A2(n_116),
.B1(n_133),
.B2(n_25),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_161),
.A3(n_150),
.B1(n_137),
.B2(n_148),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_212),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_203),
.B(n_186),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_180),
.A2(n_148),
.B1(n_163),
.B2(n_157),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_216),
.B1(n_218),
.B2(n_182),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_193),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_153),
.B(n_157),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_207),
.A2(n_211),
.B(n_214),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_173),
.A2(n_163),
.B(n_6),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_190),
.A2(n_5),
.A3(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_11),
.B(n_12),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_169),
.A2(n_25),
.B1(n_13),
.B2(n_14),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_167),
.A2(n_25),
.B1(n_14),
.B2(n_15),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_213),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_220),
.A2(n_225),
.B1(n_228),
.B2(n_224),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_210),
.B(n_183),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_221),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_176),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_226),
.C(n_227),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_236),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_189),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_184),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_174),
.C(n_168),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_231),
.C(n_211),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_196),
.A2(n_194),
.B1(n_195),
.B2(n_167),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_177),
.Y(n_231)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_170),
.B1(n_167),
.B2(n_193),
.Y(n_233)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_234),
.B(n_235),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_219),
.B(n_179),
.Y(n_235)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_240),
.A2(n_243),
.B1(n_245),
.B2(n_248),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_196),
.B1(n_218),
.B2(n_204),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_216),
.B1(n_203),
.B2(n_209),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_246),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_201),
.B1(n_208),
.B2(n_168),
.Y(n_248)
);

OAI321xp33_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_202),
.A3(n_206),
.B1(n_212),
.B2(n_192),
.C(n_214),
.Y(n_250)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_232),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_223),
.C(n_226),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_258),
.C(n_261),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_252),
.B(n_227),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_257),
.B(n_263),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_231),
.C(n_230),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_238),
.B(n_234),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_259),
.A2(n_243),
.B(n_236),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_238),
.C(n_222),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_175),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_187),
.C(n_191),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_239),
.C(n_248),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_268),
.B(n_269),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_262),
.A2(n_241),
.B1(n_251),
.B2(n_249),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_249),
.C(n_245),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_274),
.C(n_265),
.Y(n_277)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_273),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_258),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_277),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_261),
.C(n_260),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_278),
.B(n_12),
.Y(n_284)
);

BUFx4f_ASAP7_75t_SL g279 ( 
.A(n_267),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_254),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_274),
.B(n_206),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_270),
.C(n_268),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_285),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_286),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_279),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_15),
.B(n_16),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_280),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_279),
.B(n_281),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_287),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_292),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_15),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_16),
.B1(n_25),
.B2(n_260),
.Y(n_296)
);


endmodule