module fake_jpeg_7778_n_105 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_105);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_49),
.B(n_54),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_35),
.B1(n_48),
.B2(n_47),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_60),
.A2(n_63),
.B1(n_65),
.B2(n_22),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_2),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_14),
.B(n_16),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_37),
.B1(n_35),
.B2(n_38),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_45),
.B1(n_41),
.B2(n_40),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_71),
.B1(n_75),
.B2(n_77),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_72),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_76),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_13),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_74),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_66),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_70),
.B1(n_69),
.B2(n_63),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_81),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_91),
.B1(n_90),
.B2(n_83),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_82),
.B1(n_92),
.B2(n_87),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_95),
.A2(n_64),
.B(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_88),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_100),
.B(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_23),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_24),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_25),
.B(n_29),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_30),
.Y(n_105)
);


endmodule