module fake_jpeg_16662_n_305 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_305);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_40),
.Y(n_102)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_44),
.Y(n_66)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_54),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_8),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_59),
.Y(n_71)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_8),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_62),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_15),
.B(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_65),
.Y(n_89)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_22),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_73),
.B(n_83),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_35),
.B1(n_37),
.B2(n_18),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_74),
.A2(n_108),
.B1(n_24),
.B2(n_33),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_37),
.B1(n_18),
.B2(n_36),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_76),
.A2(n_103),
.B1(n_30),
.B2(n_23),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_81),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_58),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_42),
.B(n_15),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_25),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_92),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_22),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_29),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_93),
.A2(n_95),
.B1(n_20),
.B2(n_1),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_64),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_20),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_29),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_26),
.Y(n_96)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_43),
.B(n_26),
.Y(n_97)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_40),
.B(n_27),
.Y(n_98)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_41),
.B(n_27),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_100),
.B(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_39),
.B(n_36),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_53),
.A2(n_18),
.B1(n_29),
.B2(n_28),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_44),
.B(n_34),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_24),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_55),
.B(n_25),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_38),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_46),
.A2(n_30),
.B1(n_34),
.B2(n_28),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_88),
.B(n_91),
.C(n_71),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_114),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_76),
.A2(n_63),
.B1(n_61),
.B2(n_38),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_107),
.B1(n_79),
.B2(n_72),
.Y(n_152)
);

OAI22x1_ASAP7_75t_L g166 ( 
.A1(n_112),
.A2(n_115),
.B1(n_145),
.B2(n_150),
.Y(n_166)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_87),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_113),
.A2(n_70),
.B1(n_87),
.B2(n_0),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_23),
.Y(n_114)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_93),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_87),
.C(n_102),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_129),
.Y(n_156)
);

NAND2xp33_ASAP7_75t_SL g120 ( 
.A(n_85),
.B(n_24),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_120),
.A2(n_121),
.B(n_128),
.Y(n_163)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_85),
.B(n_24),
.Y(n_121)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_33),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_99),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_137),
.Y(n_165)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_38),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_133),
.B(n_142),
.Y(n_175)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_80),
.B1(n_79),
.B2(n_107),
.Y(n_135)
);

AO22x1_ASAP7_75t_SL g164 ( 
.A1(n_135),
.A2(n_102),
.B1(n_78),
.B2(n_67),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_66),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_89),
.A2(n_38),
.A3(n_33),
.B1(n_32),
.B2(n_20),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_146),
.B1(n_102),
.B2(n_84),
.Y(n_167)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_140),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_93),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_33),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_84),
.B(n_20),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_144),
.B(n_147),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_95),
.B(n_9),
.Y(n_147)
);

BUFx4f_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_106),
.A2(n_11),
.B1(n_13),
.B2(n_5),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_152),
.A2(n_168),
.B1(n_172),
.B2(n_174),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_157),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_83),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_72),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_158),
.B(n_161),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_186),
.C(n_125),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_69),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_167),
.B1(n_148),
.B2(n_135),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_69),
.B1(n_70),
.B2(n_5),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_117),
.B(n_87),
.Y(n_169)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_113),
.B1(n_141),
.B2(n_134),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_112),
.A2(n_0),
.B1(n_2),
.B2(n_6),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_145),
.A2(n_0),
.B1(n_2),
.B2(n_6),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_127),
.B(n_12),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_178),
.B(n_181),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_0),
.Y(n_180)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_13),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_120),
.A2(n_121),
.B1(n_135),
.B2(n_116),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_182),
.A2(n_168),
.B1(n_158),
.B2(n_152),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_14),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_136),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_110),
.B(n_14),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_189),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_119),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_SL g232 ( 
.A1(n_191),
.A2(n_195),
.B(n_205),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_171),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_194),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_179),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_166),
.A2(n_135),
.B1(n_131),
.B2(n_149),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_196),
.A2(n_202),
.B1(n_210),
.B2(n_216),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_148),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_201),
.C(n_190),
.Y(n_235)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_166),
.A2(n_139),
.B1(n_146),
.B2(n_118),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_182),
.A2(n_2),
.B(n_163),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_203),
.A2(n_215),
.B(n_211),
.Y(n_241)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_179),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_206),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_156),
.B(n_155),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_153),
.Y(n_207)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_177),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_213),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_159),
.A2(n_161),
.B1(n_167),
.B2(n_151),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_217),
.B1(n_192),
.B2(n_187),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_173),
.Y(n_214)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_176),
.A2(n_164),
.B(n_157),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_162),
.A2(n_151),
.B1(n_164),
.B2(n_172),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_173),
.A2(n_180),
.B1(n_174),
.B2(n_183),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_215),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_222),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_186),
.Y(n_219)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_203),
.A2(n_177),
.B(n_154),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_220),
.A2(n_241),
.B(n_199),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_200),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_154),
.B(n_207),
.Y(n_224)
);

NAND3xp33_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_233),
.C(n_227),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_226),
.A2(n_232),
.B1(n_218),
.B2(n_238),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_236),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_202),
.A2(n_210),
.B(n_195),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_231),
.A2(n_212),
.B(n_217),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_211),
.Y(n_234)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_242),
.C(n_219),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_193),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_216),
.B(n_192),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_223),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_204),
.Y(n_240)
);

AO221x1_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_214),
.B1(n_209),
.B2(n_199),
.C(n_201),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_198),
.B(n_190),
.Y(n_242)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_243),
.A2(n_245),
.B(n_249),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_252),
.C(n_248),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_247),
.A2(n_245),
.B1(n_258),
.B2(n_260),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_233),
.B(n_228),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_257),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_234),
.C(n_237),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_246),
.C(n_248),
.Y(n_264)
);

AOI322xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_241),
.A3(n_231),
.B1(n_226),
.B2(n_220),
.C1(n_228),
.C2(n_229),
.Y(n_253)
);

OA21x2_ASAP7_75t_SL g270 ( 
.A1(n_253),
.A2(n_260),
.B(n_244),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_220),
.A2(n_229),
.B(n_227),
.C(n_236),
.Y(n_257)
);

AND2x4_ASAP7_75t_SL g258 ( 
.A(n_222),
.B(n_240),
.Y(n_258)
);

AO21x1_ASAP7_75t_L g266 ( 
.A1(n_258),
.A2(n_254),
.B(n_251),
.Y(n_266)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_221),
.Y(n_259)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

OA21x2_ASAP7_75t_SL g260 ( 
.A1(n_225),
.A2(n_239),
.B(n_221),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_258),
.Y(n_269)
);

OAI321xp33_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_223),
.A3(n_225),
.B1(n_239),
.B2(n_261),
.C(n_254),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_262),
.A2(n_270),
.B1(n_273),
.B2(n_255),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_271),
.C(n_256),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_274),
.Y(n_280)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_259),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_272),
.B(n_255),
.Y(n_285)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_276),
.C(n_279),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_247),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_257),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_281),
.B(n_262),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_256),
.C(n_250),
.Y(n_279)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_263),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_283),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_270),
.C(n_263),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_266),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_278),
.A2(n_272),
.B1(n_267),
.B2(n_265),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_287),
.A2(n_269),
.B1(n_284),
.B2(n_292),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_293),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_273),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_290),
.C(n_277),
.Y(n_295)
);

AOI21xp33_ASAP7_75t_SL g290 ( 
.A1(n_276),
.A2(n_266),
.B(n_268),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_295),
.A2(n_286),
.B1(n_287),
.B2(n_294),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_267),
.Y(n_296)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_296),
.Y(n_301)
);

NAND2x1_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_284),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_298),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_301),
.A2(n_296),
.B(n_297),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_303),
.B(n_300),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_302),
.Y(n_305)
);


endmodule