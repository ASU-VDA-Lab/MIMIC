module fake_netlist_5_617_n_1968 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1968);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1968;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_696;
wire n_550;
wire n_897;
wire n_215;
wire n_798;
wire n_196;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_1163;
wire n_906;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_192;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1944;
wire n_909;
wire n_1817;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g189 ( 
.A(n_65),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_89),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_39),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_18),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_35),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_167),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_144),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_59),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_140),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_42),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_175),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_128),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_72),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_80),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_26),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_44),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_164),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_24),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_0),
.Y(n_210)
);

BUFx2_ASAP7_75t_SL g211 ( 
.A(n_156),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_102),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_143),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_78),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_11),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_174),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_3),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_176),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_107),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_75),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_170),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_124),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_31),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_57),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_147),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_37),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_16),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_40),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_20),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_70),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_169),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_136),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_112),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_94),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_9),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_52),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_74),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_68),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_64),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_114),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_4),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_118),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_184),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_51),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_104),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_125),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_39),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_15),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_105),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_101),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_91),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_186),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_163),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_178),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_11),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_151),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_88),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_76),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_171),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_132),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_15),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_30),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_109),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_90),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_162),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_23),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_134),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_10),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_79),
.Y(n_270)
);

BUFx8_ASAP7_75t_SL g271 ( 
.A(n_4),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_8),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_7),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_152),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_160),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_36),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_64),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_21),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_99),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_123),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_57),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_87),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_34),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_31),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_172),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_86),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_155),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_8),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_20),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_95),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_121),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_137),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_3),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_179),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_111),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_146),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_84),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_29),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_182),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_117),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_93),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_6),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_51),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_13),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_29),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_52),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_7),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_53),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_63),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_122),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_138),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_28),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_38),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_139),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_166),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_131),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_185),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_98),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_65),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_10),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_133),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_36),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_71),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_23),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_17),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_21),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_100),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_54),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_58),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_41),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_27),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_62),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_41),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_53),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_18),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_24),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_165),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_14),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_44),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_129),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_153),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_187),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_119),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_61),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_25),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_127),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_82),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_43),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_183),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_14),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_54),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_159),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_142),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_45),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_60),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_110),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_63),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_5),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_32),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_6),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_92),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_34),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_47),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_13),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_12),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_145),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_62),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_154),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_5),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_130),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_55),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_26),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_116),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_32),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_81),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_362),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_271),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_340),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_270),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_190),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_362),
.Y(n_381)
);

BUFx2_ASAP7_75t_SL g382 ( 
.A(n_291),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_362),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_362),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_198),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_328),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_192),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_197),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_362),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_200),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_287),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_213),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_263),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_202),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_302),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_255),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_263),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_263),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_204),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_191),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_322),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_322),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_205),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_322),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_363),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_363),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_213),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_196),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_363),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_208),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_307),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_307),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_308),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_308),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_267),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_213),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_267),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_267),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_191),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_288),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_288),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_212),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_288),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_330),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_330),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_260),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_330),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_214),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_338),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_216),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_338),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_338),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_189),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_189),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_220),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_219),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_221),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_201),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_201),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_218),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_222),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_260),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_207),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_199),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_234),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_361),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_206),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_238),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_207),
.Y(n_452)
);

CKINVDCx14_ASAP7_75t_R g453 ( 
.A(n_361),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_239),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_209),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_241),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_222),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_243),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_210),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_246),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_247),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_302),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_210),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_224),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_219),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_224),
.Y(n_466)
);

INVxp33_ASAP7_75t_SL g467 ( 
.A(n_215),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_251),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_225),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_225),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_222),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_380),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_398),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_376),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_398),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_386),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_404),
.B(n_219),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_438),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_376),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_381),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_398),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_398),
.Y(n_483)
);

NOR2x1_ASAP7_75t_L g484 ( 
.A(n_394),
.B(n_317),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_381),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_388),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_383),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_398),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_394),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_394),
.A2(n_317),
.B(n_266),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_438),
.B(n_291),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_404),
.B(n_317),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_409),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_409),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_409),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_L g496 ( 
.A(n_417),
.B(n_336),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_418),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_383),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_438),
.B(n_301),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_384),
.B(n_317),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_453),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_389),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_396),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_384),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_401),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_410),
.A2(n_195),
.B1(n_312),
.B2(n_217),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_418),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_418),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_390),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_410),
.A2(n_371),
.B1(n_303),
.B2(n_236),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_443),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_443),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_443),
.Y(n_513)
);

OA21x2_ASAP7_75t_L g514 ( 
.A1(n_457),
.A2(n_229),
.B(n_227),
.Y(n_514)
);

OA21x2_ASAP7_75t_L g515 ( 
.A1(n_457),
.A2(n_229),
.B(n_227),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_390),
.B(n_301),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_457),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_465),
.B(n_253),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_391),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_465),
.B(n_254),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_471),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_379),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_471),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_471),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_391),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_435),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_395),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_385),
.A2(n_193),
.B1(n_336),
.B2(n_354),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_393),
.B(n_302),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_465),
.B(n_257),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_447),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_408),
.B(n_261),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_435),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_395),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_436),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_436),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_399),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_440),
.Y(n_538)
);

OA21x2_ASAP7_75t_L g539 ( 
.A1(n_399),
.A2(n_256),
.B(n_230),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_382),
.B(n_346),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_400),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_440),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_400),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_441),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_397),
.A2(n_462),
.B1(n_392),
.B2(n_442),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_403),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_441),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_403),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_455),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_406),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_446),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_506),
.A2(n_402),
.B1(n_428),
.B2(n_421),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_L g553 ( 
.A(n_492),
.B(n_449),
.C(n_444),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_493),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_479),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_479),
.B(n_405),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_493),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g558 ( 
.A(n_479),
.B(n_412),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_501),
.B(n_393),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_518),
.B(n_424),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_514),
.Y(n_561)
);

INVxp33_ASAP7_75t_SL g562 ( 
.A(n_545),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_478),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_525),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_492),
.B(n_408),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_525),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_518),
.B(n_430),
.Y(n_567)
);

NOR2x1p5_ASAP7_75t_L g568 ( 
.A(n_472),
.B(n_377),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_514),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_525),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_520),
.B(n_437),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_525),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_514),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_SL g574 ( 
.A1(n_506),
.A2(n_462),
.B1(n_397),
.B2(n_432),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_514),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_501),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_514),
.Y(n_577)
);

AND3x1_ASAP7_75t_L g578 ( 
.A(n_510),
.B(n_387),
.C(n_445),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_514),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_493),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_515),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_515),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_501),
.B(n_439),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_515),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_515),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_482),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_528),
.A2(n_510),
.B1(n_378),
.B2(n_549),
.Y(n_587)
);

AO22x2_ASAP7_75t_L g588 ( 
.A1(n_528),
.A2(n_266),
.B1(n_279),
.B2(n_264),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_493),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_532),
.B(n_467),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_520),
.B(n_451),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_486),
.B(n_454),
.Y(n_592)
);

INVxp67_ASAP7_75t_SL g593 ( 
.A(n_475),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_515),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_549),
.A2(n_228),
.B1(n_240),
.B2(n_237),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_482),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_515),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_539),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_494),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_R g600 ( 
.A(n_549),
.B(n_455),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_532),
.B(n_456),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_530),
.B(n_492),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_494),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_494),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_539),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_502),
.B(n_460),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_478),
.A2(n_382),
.B1(n_230),
.B2(n_273),
.Y(n_607)
);

AO22x2_ASAP7_75t_L g608 ( 
.A1(n_529),
.A2(n_264),
.B1(n_279),
.B2(n_266),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_539),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_494),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_482),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_539),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_539),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_539),
.Y(n_614)
);

BUFx10_ASAP7_75t_L g615 ( 
.A(n_503),
.Y(n_615)
);

CKINVDCx11_ASAP7_75t_R g616 ( 
.A(n_477),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_505),
.B(n_461),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_482),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_497),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_482),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_540),
.B(n_448),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_530),
.B(n_450),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_497),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_497),
.Y(n_624)
);

NAND3xp33_ASAP7_75t_L g625 ( 
.A(n_491),
.B(n_419),
.C(n_417),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_529),
.A2(n_245),
.B1(n_248),
.B2(n_242),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_540),
.B(n_231),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_531),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_478),
.A2(n_256),
.B1(n_283),
.B2(n_273),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_474),
.Y(n_630)
);

AND3x2_ASAP7_75t_L g631 ( 
.A(n_522),
.B(n_279),
.C(n_264),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_497),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_474),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_507),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_531),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_522),
.B(n_458),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_480),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_482),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_482),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_522),
.B(n_468),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_480),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_507),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_491),
.B(n_265),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_499),
.B(n_232),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_516),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_499),
.B(n_419),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_526),
.B(n_420),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_516),
.B(n_274),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_507),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_481),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_507),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_511),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_477),
.Y(n_653)
);

INVx5_ASAP7_75t_L g654 ( 
.A(n_482),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_481),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_495),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_511),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_545),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_511),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_513),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_516),
.B(n_280),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_513),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_495),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_495),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_485),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_495),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_516),
.B(n_285),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_485),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_513),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_490),
.Y(n_670)
);

NOR2x1p5_ASAP7_75t_L g671 ( 
.A(n_526),
.B(n_283),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_533),
.B(n_420),
.Y(n_672)
);

AND3x1_ASAP7_75t_L g673 ( 
.A(n_533),
.B(n_293),
.C(n_289),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_535),
.B(n_286),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_535),
.B(n_290),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_487),
.Y(n_676)
);

BUFx10_ASAP7_75t_L g677 ( 
.A(n_500),
.Y(n_677)
);

INVxp33_ASAP7_75t_L g678 ( 
.A(n_551),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_513),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_517),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_517),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_536),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_500),
.A2(n_364),
.B1(n_289),
.B2(n_293),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_496),
.A2(n_319),
.B1(n_324),
.B2(n_325),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_536),
.B(n_294),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_500),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_500),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_500),
.A2(n_364),
.B1(n_313),
.B2(n_348),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_517),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_487),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_538),
.B(n_422),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_517),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_498),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_523),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_538),
.B(n_295),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_542),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_498),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_475),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_542),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_L g700 ( 
.A(n_484),
.B(n_255),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_495),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_523),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_635),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_584),
.Y(n_704)
);

NOR2xp67_ASAP7_75t_L g705 ( 
.A(n_590),
.B(n_544),
.Y(n_705)
);

BUFx6f_ASAP7_75t_SL g706 ( 
.A(n_615),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_687),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_563),
.B(n_370),
.Y(n_708)
);

O2A1O1Ixp5_ASAP7_75t_L g709 ( 
.A1(n_598),
.A2(n_315),
.B(n_318),
.C(n_314),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_565),
.B(n_504),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_687),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_563),
.B(n_299),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_635),
.B(n_422),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_565),
.B(n_300),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_565),
.B(n_504),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_600),
.Y(n_716)
);

NOR2x1p5_ASAP7_75t_L g717 ( 
.A(n_622),
.B(n_249),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_565),
.B(n_509),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_601),
.B(n_509),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_687),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_584),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_628),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_628),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_602),
.A2(n_310),
.B1(n_316),
.B2(n_311),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_627),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_677),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_678),
.B(n_682),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_699),
.B(n_423),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_555),
.B(n_645),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_576),
.Y(n_730)
);

HB1xp67_ASAP7_75t_L g731 ( 
.A(n_653),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_555),
.B(n_519),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_686),
.B(n_255),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_553),
.B(n_262),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_696),
.B(n_537),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_696),
.B(n_537),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_677),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_686),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_584),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_691),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_553),
.B(n_269),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_646),
.B(n_537),
.Y(n_742)
);

INVxp33_ASAP7_75t_L g743 ( 
.A(n_616),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_644),
.B(n_537),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_699),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_691),
.B(n_423),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_560),
.B(n_272),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_567),
.B(n_276),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_677),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_630),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_598),
.A2(n_490),
.B(n_315),
.C(n_318),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_571),
.B(n_591),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_561),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_630),
.Y(n_754)
);

NOR2x1p5_ASAP7_75t_L g755 ( 
.A(n_556),
.B(n_277),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_561),
.B(n_537),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_633),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_621),
.B(n_278),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_615),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_569),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_569),
.B(n_475),
.Y(n_761)
);

AND2x6_ASAP7_75t_L g762 ( 
.A(n_573),
.B(n_575),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_615),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_L g764 ( 
.A(n_670),
.B(n_342),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_573),
.B(n_475),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_626),
.B(n_281),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_575),
.B(n_475),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_577),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_607),
.B(n_352),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_577),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_605),
.B(n_255),
.Y(n_771)
);

NOR3xp33_ASAP7_75t_L g772 ( 
.A(n_574),
.B(n_496),
.C(n_426),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_626),
.B(n_353),
.Y(n_773)
);

BUFx5_ASAP7_75t_L g774 ( 
.A(n_579),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_579),
.B(n_476),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_581),
.B(n_476),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_581),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_677),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_643),
.B(n_284),
.Y(n_779)
);

BUFx6f_ASAP7_75t_SL g780 ( 
.A(n_615),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_605),
.A2(n_331),
.B1(n_355),
.B2(n_354),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_582),
.B(n_476),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_671),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_593),
.A2(n_484),
.B(n_483),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_582),
.B(n_585),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_595),
.B(n_356),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_585),
.B(n_476),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_698),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_671),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_595),
.B(n_298),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_594),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_587),
.B(n_366),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_587),
.B(n_425),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_592),
.B(n_304),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_684),
.B(n_368),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_684),
.B(n_373),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_594),
.B(n_476),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_631),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_629),
.B(n_552),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_606),
.B(n_305),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_617),
.B(n_375),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_597),
.B(n_488),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_558),
.A2(n_211),
.B1(n_321),
.B2(n_297),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_637),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_597),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_609),
.B(n_255),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_583),
.B(n_306),
.Y(n_807)
);

NOR2xp67_ASAP7_75t_L g808 ( 
.A(n_625),
.B(n_544),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_673),
.B(n_648),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_559),
.B(n_425),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_608),
.A2(n_612),
.B1(n_614),
.B2(n_613),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_673),
.B(n_255),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_612),
.B(n_314),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_613),
.B(n_314),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_637),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_608),
.A2(n_211),
.B1(n_347),
.B2(n_343),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_641),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_698),
.Y(n_818)
);

INVx8_ASAP7_75t_L g819 ( 
.A(n_670),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_641),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_578),
.B(n_426),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_650),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_674),
.B(n_309),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_614),
.B(n_488),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_650),
.Y(n_825)
);

NOR2xp67_ASAP7_75t_L g826 ( 
.A(n_625),
.B(n_547),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_670),
.B(n_315),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_655),
.B(n_488),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_698),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_665),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_665),
.B(n_488),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_668),
.B(n_488),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_568),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_608),
.A2(n_318),
.B1(n_327),
.B2(n_337),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_608),
.A2(n_327),
.B1(n_337),
.B2(n_259),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_578),
.B(n_427),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_661),
.B(n_667),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_670),
.Y(n_838)
);

NAND2xp33_ASAP7_75t_L g839 ( 
.A(n_670),
.B(n_327),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_596),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_668),
.B(n_194),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_647),
.B(n_427),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_675),
.B(n_320),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_676),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_676),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_690),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_690),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_693),
.B(n_547),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_588),
.A2(n_313),
.B1(n_355),
.B2(n_326),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_685),
.A2(n_282),
.B1(n_349),
.B2(n_347),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_695),
.B(n_329),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_697),
.B(n_194),
.Y(n_852)
);

AND2x4_ASAP7_75t_SL g853 ( 
.A(n_683),
.B(n_302),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_588),
.A2(n_275),
.B1(n_349),
.B2(n_343),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_697),
.B(n_203),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_596),
.B(n_203),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_564),
.Y(n_857)
);

NAND2xp33_ASAP7_75t_L g858 ( 
.A(n_688),
.B(n_223),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_596),
.B(n_226),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_596),
.B(n_233),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_588),
.Y(n_861)
);

NAND2xp33_ASAP7_75t_L g862 ( 
.A(n_611),
.B(n_618),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_611),
.B(n_235),
.Y(n_863)
);

BUFx8_ASAP7_75t_SL g864 ( 
.A(n_562),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_611),
.B(n_235),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_672),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_618),
.B(n_244),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_752),
.A2(n_719),
.B1(n_725),
.B2(n_721),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_838),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_708),
.B(n_618),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_825),
.Y(n_871)
);

AND2x6_ASAP7_75t_SL g872 ( 
.A(n_790),
.B(n_326),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_722),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_708),
.B(n_618),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_866),
.B(n_620),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_825),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_845),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_705),
.B(n_620),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_783),
.B(n_568),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_747),
.B(n_620),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_716),
.B(n_658),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_838),
.B(n_620),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_846),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_747),
.B(n_638),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_727),
.B(n_636),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_748),
.B(n_638),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_748),
.A2(n_640),
.B1(n_588),
.B2(n_700),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_707),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_774),
.B(n_638),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_846),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_848),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_774),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_848),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_745),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_857),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_728),
.Y(n_896)
);

AND2x6_ASAP7_75t_L g897 ( 
.A(n_838),
.B(n_704),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_766),
.A2(n_639),
.B1(n_638),
.B2(n_701),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_857),
.Y(n_899)
);

OR2x6_ASAP7_75t_L g900 ( 
.A(n_723),
.B(n_244),
.Y(n_900)
);

OR2x6_ASAP7_75t_L g901 ( 
.A(n_730),
.B(n_250),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_738),
.Y(n_902)
);

BUFx4f_ASAP7_75t_L g903 ( 
.A(n_793),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_766),
.A2(n_639),
.B1(n_701),
.B2(n_656),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_774),
.B(n_639),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_711),
.A2(n_639),
.B1(n_701),
.B2(n_656),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_703),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_774),
.B(n_656),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_774),
.Y(n_909)
);

NOR2xp67_ASAP7_75t_L g910 ( 
.A(n_759),
.B(n_429),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_720),
.A2(n_666),
.B1(n_701),
.B2(n_656),
.Y(n_911)
);

INVxp67_ASAP7_75t_SL g912 ( 
.A(n_838),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_713),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_750),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_861),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_731),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_827),
.A2(n_490),
.B(n_564),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_819),
.A2(n_785),
.B(n_729),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_706),
.Y(n_919)
);

NOR2x1p5_ASAP7_75t_L g920 ( 
.A(n_833),
.B(n_429),
.Y(n_920)
);

INVx5_ASAP7_75t_L g921 ( 
.A(n_762),
.Y(n_921)
);

INVxp33_ASAP7_75t_L g922 ( 
.A(n_734),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_704),
.B(n_663),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_707),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_810),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_717),
.Y(n_926)
);

INVx8_ASAP7_75t_L g927 ( 
.A(n_762),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_754),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_842),
.B(n_753),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_753),
.B(n_663),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_760),
.B(n_663),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_819),
.A2(n_664),
.B(n_654),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_757),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_746),
.B(n_740),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_760),
.B(n_666),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_721),
.B(n_666),
.Y(n_936)
);

INVx5_ASAP7_75t_L g937 ( 
.A(n_762),
.Y(n_937)
);

INVxp67_ASAP7_75t_SL g938 ( 
.A(n_768),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_739),
.B(n_666),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_734),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_707),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_768),
.B(n_770),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_706),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_781),
.A2(n_348),
.B1(n_331),
.B2(n_250),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_770),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_707),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_819),
.A2(n_839),
.B(n_862),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_804),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_726),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_777),
.B(n_566),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_791),
.B(n_566),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_788),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_815),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_SL g954 ( 
.A1(n_790),
.A2(n_357),
.B1(n_332),
.B2(n_333),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_780),
.Y(n_955)
);

INVx5_ASAP7_75t_L g956 ( 
.A(n_762),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_817),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_788),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_789),
.B(n_431),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_791),
.B(n_570),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_820),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_798),
.B(n_818),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_822),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_726),
.B(n_664),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_805),
.B(n_570),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_809),
.A2(n_268),
.B1(n_259),
.B2(n_258),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_726),
.B(n_664),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_818),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_829),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_781),
.A2(n_252),
.B1(n_341),
.B2(n_323),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_755),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_805),
.B(n_572),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_726),
.B(n_664),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_830),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_844),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_778),
.B(n_572),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_L g977 ( 
.A(n_741),
.B(n_335),
.C(n_334),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_847),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_808),
.B(n_589),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_828),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_840),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_826),
.B(n_589),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_778),
.B(n_554),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_758),
.A2(n_252),
.B1(n_258),
.B2(n_268),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_762),
.Y(n_985)
);

INVx4_ASAP7_75t_L g986 ( 
.A(n_778),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_758),
.A2(n_275),
.B1(n_282),
.B2(n_292),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_761),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_772),
.B(n_431),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_840),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_799),
.A2(n_292),
.B1(n_341),
.B2(n_296),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_778),
.B(n_554),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_831),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_765),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_L g995 ( 
.A1(n_849),
.A2(n_741),
.B1(n_834),
.B2(n_835),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_744),
.B(n_599),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_821),
.B(n_433),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_836),
.B(n_433),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_832),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_742),
.B(n_599),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_710),
.B(n_603),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_715),
.B(n_554),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_837),
.A2(n_296),
.B1(n_297),
.B2(n_321),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_718),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_864),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_732),
.B(n_603),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_767),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_737),
.B(n_749),
.Y(n_1008)
);

BUFx4f_ASAP7_75t_L g1009 ( 
.A(n_853),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_792),
.B(n_339),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_775),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_849),
.A2(n_323),
.B1(n_551),
.B2(n_434),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_773),
.B(n_344),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_853),
.A2(n_434),
.B(n_470),
.C(n_469),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_786),
.B(n_807),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_776),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_735),
.Y(n_1017)
);

CKINVDCx6p67_ASAP7_75t_R g1018 ( 
.A(n_763),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_840),
.Y(n_1019)
);

NAND2xp33_ASAP7_75t_SL g1020 ( 
.A(n_811),
.B(n_345),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_737),
.B(n_623),
.Y(n_1021)
);

AOI21x1_ASAP7_75t_L g1022 ( 
.A1(n_771),
.A2(n_632),
.B(n_624),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_736),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_841),
.B(n_624),
.Y(n_1024)
);

OR2x4_ASAP7_75t_L g1025 ( 
.A(n_807),
.B(n_446),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_840),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_852),
.B(n_632),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_756),
.B(n_634),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_782),
.Y(n_1029)
);

INVx5_ASAP7_75t_L g1030 ( 
.A(n_709),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_787),
.Y(n_1031)
);

BUFx4f_ASAP7_75t_L g1032 ( 
.A(n_743),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_794),
.B(n_452),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_797),
.B(n_634),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_802),
.Y(n_1035)
);

INVx5_ASAP7_75t_L g1036 ( 
.A(n_764),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_856),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_800),
.B(n_350),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_800),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_824),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_714),
.B(n_642),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_712),
.B(n_459),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_865),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_855),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_779),
.B(n_642),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_816),
.B(n_557),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_949),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_916),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_1015),
.A2(n_823),
.B(n_843),
.C(n_851),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_922),
.B(n_1039),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_903),
.B(n_779),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_903),
.B(n_823),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_940),
.B(n_843),
.Y(n_1053)
);

BUFx4f_ASAP7_75t_L g1054 ( 
.A(n_1018),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_947),
.A2(n_827),
.B(n_806),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_940),
.B(n_851),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_885),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_894),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1038),
.A2(n_796),
.B1(n_795),
.B2(n_724),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_868),
.B(n_854),
.Y(n_1060)
);

NAND2x1p5_ASAP7_75t_L g1061 ( 
.A(n_986),
.B(n_859),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_938),
.A2(n_806),
.B(n_771),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_962),
.B(n_801),
.Y(n_1063)
);

NOR3xp33_ASAP7_75t_L g1064 ( 
.A(n_1038),
.B(n_769),
.C(n_858),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_880),
.A2(n_814),
.B(n_813),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_1005),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_884),
.A2(n_814),
.B(n_813),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_SL g1068 ( 
.A1(n_1015),
.A2(n_812),
.B(n_751),
.C(n_860),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_915),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_881),
.B(n_803),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_R g1071 ( 
.A(n_919),
.B(n_351),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_1010),
.A2(n_863),
.B(n_860),
.C(n_859),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_1010),
.A2(n_850),
.B(n_784),
.C(n_733),
.Y(n_1073)
);

NAND2xp33_ASAP7_75t_L g1074 ( 
.A(n_949),
.B(n_863),
.Y(n_1074)
);

BUFx5_ASAP7_75t_L g1075 ( 
.A(n_897),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_1014),
.A2(n_867),
.B(n_733),
.C(n_470),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_995),
.A2(n_867),
.B1(n_359),
.B2(n_360),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_SL g1078 ( 
.A1(n_1014),
.A2(n_557),
.B(n_580),
.C(n_604),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1004),
.B(n_651),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_873),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_915),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_894),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_995),
.A2(n_358),
.B1(n_365),
.B2(n_367),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_1013),
.A2(n_369),
.B(n_372),
.C(n_406),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_879),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_917),
.A2(n_649),
.B(n_557),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_934),
.B(n_651),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_997),
.B(n_652),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_871),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_886),
.A2(n_654),
.B(n_586),
.Y(n_1090)
);

AO32x1_ASAP7_75t_L g1091 ( 
.A1(n_876),
.A2(n_469),
.A3(n_466),
.B1(n_464),
.B2(n_463),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_881),
.B(n_0),
.Y(n_1092)
);

OR2x6_ASAP7_75t_L g1093 ( 
.A(n_927),
.B(n_913),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_896),
.B(n_1033),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_988),
.A2(n_649),
.B(n_580),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_896),
.B(n_1),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_925),
.B(n_1009),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_907),
.Y(n_1098)
);

OR2x6_ASAP7_75t_L g1099 ( 
.A(n_927),
.B(n_459),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_920),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_1009),
.B(n_652),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_949),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_877),
.Y(n_1103)
);

NOR2x1_ASAP7_75t_R g1104 ( 
.A(n_943),
.B(n_463),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_929),
.B(n_702),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_964),
.A2(n_654),
.B(n_586),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_970),
.A2(n_466),
.B1(n_464),
.B2(n_407),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_1025),
.B(n_1),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_890),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1025),
.B(n_2),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_970),
.A2(n_407),
.B1(n_411),
.B2(n_413),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_962),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_924),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_887),
.A2(n_411),
.B(n_413),
.C(n_414),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_945),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_879),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_964),
.A2(n_654),
.B(n_586),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_998),
.B(n_657),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_989),
.B(n_414),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_914),
.A2(n_415),
.B(n_416),
.C(n_692),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_959),
.B(n_541),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_944),
.A2(n_991),
.B1(n_1012),
.B2(n_942),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1029),
.B(n_657),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_944),
.A2(n_702),
.B1(n_694),
.B2(n_689),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_954),
.A2(n_694),
.B1(n_689),
.B2(n_681),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1031),
.B(n_659),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_928),
.A2(n_681),
.B(n_659),
.C(n_679),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_900),
.Y(n_1128)
);

NOR2x1_ASAP7_75t_SL g1129 ( 
.A(n_921),
.B(n_586),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_933),
.A2(n_660),
.B(n_679),
.C(n_669),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_967),
.A2(n_654),
.B(n_586),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_949),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_921),
.B(n_662),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_973),
.A2(n_654),
.B(n_586),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_954),
.A2(n_543),
.B1(n_548),
.B2(n_541),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1035),
.B(n_580),
.Y(n_1136)
);

NAND2x1p5_ASAP7_75t_L g1137 ( 
.A(n_986),
.B(n_604),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_901),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1017),
.B(n_604),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1023),
.B(n_610),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_924),
.Y(n_1141)
);

OAI21xp33_ASAP7_75t_L g1142 ( 
.A1(n_984),
.A2(n_680),
.B(n_649),
.Y(n_1142)
);

AOI21x1_ASAP7_75t_L g1143 ( 
.A1(n_976),
.A2(n_680),
.B(n_619),
.Y(n_1143)
);

CKINVDCx20_ASAP7_75t_R g1144 ( 
.A(n_1005),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_908),
.A2(n_524),
.B(n_523),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_889),
.A2(n_524),
.B(n_523),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_959),
.B(n_541),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1042),
.B(n_541),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_948),
.A2(n_680),
.B(n_619),
.C(n_610),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_921),
.B(n_610),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_891),
.B(n_2),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_900),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_900),
.Y(n_1153)
);

BUFx2_ASAP7_75t_SL g1154 ( 
.A(n_921),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_1032),
.Y(n_1155)
);

NAND3xp33_ASAP7_75t_SL g1156 ( 
.A(n_987),
.B(n_548),
.C(n_543),
.Y(n_1156)
);

NOR3xp33_ASAP7_75t_SL g1157 ( 
.A(n_955),
.B(n_9),
.C(n_12),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_924),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_893),
.B(n_17),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1042),
.B(n_543),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1040),
.B(n_619),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_1032),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_905),
.A2(n_524),
.B(n_495),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_883),
.Y(n_1164)
);

NAND3xp33_ASAP7_75t_L g1165 ( 
.A(n_977),
.B(n_550),
.C(n_527),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_952),
.A2(n_958),
.B1(n_910),
.B2(n_1044),
.Y(n_1166)
);

NOR3xp33_ASAP7_75t_SL g1167 ( 
.A(n_1020),
.B(n_19),
.C(n_22),
.Y(n_1167)
);

INVx6_ASAP7_75t_L g1168 ( 
.A(n_924),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_952),
.B(n_19),
.Y(n_1169)
);

NAND2xp33_ASAP7_75t_SL g1170 ( 
.A(n_971),
.B(n_550),
.Y(n_1170)
);

AOI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_958),
.A2(n_548),
.B1(n_543),
.B2(n_546),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_918),
.A2(n_524),
.B(n_495),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_901),
.B(n_548),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_901),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_902),
.B(n_22),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_953),
.B(n_27),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_R g1177 ( 
.A(n_1020),
.B(n_103),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_957),
.B(n_30),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_912),
.A2(n_512),
.B(n_495),
.Y(n_1179)
);

CKINVDCx8_ASAP7_75t_R g1180 ( 
.A(n_872),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_988),
.B(n_546),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_961),
.B(n_33),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_963),
.B(n_33),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_974),
.B(n_35),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_937),
.B(n_550),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_912),
.A2(n_512),
.B(n_508),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_975),
.A2(n_473),
.B(n_483),
.C(n_489),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_978),
.Y(n_1188)
);

NOR2x1_ASAP7_75t_SL g1189 ( 
.A(n_937),
.B(n_473),
.Y(n_1189)
);

AO32x1_ASAP7_75t_L g1190 ( 
.A1(n_1037),
.A2(n_473),
.A3(n_483),
.B1(n_40),
.B2(n_42),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1045),
.A2(n_512),
.B(n_508),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_941),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_892),
.A2(n_512),
.B(n_508),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_941),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_926),
.A2(n_473),
.B(n_483),
.C(n_489),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_994),
.B(n_546),
.Y(n_1196)
);

CKINVDCx6p67_ASAP7_75t_R g1197 ( 
.A(n_1155),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1143),
.A2(n_1022),
.B(n_976),
.Y(n_1198)
);

AOI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1055),
.A2(n_874),
.B(n_870),
.Y(n_1199)
);

AOI221x1_ASAP7_75t_L g1200 ( 
.A1(n_1049),
.A2(n_1000),
.B1(n_980),
.B2(n_993),
.C(n_999),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_SL g1201 ( 
.A1(n_1073),
.A2(n_1046),
.B(n_875),
.C(n_983),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_1114),
.A2(n_892),
.A3(n_909),
.B(n_1021),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1048),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1052),
.B(n_966),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1070),
.B(n_994),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1058),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1172),
.A2(n_983),
.B(n_992),
.Y(n_1207)
);

INVx4_ASAP7_75t_L g1208 ( 
.A(n_1113),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1057),
.B(n_1041),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1163),
.A2(n_1086),
.B(n_1191),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_1113),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1094),
.B(n_1007),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1188),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1059),
.A2(n_956),
.B1(n_937),
.B2(n_1036),
.Y(n_1214)
);

AOI21x1_ASAP7_75t_SL g1215 ( 
.A1(n_1060),
.A2(n_878),
.B(n_1008),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1086),
.A2(n_1002),
.B(n_935),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1065),
.A2(n_996),
.B(n_1046),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1193),
.A2(n_1002),
.B(n_931),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_SL g1219 ( 
.A1(n_1051),
.A2(n_882),
.B(n_979),
.C(n_982),
.Y(n_1219)
);

AO31x2_ASAP7_75t_L g1220 ( 
.A1(n_1067),
.A2(n_909),
.A3(n_1007),
.B(n_1011),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1089),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_1066),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1092),
.A2(n_991),
.B1(n_1003),
.B2(n_1043),
.Y(n_1223)
);

NAND2x1p5_ASAP7_75t_L g1224 ( 
.A(n_1113),
.B(n_937),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1145),
.A2(n_930),
.B(n_960),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1062),
.A2(n_1036),
.B(n_956),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1103),
.Y(n_1227)
);

OA21x2_ASAP7_75t_L g1228 ( 
.A1(n_1165),
.A2(n_1027),
.B(n_1024),
.Y(n_1228)
);

OR2x6_ASAP7_75t_L g1229 ( 
.A(n_1099),
.B(n_927),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1158),
.Y(n_1230)
);

AOI221xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1077),
.A2(n_1012),
.B1(n_1006),
.B2(n_1001),
.C(n_1011),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1053),
.B(n_1016),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1068),
.A2(n_1028),
.B(n_1034),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1109),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1072),
.A2(n_1036),
.B(n_956),
.Y(n_1235)
);

AO22x2_ASAP7_75t_L g1236 ( 
.A1(n_1083),
.A2(n_1077),
.B1(n_1056),
.B2(n_1122),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1085),
.B(n_1116),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1122),
.A2(n_1016),
.A3(n_972),
.B(n_951),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1121),
.B(n_968),
.Y(n_1239)
);

AOI221xp5_ASAP7_75t_L g1240 ( 
.A1(n_1083),
.A2(n_895),
.B1(n_899),
.B2(n_950),
.C(n_965),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1146),
.A2(n_904),
.B(n_898),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_SL g1242 ( 
.A1(n_1189),
.A2(n_911),
.B(n_906),
.Y(n_1242)
);

AOI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1090),
.A2(n_1008),
.B(n_882),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1147),
.B(n_969),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1166),
.A2(n_956),
.B1(n_1036),
.B2(n_985),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1064),
.A2(n_985),
.B(n_888),
.C(n_946),
.Y(n_1246)
);

BUFx4_ASAP7_75t_SL g1247 ( 
.A(n_1144),
.Y(n_1247)
);

O2A1O1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1084),
.A2(n_939),
.B(n_923),
.C(n_936),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1074),
.A2(n_932),
.B(n_869),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1181),
.A2(n_1196),
.B(n_1095),
.Y(n_1250)
);

AOI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1105),
.A2(n_923),
.B(n_936),
.Y(n_1251)
);

INVx5_ASAP7_75t_L g1252 ( 
.A(n_1158),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1105),
.A2(n_869),
.B(n_1088),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1082),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1119),
.B(n_946),
.Y(n_1255)
);

AO21x1_ASAP7_75t_L g1256 ( 
.A1(n_1187),
.A2(n_1030),
.B(n_897),
.Y(n_1256)
);

INVxp67_ASAP7_75t_SL g1257 ( 
.A(n_1192),
.Y(n_1257)
);

CKINVDCx11_ASAP7_75t_R g1258 ( 
.A(n_1180),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1108),
.A2(n_1030),
.B(n_1026),
.C(n_981),
.Y(n_1259)
);

AO22x2_ASAP7_75t_L g1260 ( 
.A1(n_1138),
.A2(n_1026),
.B1(n_981),
.B2(n_990),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1162),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1115),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1054),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1118),
.A2(n_869),
.B(n_1030),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1095),
.A2(n_1030),
.B(n_897),
.Y(n_1265)
);

AOI21xp33_ASAP7_75t_L g1266 ( 
.A1(n_1050),
.A2(n_990),
.B(n_1019),
.Y(n_1266)
);

XOR2x2_ASAP7_75t_L g1267 ( 
.A(n_1100),
.B(n_37),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1125),
.A2(n_897),
.B(n_489),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1069),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1081),
.Y(n_1270)
);

A2O1A1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1110),
.A2(n_869),
.B(n_1019),
.C(n_897),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1098),
.B(n_1080),
.Y(n_1272)
);

INVx4_ASAP7_75t_L g1273 ( 
.A(n_1158),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1179),
.A2(n_1186),
.B(n_1117),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1194),
.B(n_1019),
.Y(n_1275)
);

NOR2xp67_ASAP7_75t_L g1276 ( 
.A(n_1047),
.B(n_1019),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1136),
.A2(n_508),
.B(n_512),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1112),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1096),
.A2(n_550),
.B1(n_546),
.B2(n_534),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1161),
.A2(n_508),
.B(n_512),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1148),
.B(n_38),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1093),
.A2(n_521),
.B1(n_489),
.B2(n_512),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1176),
.A2(n_521),
.B(n_489),
.C(n_550),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1160),
.B(n_43),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1106),
.A2(n_1131),
.B(n_1134),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1087),
.B(n_546),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1164),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1128),
.B(n_45),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1054),
.B(n_550),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1063),
.B(n_1173),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1178),
.A2(n_521),
.B(n_546),
.C(n_534),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1093),
.A2(n_521),
.B1(n_512),
.B2(n_508),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1063),
.B(n_108),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_SL g1294 ( 
.A(n_1104),
.B(n_46),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1152),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1139),
.A2(n_508),
.B(n_521),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1182),
.B(n_546),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1168),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1139),
.A2(n_508),
.B(n_546),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1149),
.A2(n_1140),
.B(n_1076),
.Y(n_1300)
);

AOI221x1_ASAP7_75t_L g1301 ( 
.A1(n_1183),
.A2(n_550),
.B1(n_534),
.B2(n_527),
.C(n_49),
.Y(n_1301)
);

OAI21xp33_ASAP7_75t_L g1302 ( 
.A1(n_1184),
.A2(n_550),
.B(n_534),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1140),
.A2(n_534),
.B(n_527),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1169),
.B(n_46),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1127),
.A2(n_97),
.B(n_188),
.Y(n_1305)
);

O2A1O1Ixp5_ASAP7_75t_L g1306 ( 
.A1(n_1170),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_1306)
);

AOI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1101),
.A2(n_534),
.B(n_527),
.Y(n_1307)
);

INVx8_ASAP7_75t_L g1308 ( 
.A(n_1093),
.Y(n_1308)
);

AND2x2_ASAP7_75t_SL g1309 ( 
.A(n_1153),
.B(n_48),
.Y(n_1309)
);

AOI211x1_ASAP7_75t_L g1310 ( 
.A1(n_1097),
.A2(n_50),
.B(n_55),
.C(n_56),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1175),
.B(n_527),
.Y(n_1311)
);

OA21x2_ASAP7_75t_L g1312 ( 
.A1(n_1142),
.A2(n_534),
.B(n_527),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1123),
.Y(n_1313)
);

INVx5_ASAP7_75t_L g1314 ( 
.A(n_1168),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1124),
.A2(n_534),
.B(n_527),
.Y(n_1315)
);

OA21x2_ASAP7_75t_L g1316 ( 
.A1(n_1135),
.A2(n_527),
.B(n_113),
.Y(n_1316)
);

AOI21xp33_ASAP7_75t_L g1317 ( 
.A1(n_1151),
.A2(n_50),
.B(n_56),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1174),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1130),
.A2(n_115),
.B(n_181),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1061),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1124),
.A2(n_61),
.A3(n_66),
.B(n_67),
.Y(n_1321)
);

AOI221x1_ASAP7_75t_L g1322 ( 
.A1(n_1159),
.A2(n_69),
.B1(n_73),
.B2(n_77),
.C(n_83),
.Y(n_1322)
);

AO21x1_ASAP7_75t_L g1323 ( 
.A1(n_1195),
.A2(n_85),
.B(n_96),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1079),
.B(n_106),
.Y(n_1324)
);

AO21x2_ASAP7_75t_L g1325 ( 
.A1(n_1078),
.A2(n_120),
.B(n_126),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1126),
.A2(n_135),
.B(n_141),
.Y(n_1326)
);

A2O1A1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1167),
.A2(n_148),
.B(n_149),
.C(n_157),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1150),
.A2(n_158),
.B(n_161),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1157),
.B(n_168),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1120),
.Y(n_1330)
);

INVx1_ASAP7_75t_SL g1331 ( 
.A(n_1168),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1047),
.Y(n_1332)
);

AOI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1185),
.A2(n_1133),
.B(n_1099),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1141),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1141),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1071),
.B(n_1099),
.Y(n_1336)
);

O2A1O1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1107),
.A2(n_1156),
.B(n_1111),
.C(n_1061),
.Y(n_1337)
);

OR2x6_ASAP7_75t_L g1338 ( 
.A(n_1154),
.B(n_1132),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1171),
.A2(n_1137),
.B(n_1111),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1129),
.A2(n_1075),
.B(n_1091),
.Y(n_1340)
);

INVx4_ASAP7_75t_L g1341 ( 
.A(n_1102),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1102),
.B(n_1132),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1091),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1091),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1075),
.A2(n_1190),
.B(n_1177),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1075),
.B(n_1190),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1190),
.A2(n_1049),
.B(n_940),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1075),
.B(n_1039),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1075),
.B(n_1085),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1075),
.A2(n_1070),
.B1(n_1039),
.B2(n_1092),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_SL g1351 ( 
.A(n_1155),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1048),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1049),
.A2(n_819),
.B(n_838),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1143),
.A2(n_1172),
.B(n_1055),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1213),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1252),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1204),
.A2(n_1350),
.B1(n_1293),
.B2(n_1236),
.Y(n_1357)
);

AO21x2_ASAP7_75t_L g1358 ( 
.A1(n_1347),
.A2(n_1235),
.B(n_1340),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1205),
.B(n_1212),
.Y(n_1359)
);

NOR2xp67_ASAP7_75t_L g1360 ( 
.A(n_1272),
.B(n_1352),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1221),
.Y(n_1361)
);

AO31x2_ASAP7_75t_L g1362 ( 
.A1(n_1343),
.A2(n_1344),
.A3(n_1200),
.B(n_1301),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1290),
.B(n_1209),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1285),
.A2(n_1207),
.B(n_1218),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1349),
.B(n_1293),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1227),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1224),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1234),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1225),
.A2(n_1198),
.B(n_1226),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1353),
.A2(n_1199),
.B(n_1243),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1265),
.A2(n_1249),
.B(n_1305),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1232),
.B(n_1313),
.Y(n_1372)
);

NAND2x1p5_ASAP7_75t_L g1373 ( 
.A(n_1252),
.B(n_1314),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_SL g1374 ( 
.A1(n_1323),
.A2(n_1256),
.B(n_1333),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1223),
.A2(n_1278),
.B1(n_1236),
.B2(n_1257),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1319),
.A2(n_1217),
.B(n_1307),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1347),
.A2(n_1231),
.B(n_1346),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1247),
.Y(n_1378)
);

AOI221x1_ASAP7_75t_L g1379 ( 
.A1(n_1317),
.A2(n_1320),
.B1(n_1260),
.B2(n_1327),
.C(n_1259),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1287),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1264),
.A2(n_1216),
.B(n_1299),
.Y(n_1381)
);

NOR2x1_ASAP7_75t_L g1382 ( 
.A(n_1338),
.B(n_1263),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1348),
.A2(n_1253),
.B(n_1251),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1233),
.A2(n_1241),
.B(n_1280),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1278),
.A2(n_1206),
.B1(n_1271),
.B2(n_1254),
.Y(n_1385)
);

AO21x2_ASAP7_75t_L g1386 ( 
.A1(n_1241),
.A2(n_1233),
.B(n_1303),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1281),
.B(n_1318),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1277),
.A2(n_1296),
.B(n_1315),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1255),
.B(n_1239),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1261),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1302),
.A2(n_1229),
.B1(n_1295),
.B2(n_1270),
.Y(n_1391)
);

OAI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1294),
.A2(n_1322),
.B1(n_1304),
.B2(n_1288),
.Y(n_1392)
);

O2A1O1Ixp33_ASAP7_75t_SL g1393 ( 
.A1(n_1246),
.A2(n_1324),
.B(n_1337),
.C(n_1291),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1284),
.B(n_1309),
.Y(n_1394)
);

NAND2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1252),
.B(n_1314),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1329),
.B(n_1269),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1315),
.A2(n_1345),
.B(n_1303),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1250),
.A2(n_1300),
.B(n_1312),
.Y(n_1398)
);

AO21x2_ASAP7_75t_L g1399 ( 
.A1(n_1300),
.A2(n_1250),
.B(n_1339),
.Y(n_1399)
);

AO31x2_ASAP7_75t_L g1400 ( 
.A1(n_1283),
.A2(n_1330),
.A3(n_1297),
.B(n_1311),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1312),
.A2(n_1242),
.B(n_1248),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1339),
.A2(n_1268),
.B(n_1286),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1244),
.B(n_1237),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1262),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1332),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1229),
.A2(n_1275),
.B1(n_1203),
.B2(n_1245),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1331),
.B(n_1342),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1260),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_SL g1409 ( 
.A1(n_1222),
.A2(n_1310),
.B1(n_1294),
.B2(n_1267),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1268),
.A2(n_1316),
.B(n_1228),
.Y(n_1410)
);

CKINVDCx11_ASAP7_75t_R g1411 ( 
.A(n_1258),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1240),
.A2(n_1316),
.B1(n_1336),
.B2(n_1308),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1334),
.Y(n_1413)
);

AO22x2_ASAP7_75t_L g1414 ( 
.A1(n_1335),
.A2(n_1231),
.B1(n_1289),
.B2(n_1331),
.Y(n_1414)
);

OAI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1229),
.A2(n_1279),
.B1(n_1308),
.B2(n_1197),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1338),
.Y(n_1416)
);

AO21x2_ASAP7_75t_L g1417 ( 
.A1(n_1201),
.A2(n_1279),
.B(n_1219),
.Y(n_1417)
);

AO21x1_ASAP7_75t_L g1418 ( 
.A1(n_1326),
.A2(n_1266),
.B(n_1328),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1308),
.A2(n_1349),
.B1(n_1351),
.B2(n_1228),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1220),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1338),
.A2(n_1325),
.B(n_1224),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1220),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1292),
.A2(n_1282),
.B(n_1306),
.Y(n_1423)
);

AO21x2_ASAP7_75t_L g1424 ( 
.A1(n_1325),
.A2(n_1276),
.B(n_1238),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1341),
.Y(n_1425)
);

AOI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1351),
.A2(n_1237),
.B1(n_1276),
.B2(n_1341),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1208),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1211),
.Y(n_1428)
);

OAI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1314),
.A2(n_1208),
.B1(n_1273),
.B2(n_1298),
.Y(n_1429)
);

AO21x2_ASAP7_75t_L g1430 ( 
.A1(n_1238),
.A2(n_1202),
.B(n_1321),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1211),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1273),
.A2(n_1238),
.B(n_1202),
.Y(n_1432)
);

AOI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1202),
.A2(n_1321),
.B(n_1230),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1321),
.A2(n_1230),
.B(n_1298),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1230),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1298),
.B(n_1284),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1350),
.A2(n_1039),
.B1(n_903),
.B2(n_1049),
.Y(n_1437)
);

CKINVDCx8_ASAP7_75t_R g1438 ( 
.A(n_1203),
.Y(n_1438)
);

OAI221xp5_ASAP7_75t_L g1439 ( 
.A1(n_1350),
.A2(n_1049),
.B1(n_1038),
.B2(n_1039),
.C(n_1015),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1203),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1213),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1213),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1206),
.Y(n_1443)
);

AO31x2_ASAP7_75t_L g1444 ( 
.A1(n_1343),
.A2(n_1344),
.A3(n_1200),
.B(n_1301),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1350),
.A2(n_1049),
.B(n_1038),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1215),
.A2(n_1274),
.B(n_1354),
.Y(n_1446)
);

O2A1O1Ixp33_ASAP7_75t_SL g1447 ( 
.A1(n_1327),
.A2(n_1049),
.B(n_1271),
.C(n_1015),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1224),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1215),
.A2(n_1274),
.B(n_1354),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1284),
.B(n_1204),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1235),
.A2(n_1049),
.B(n_1226),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1350),
.A2(n_1049),
.B(n_1038),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1215),
.A2(n_1274),
.B(n_1354),
.Y(n_1453)
);

CKINVDCx11_ASAP7_75t_R g1454 ( 
.A(n_1258),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1213),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1350),
.A2(n_1039),
.B1(n_903),
.B2(n_1049),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1213),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1205),
.B(n_1039),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1349),
.B(n_1293),
.Y(n_1459)
);

NOR2xp67_ASAP7_75t_L g1460 ( 
.A(n_1272),
.B(n_1080),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1350),
.A2(n_1039),
.B1(n_903),
.B2(n_1049),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1215),
.A2(n_1274),
.B(n_1354),
.Y(n_1462)
);

NAND3xp33_ASAP7_75t_SL g1463 ( 
.A(n_1350),
.B(n_1039),
.C(n_1049),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1213),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1350),
.B(n_1049),
.Y(n_1465)
);

NAND2xp33_ASAP7_75t_SL g1466 ( 
.A(n_1214),
.B(n_1039),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1224),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1205),
.B(n_1039),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1203),
.Y(n_1469)
);

BUFx8_ASAP7_75t_SL g1470 ( 
.A(n_1222),
.Y(n_1470)
);

AO21x2_ASAP7_75t_L g1471 ( 
.A1(n_1347),
.A2(n_1235),
.B(n_1340),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1350),
.A2(n_1049),
.B(n_1038),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1213),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1347),
.A2(n_1200),
.B(n_1210),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1205),
.B(n_1039),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1302),
.A2(n_1049),
.B(n_1015),
.C(n_1092),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1215),
.A2(n_1354),
.B(n_1274),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1290),
.B(n_1205),
.Y(n_1478)
);

OAI222xp33_ASAP7_75t_L g1479 ( 
.A1(n_1350),
.A2(n_1039),
.B1(n_954),
.B2(n_574),
.C1(n_940),
.C2(n_1059),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1260),
.Y(n_1480)
);

CKINVDCx14_ASAP7_75t_R g1481 ( 
.A(n_1222),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1213),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1261),
.Y(n_1483)
);

AO21x2_ASAP7_75t_L g1484 ( 
.A1(n_1347),
.A2(n_1235),
.B(n_1340),
.Y(n_1484)
);

A2O1A1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1302),
.A2(n_1049),
.B(n_1015),
.C(n_1092),
.Y(n_1485)
);

AO22x2_ASAP7_75t_L g1486 ( 
.A1(n_1301),
.A2(n_1347),
.B1(n_1310),
.B2(n_1322),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1260),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1284),
.B(n_1204),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1205),
.B(n_1039),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1347),
.A2(n_1235),
.B(n_1340),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1215),
.A2(n_1274),
.B(n_1354),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1347),
.A2(n_1200),
.B(n_1210),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1235),
.A2(n_1049),
.B(n_1226),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_SL g1494 ( 
.A1(n_1323),
.A2(n_1256),
.B(n_1333),
.Y(n_1494)
);

OA21x2_ASAP7_75t_L g1495 ( 
.A1(n_1347),
.A2(n_1200),
.B(n_1210),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1478),
.B(n_1359),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1363),
.B(n_1458),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1450),
.B(n_1488),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1368),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1445),
.A2(n_1472),
.B(n_1452),
.Y(n_1500)
);

NOR2xp67_ASAP7_75t_L g1501 ( 
.A(n_1460),
.B(n_1360),
.Y(n_1501)
);

OA21x2_ASAP7_75t_L g1502 ( 
.A1(n_1401),
.A2(n_1410),
.B(n_1451),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1468),
.B(n_1475),
.Y(n_1503)
);

OAI31xp33_ASAP7_75t_SL g1504 ( 
.A1(n_1439),
.A2(n_1463),
.A3(n_1456),
.B(n_1437),
.Y(n_1504)
);

AOI21x1_ASAP7_75t_SL g1505 ( 
.A1(n_1396),
.A2(n_1489),
.B(n_1487),
.Y(n_1505)
);

OA21x2_ASAP7_75t_L g1506 ( 
.A1(n_1401),
.A2(n_1410),
.B(n_1493),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1476),
.A2(n_1485),
.B1(n_1392),
.B2(n_1357),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1476),
.A2(n_1485),
.B1(n_1392),
.B2(n_1461),
.Y(n_1508)
);

AOI21x1_ASAP7_75t_SL g1509 ( 
.A1(n_1480),
.A2(n_1487),
.B(n_1420),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1380),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1440),
.Y(n_1511)
);

NOR2xp67_ASAP7_75t_L g1512 ( 
.A(n_1404),
.B(n_1390),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1480),
.Y(n_1513)
);

OA21x2_ASAP7_75t_L g1514 ( 
.A1(n_1432),
.A2(n_1370),
.B(n_1398),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1370),
.A2(n_1398),
.B(n_1384),
.Y(n_1515)
);

AND2x2_ASAP7_75t_SL g1516 ( 
.A(n_1419),
.B(n_1412),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1411),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1389),
.B(n_1372),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1438),
.A2(n_1426),
.B1(n_1382),
.B2(n_1385),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_SL g1520 ( 
.A1(n_1373),
.A2(n_1395),
.B(n_1465),
.Y(n_1520)
);

O2A1O1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1479),
.A2(n_1447),
.B(n_1393),
.C(n_1375),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1387),
.B(n_1407),
.Y(n_1522)
);

OAI31xp33_ASAP7_75t_L g1523 ( 
.A1(n_1409),
.A2(n_1466),
.A3(n_1415),
.B(n_1394),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1365),
.B(n_1459),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1481),
.A2(n_1378),
.B1(n_1483),
.B2(n_1443),
.Y(n_1525)
);

AOI21x1_ASAP7_75t_SL g1526 ( 
.A1(n_1420),
.A2(n_1403),
.B(n_1486),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1469),
.A2(n_1419),
.B1(n_1391),
.B2(n_1406),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1405),
.B(n_1366),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1415),
.A2(n_1481),
.B1(n_1416),
.B2(n_1459),
.Y(n_1529)
);

O2A1O1Ixp5_ASAP7_75t_L g1530 ( 
.A1(n_1418),
.A2(n_1466),
.B(n_1433),
.C(n_1421),
.Y(n_1530)
);

AOI21x1_ASAP7_75t_SL g1531 ( 
.A1(n_1486),
.A2(n_1365),
.B(n_1436),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1441),
.B(n_1455),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_SL g1533 ( 
.A1(n_1373),
.A2(n_1395),
.B(n_1356),
.Y(n_1533)
);

AOI21x1_ASAP7_75t_SL g1534 ( 
.A1(n_1379),
.A2(n_1374),
.B(n_1494),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1455),
.B(n_1464),
.Y(n_1535)
);

INVx3_ASAP7_75t_SL g1536 ( 
.A(n_1378),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_1356),
.Y(n_1537)
);

A2O1A1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1402),
.A2(n_1423),
.B(n_1397),
.C(n_1384),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1411),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1454),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1408),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1355),
.A2(n_1457),
.B1(n_1473),
.B2(n_1442),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1464),
.B(n_1482),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1482),
.B(n_1361),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1428),
.B(n_1435),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1429),
.A2(n_1414),
.B1(n_1425),
.B2(n_1467),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1413),
.B(n_1399),
.Y(n_1547)
);

OA21x2_ASAP7_75t_L g1548 ( 
.A1(n_1397),
.A2(n_1388),
.B(n_1491),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1434),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1367),
.B(n_1467),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1431),
.B(n_1427),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1422),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1425),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1427),
.B(n_1448),
.Y(n_1554)
);

O2A1O1Ixp5_ASAP7_75t_L g1555 ( 
.A1(n_1383),
.A2(n_1422),
.B(n_1429),
.C(n_1448),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1470),
.B(n_1367),
.Y(n_1556)
);

AOI21x1_ASAP7_75t_SL g1557 ( 
.A1(n_1414),
.A2(n_1417),
.B(n_1400),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1470),
.B(n_1356),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1356),
.B(n_1377),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1400),
.B(n_1377),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1454),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1400),
.B(n_1377),
.Y(n_1562)
);

O2A1O1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1386),
.A2(n_1417),
.B(n_1358),
.C(n_1471),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1400),
.B(n_1430),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1474),
.A2(n_1495),
.B1(n_1492),
.B2(n_1386),
.Y(n_1565)
);

AOI21x1_ASAP7_75t_SL g1566 ( 
.A1(n_1424),
.A2(n_1362),
.B(n_1444),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1474),
.A2(n_1495),
.B(n_1492),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1492),
.B(n_1402),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1423),
.A2(n_1490),
.B1(n_1358),
.B2(n_1471),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1484),
.A2(n_1362),
.B1(n_1444),
.B2(n_1376),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1362),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1444),
.A2(n_1376),
.B1(n_1371),
.B2(n_1381),
.Y(n_1572)
);

BUFx5_ASAP7_75t_L g1573 ( 
.A(n_1477),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1446),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1446),
.B(n_1453),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1449),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1449),
.B(n_1462),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1369),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1364),
.B(n_1365),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1368),
.Y(n_1580)
);

O2A1O1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1479),
.A2(n_1049),
.B(n_1439),
.C(n_1445),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1478),
.B(n_1359),
.Y(n_1582)
);

OAI211xp5_ASAP7_75t_L g1583 ( 
.A1(n_1445),
.A2(n_574),
.B(n_954),
.C(n_1038),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1480),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1365),
.B(n_1459),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1363),
.B(n_1387),
.Y(n_1586)
);

AOI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1445),
.A2(n_1049),
.B(n_1452),
.Y(n_1587)
);

CKINVDCx16_ASAP7_75t_R g1588 ( 
.A(n_1481),
.Y(n_1588)
);

AOI21x1_ASAP7_75t_SL g1589 ( 
.A1(n_1396),
.A2(n_1346),
.B(n_1458),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_SL g1590 ( 
.A1(n_1445),
.A2(n_1049),
.B(n_1452),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1363),
.B(n_1387),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1411),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1450),
.B(n_1488),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1365),
.B(n_1459),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1445),
.A2(n_1049),
.B(n_1452),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1363),
.B(n_1387),
.Y(n_1596)
);

OA21x2_ASAP7_75t_L g1597 ( 
.A1(n_1401),
.A2(n_1410),
.B(n_1451),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1450),
.B(n_1488),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_SL g1599 ( 
.A1(n_1445),
.A2(n_1049),
.B(n_1452),
.Y(n_1599)
);

O2A1O1Ixp5_ASAP7_75t_L g1600 ( 
.A1(n_1445),
.A2(n_1472),
.B(n_1452),
.C(n_1049),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1450),
.B(n_1488),
.Y(n_1601)
);

AOI211xp5_ASAP7_75t_L g1602 ( 
.A1(n_1479),
.A2(n_1038),
.B(n_766),
.C(n_1049),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1450),
.B(n_1488),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1478),
.B(n_1359),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1478),
.B(n_1359),
.Y(n_1605)
);

AOI21x1_ASAP7_75t_SL g1606 ( 
.A1(n_1396),
.A2(n_1346),
.B(n_1458),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1450),
.B(n_1488),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1478),
.B(n_1359),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1443),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1541),
.Y(n_1610)
);

OA21x2_ASAP7_75t_L g1611 ( 
.A1(n_1538),
.A2(n_1500),
.B(n_1530),
.Y(n_1611)
);

INVxp33_ASAP7_75t_L g1612 ( 
.A(n_1556),
.Y(n_1612)
);

OR2x6_ASAP7_75t_L g1613 ( 
.A(n_1590),
.B(n_1599),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1541),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1552),
.Y(n_1615)
);

AO21x1_ASAP7_75t_SL g1616 ( 
.A1(n_1571),
.A2(n_1559),
.B(n_1547),
.Y(n_1616)
);

AOI221xp5_ASAP7_75t_L g1617 ( 
.A1(n_1581),
.A2(n_1508),
.B1(n_1602),
.B2(n_1507),
.C(n_1600),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1513),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1513),
.B(n_1584),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1568),
.B(n_1499),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1576),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1552),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1579),
.Y(n_1623)
);

AO31x2_ASAP7_75t_L g1624 ( 
.A1(n_1570),
.A2(n_1569),
.A3(n_1565),
.B(n_1572),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1579),
.B(n_1549),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1584),
.B(n_1560),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_SL g1627 ( 
.A1(n_1583),
.A2(n_1516),
.B1(n_1595),
.B2(n_1587),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1510),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1580),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1577),
.B(n_1574),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1522),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1511),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1528),
.Y(n_1633)
);

OA21x2_ASAP7_75t_L g1634 ( 
.A1(n_1555),
.A2(n_1562),
.B(n_1564),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1516),
.B(n_1544),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1535),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1498),
.B(n_1593),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1575),
.Y(n_1638)
);

OR2x6_ASAP7_75t_L g1639 ( 
.A(n_1520),
.B(n_1563),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1578),
.Y(n_1640)
);

OR2x6_ASAP7_75t_L g1641 ( 
.A(n_1567),
.B(n_1521),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1548),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1566),
.A2(n_1557),
.B(n_1502),
.Y(n_1643)
);

AO21x2_ASAP7_75t_L g1644 ( 
.A1(n_1546),
.A2(n_1527),
.B(n_1542),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_1586),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1598),
.B(n_1601),
.Y(n_1646)
);

OR2x6_ASAP7_75t_L g1647 ( 
.A(n_1533),
.B(n_1529),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1591),
.B(n_1596),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1532),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1548),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1603),
.B(n_1607),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1543),
.Y(n_1652)
);

BUFx12f_ASAP7_75t_L g1653 ( 
.A(n_1517),
.Y(n_1653)
);

OAI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1519),
.A2(n_1588),
.B1(n_1501),
.B2(n_1503),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1515),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1523),
.A2(n_1525),
.B1(n_1497),
.B2(n_1594),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1515),
.Y(n_1657)
);

OAI221xp5_ASAP7_75t_L g1658 ( 
.A1(n_1504),
.A2(n_1496),
.B1(n_1608),
.B2(n_1605),
.C(n_1604),
.Y(n_1658)
);

OAI21x1_ASAP7_75t_L g1659 ( 
.A1(n_1502),
.A2(n_1506),
.B(n_1597),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1514),
.B(n_1545),
.Y(n_1660)
);

OAI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1518),
.A2(n_1512),
.B(n_1582),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1609),
.B(n_1536),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1610),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1657),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1610),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1617),
.A2(n_1627),
.B(n_1613),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1623),
.B(n_1585),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1614),
.Y(n_1668)
);

OAI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1617),
.A2(n_1534),
.B(n_1551),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1660),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1630),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1660),
.B(n_1573),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1653),
.Y(n_1673)
);

CKINVDCx20_ASAP7_75t_R g1674 ( 
.A(n_1653),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1620),
.B(n_1524),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1618),
.Y(n_1676)
);

INVx4_ASAP7_75t_L g1677 ( 
.A(n_1613),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1626),
.B(n_1553),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1633),
.B(n_1554),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1614),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1628),
.Y(n_1681)
);

OR2x6_ASAP7_75t_L g1682 ( 
.A(n_1639),
.B(n_1550),
.Y(n_1682)
);

OAI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1613),
.A2(n_1534),
.B(n_1550),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1619),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1613),
.A2(n_1558),
.B1(n_1536),
.B2(n_1539),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1628),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1638),
.B(n_1537),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1629),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1629),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1638),
.B(n_1526),
.Y(n_1690)
);

INVx3_ASAP7_75t_L g1691 ( 
.A(n_1655),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1619),
.B(n_1509),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1638),
.B(n_1509),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1621),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1623),
.B(n_1531),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1624),
.B(n_1634),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_1625),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1624),
.B(n_1589),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1636),
.B(n_1606),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1636),
.B(n_1505),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1630),
.B(n_1531),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1680),
.Y(n_1702)
);

OAI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1666),
.A2(n_1613),
.B1(n_1658),
.B2(n_1661),
.C(n_1656),
.Y(n_1703)
);

NAND3xp33_ASAP7_75t_L g1704 ( 
.A(n_1666),
.B(n_1658),
.C(n_1661),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1680),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1667),
.B(n_1625),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_SL g1707 ( 
.A1(n_1677),
.A2(n_1644),
.B1(n_1641),
.B2(n_1647),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1664),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1681),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1694),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1675),
.B(n_1631),
.Y(n_1711)
);

OR2x6_ASAP7_75t_L g1712 ( 
.A(n_1682),
.B(n_1639),
.Y(n_1712)
);

AOI33xp33_ASAP7_75t_L g1713 ( 
.A1(n_1685),
.A2(n_1654),
.A3(n_1631),
.B1(n_1635),
.B2(n_1651),
.B3(n_1637),
.Y(n_1713)
);

NOR3xp33_ASAP7_75t_L g1714 ( 
.A(n_1669),
.B(n_1662),
.C(n_1645),
.Y(n_1714)
);

NAND4xp25_ASAP7_75t_L g1715 ( 
.A(n_1669),
.B(n_1648),
.C(n_1632),
.D(n_1635),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1664),
.Y(n_1716)
);

OAI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1699),
.A2(n_1612),
.B(n_1641),
.Y(n_1717)
);

OAI33xp33_ASAP7_75t_L g1718 ( 
.A1(n_1692),
.A2(n_1648),
.A3(n_1649),
.B1(n_1652),
.B2(n_1615),
.B3(n_1622),
.Y(n_1718)
);

AOI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1682),
.A2(n_1639),
.B(n_1641),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1679),
.B(n_1632),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1679),
.B(n_1632),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1676),
.B(n_1700),
.Y(n_1722)
);

OR2x6_ASAP7_75t_L g1723 ( 
.A(n_1682),
.B(n_1639),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1681),
.Y(n_1724)
);

AOI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1696),
.A2(n_1646),
.B1(n_1651),
.B2(n_1637),
.C(n_1644),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1686),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_R g1727 ( 
.A(n_1674),
.B(n_1540),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1675),
.B(n_1623),
.Y(n_1728)
);

OA21x2_ASAP7_75t_L g1729 ( 
.A1(n_1696),
.A2(n_1659),
.B(n_1642),
.Y(n_1729)
);

AOI221x1_ASAP7_75t_SL g1730 ( 
.A1(n_1663),
.A2(n_1652),
.B1(n_1649),
.B2(n_1630),
.C(n_1625),
.Y(n_1730)
);

INVx3_ASAP7_75t_L g1731 ( 
.A(n_1697),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1677),
.A2(n_1647),
.B1(n_1644),
.B2(n_1641),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1686),
.Y(n_1733)
);

AOI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1677),
.A2(n_1647),
.B1(n_1644),
.B2(n_1641),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_R g1735 ( 
.A(n_1674),
.B(n_1561),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1688),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1675),
.B(n_1640),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1676),
.B(n_1684),
.Y(n_1738)
);

OAI21xp33_ASAP7_75t_L g1739 ( 
.A1(n_1698),
.A2(n_1639),
.B(n_1647),
.Y(n_1739)
);

NOR2x1_ASAP7_75t_SL g1740 ( 
.A(n_1682),
.B(n_1616),
.Y(n_1740)
);

NAND2xp33_ASAP7_75t_R g1741 ( 
.A(n_1673),
.B(n_1640),
.Y(n_1741)
);

OAI322xp33_ASAP7_75t_L g1742 ( 
.A1(n_1696),
.A2(n_1692),
.A3(n_1670),
.B1(n_1698),
.B2(n_1665),
.C1(n_1663),
.C2(n_1668),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1688),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1689),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1670),
.B(n_1625),
.Y(n_1745)
);

BUFx3_ASAP7_75t_L g1746 ( 
.A(n_1673),
.Y(n_1746)
);

BUFx3_ASAP7_75t_L g1747 ( 
.A(n_1687),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1709),
.Y(n_1748)
);

INVxp67_ASAP7_75t_SL g1749 ( 
.A(n_1741),
.Y(n_1749)
);

INVx4_ASAP7_75t_SL g1750 ( 
.A(n_1746),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1724),
.Y(n_1751)
);

INVx3_ASAP7_75t_L g1752 ( 
.A(n_1729),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1726),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1704),
.A2(n_1703),
.B(n_1714),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1706),
.B(n_1671),
.Y(n_1755)
);

NAND3xp33_ASAP7_75t_L g1756 ( 
.A(n_1714),
.B(n_1692),
.C(n_1685),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1733),
.Y(n_1757)
);

INVx2_ASAP7_75t_SL g1758 ( 
.A(n_1706),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1729),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_1727),
.Y(n_1760)
);

INVx1_ASAP7_75t_SL g1761 ( 
.A(n_1727),
.Y(n_1761)
);

OA21x2_ASAP7_75t_L g1762 ( 
.A1(n_1739),
.A2(n_1650),
.B(n_1643),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1747),
.B(n_1671),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1736),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1743),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_1746),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1740),
.B(n_1695),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1744),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1702),
.Y(n_1769)
);

OAI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1707),
.A2(n_1683),
.B(n_1693),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1717),
.A2(n_1683),
.B(n_1693),
.Y(n_1771)
);

INVxp67_ASAP7_75t_SL g1772 ( 
.A(n_1741),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1705),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1710),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1738),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1708),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1722),
.B(n_1684),
.Y(n_1777)
);

INVxp67_ASAP7_75t_L g1778 ( 
.A(n_1720),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1730),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1713),
.B(n_1677),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_L g1781 ( 
.A(n_1725),
.B(n_1693),
.C(n_1611),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1716),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1749),
.B(n_1731),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1772),
.B(n_1731),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1777),
.B(n_1715),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1769),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1769),
.Y(n_1787)
);

NAND2xp33_ASAP7_75t_SL g1788 ( 
.A(n_1766),
.B(n_1735),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1767),
.B(n_1747),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1777),
.B(n_1745),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1779),
.B(n_1678),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1767),
.B(n_1728),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_1766),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1775),
.B(n_1774),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1754),
.B(n_1713),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1767),
.B(n_1712),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1748),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1774),
.B(n_1678),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1748),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1778),
.B(n_1711),
.Y(n_1800)
);

INVx2_ASAP7_75t_SL g1801 ( 
.A(n_1766),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1752),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1756),
.B(n_1721),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1766),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1767),
.B(n_1712),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1752),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1751),
.Y(n_1807)
);

NOR3xp33_ASAP7_75t_L g1808 ( 
.A(n_1781),
.B(n_1718),
.C(n_1677),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1773),
.B(n_1665),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1750),
.B(n_1712),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1760),
.Y(n_1811)
);

OAI21x1_ASAP7_75t_L g1812 ( 
.A1(n_1752),
.A2(n_1691),
.B(n_1719),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1751),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1780),
.B(n_1737),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1758),
.B(n_1723),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1752),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1759),
.Y(n_1817)
);

AND2x4_ASAP7_75t_SL g1818 ( 
.A(n_1766),
.B(n_1682),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1758),
.B(n_1723),
.Y(n_1819)
);

NOR2xp33_ASAP7_75t_SL g1820 ( 
.A(n_1761),
.B(n_1653),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1750),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1766),
.B(n_1672),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1773),
.Y(n_1823)
);

OAI31xp33_ASAP7_75t_L g1824 ( 
.A1(n_1763),
.A2(n_1690),
.A3(n_1701),
.B(n_1695),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1786),
.Y(n_1825)
);

AOI21xp33_ASAP7_75t_L g1826 ( 
.A1(n_1795),
.A2(n_1771),
.B(n_1770),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1797),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1797),
.Y(n_1828)
);

AOI221xp5_ASAP7_75t_L g1829 ( 
.A1(n_1808),
.A2(n_1803),
.B1(n_1788),
.B2(n_1811),
.C(n_1804),
.Y(n_1829)
);

INVx1_ASAP7_75t_SL g1830 ( 
.A(n_1811),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1783),
.B(n_1750),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1787),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1823),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1783),
.B(n_1750),
.Y(n_1834)
);

NAND3xp33_ASAP7_75t_L g1835 ( 
.A(n_1791),
.B(n_1734),
.C(n_1732),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1799),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1791),
.B(n_1753),
.Y(n_1837)
);

OAI221xp5_ASAP7_75t_L g1838 ( 
.A1(n_1820),
.A2(n_1682),
.B1(n_1762),
.B2(n_1592),
.C(n_1765),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1784),
.B(n_1750),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1793),
.B(n_1753),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1799),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1784),
.B(n_1755),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1807),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1789),
.B(n_1763),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1802),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1793),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1801),
.B(n_1757),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1801),
.B(n_1757),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1789),
.B(n_1764),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1785),
.B(n_1764),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1807),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1814),
.B(n_1765),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_SL g1853 ( 
.A(n_1820),
.B(n_1742),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1813),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1813),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1792),
.B(n_1768),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1800),
.B(n_1768),
.Y(n_1857)
);

HB1xp67_ASAP7_75t_L g1858 ( 
.A(n_1794),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1785),
.B(n_1776),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1809),
.Y(n_1860)
);

NOR2x1_ASAP7_75t_L g1861 ( 
.A(n_1821),
.B(n_1782),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1858),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1831),
.B(n_1810),
.Y(n_1863)
);

CKINVDCx16_ASAP7_75t_R g1864 ( 
.A(n_1830),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1831),
.B(n_1810),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1826),
.B(n_1842),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1834),
.B(n_1810),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1842),
.B(n_1822),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1836),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1836),
.Y(n_1870)
);

AND2x4_ASAP7_75t_SL g1871 ( 
.A(n_1834),
.B(n_1839),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1841),
.Y(n_1872)
);

INVx1_ASAP7_75t_SL g1873 ( 
.A(n_1839),
.Y(n_1873)
);

INVx1_ASAP7_75t_SL g1874 ( 
.A(n_1850),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1844),
.B(n_1810),
.Y(n_1875)
);

INVxp67_ASAP7_75t_L g1876 ( 
.A(n_1853),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1841),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1861),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1837),
.B(n_1850),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1837),
.B(n_1794),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1844),
.Y(n_1881)
);

INVx2_ASAP7_75t_SL g1882 ( 
.A(n_1846),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1859),
.B(n_1790),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_SL g1884 ( 
.A1(n_1835),
.A2(n_1818),
.B1(n_1805),
.B2(n_1796),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1829),
.B(n_1790),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1859),
.B(n_1798),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1849),
.B(n_1796),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1856),
.B(n_1792),
.Y(n_1888)
);

INVxp67_ASAP7_75t_L g1889 ( 
.A(n_1882),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1879),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1879),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1864),
.B(n_1857),
.Y(n_1892)
);

AOI221xp5_ASAP7_75t_L g1893 ( 
.A1(n_1876),
.A2(n_1825),
.B1(n_1833),
.B2(n_1832),
.C(n_1838),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1873),
.B(n_1825),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1871),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1881),
.B(n_1852),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1874),
.B(n_1832),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1871),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1882),
.B(n_1833),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1880),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1880),
.Y(n_1901)
);

INVxp67_ASAP7_75t_L g1902 ( 
.A(n_1862),
.Y(n_1902)
);

HB1xp67_ASAP7_75t_L g1903 ( 
.A(n_1878),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1866),
.B(n_1885),
.Y(n_1904)
);

O2A1O1Ixp33_ASAP7_75t_L g1905 ( 
.A1(n_1862),
.A2(n_1878),
.B(n_1870),
.C(n_1872),
.Y(n_1905)
);

NAND3xp33_ASAP7_75t_L g1906 ( 
.A(n_1884),
.B(n_1827),
.C(n_1828),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1869),
.Y(n_1907)
);

OA21x2_ASAP7_75t_L g1908 ( 
.A1(n_1869),
.A2(n_1845),
.B(n_1802),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1881),
.B(n_1849),
.Y(n_1909)
);

NAND2x1_ASAP7_75t_L g1910 ( 
.A(n_1875),
.B(n_1860),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1895),
.B(n_1863),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1904),
.B(n_1863),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1903),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1910),
.Y(n_1914)
);

INVx1_ASAP7_75t_SL g1915 ( 
.A(n_1898),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1889),
.B(n_1865),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1903),
.Y(n_1917)
);

NOR2x1p5_ASAP7_75t_L g1918 ( 
.A(n_1899),
.B(n_1865),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1908),
.Y(n_1919)
);

HB1xp67_ASAP7_75t_L g1920 ( 
.A(n_1889),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1892),
.A2(n_1867),
.B1(n_1875),
.B2(n_1887),
.Y(n_1921)
);

NAND2x1_ASAP7_75t_L g1922 ( 
.A(n_1890),
.B(n_1867),
.Y(n_1922)
);

NAND2x1p5_ASAP7_75t_L g1923 ( 
.A(n_1891),
.B(n_1883),
.Y(n_1923)
);

NAND3xp33_ASAP7_75t_SL g1924 ( 
.A(n_1923),
.B(n_1893),
.C(n_1905),
.Y(n_1924)
);

OAI211xp5_ASAP7_75t_L g1925 ( 
.A1(n_1920),
.A2(n_1905),
.B(n_1902),
.C(n_1906),
.Y(n_1925)
);

A2O1A1Ixp33_ASAP7_75t_L g1926 ( 
.A1(n_1912),
.A2(n_1902),
.B(n_1897),
.C(n_1901),
.Y(n_1926)
);

OAI211xp5_ASAP7_75t_L g1927 ( 
.A1(n_1922),
.A2(n_1894),
.B(n_1900),
.C(n_1909),
.Y(n_1927)
);

AOI221xp5_ASAP7_75t_SL g1928 ( 
.A1(n_1921),
.A2(n_1907),
.B1(n_1896),
.B2(n_1868),
.C(n_1877),
.Y(n_1928)
);

NAND4xp25_ASAP7_75t_L g1929 ( 
.A(n_1921),
.B(n_1887),
.C(n_1883),
.D(n_1877),
.Y(n_1929)
);

OAI221xp5_ASAP7_75t_L g1930 ( 
.A1(n_1923),
.A2(n_1886),
.B1(n_1824),
.B2(n_1851),
.C(n_1854),
.Y(n_1930)
);

OAI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1915),
.A2(n_1887),
.B1(n_1888),
.B2(n_1886),
.Y(n_1931)
);

OAI21xp33_ASAP7_75t_L g1932 ( 
.A1(n_1912),
.A2(n_1888),
.B(n_1872),
.Y(n_1932)
);

NOR3xp33_ASAP7_75t_L g1933 ( 
.A(n_1911),
.B(n_1870),
.C(n_1843),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1916),
.B(n_1735),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1924),
.A2(n_1914),
.B(n_1919),
.Y(n_1935)
);

OAI221xp5_ASAP7_75t_L g1936 ( 
.A1(n_1925),
.A2(n_1914),
.B1(n_1913),
.B2(n_1917),
.C(n_1919),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1934),
.Y(n_1937)
);

NAND3xp33_ASAP7_75t_L g1938 ( 
.A(n_1926),
.B(n_1916),
.C(n_1908),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1931),
.Y(n_1939)
);

OAI31xp33_ASAP7_75t_L g1940 ( 
.A1(n_1930),
.A2(n_1927),
.A3(n_1918),
.B(n_1929),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1935),
.B(n_1916),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1936),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1938),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1937),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1939),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1940),
.B(n_1932),
.Y(n_1946)
);

AND2x2_ASAP7_75t_SL g1947 ( 
.A(n_1941),
.B(n_1933),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1941),
.B(n_1860),
.Y(n_1948)
);

OAI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1943),
.A2(n_1848),
.B1(n_1840),
.B2(n_1847),
.Y(n_1949)
);

AOI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1946),
.A2(n_1928),
.B1(n_1855),
.B2(n_1843),
.Y(n_1950)
);

OAI211xp5_ASAP7_75t_L g1951 ( 
.A1(n_1942),
.A2(n_1855),
.B(n_1845),
.C(n_1824),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1948),
.Y(n_1952)
);

NAND4xp75_ASAP7_75t_L g1953 ( 
.A(n_1947),
.B(n_1945),
.C(n_1944),
.D(n_1802),
.Y(n_1953)
);

BUFx3_ASAP7_75t_L g1954 ( 
.A(n_1950),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_SL g1955 ( 
.A1(n_1952),
.A2(n_1949),
.B1(n_1951),
.B2(n_1806),
.Y(n_1955)
);

NAND3xp33_ASAP7_75t_SL g1956 ( 
.A(n_1955),
.B(n_1953),
.C(n_1954),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1956),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1956),
.Y(n_1958)
);

AOI21xp5_ASAP7_75t_L g1959 ( 
.A1(n_1957),
.A2(n_1958),
.B(n_1954),
.Y(n_1959)
);

AOI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1957),
.A2(n_1806),
.B(n_1816),
.Y(n_1960)
);

INVx4_ASAP7_75t_L g1961 ( 
.A(n_1959),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1960),
.B(n_1806),
.Y(n_1962)
);

OAI22xp5_ASAP7_75t_SL g1963 ( 
.A1(n_1961),
.A2(n_1816),
.B1(n_1817),
.B2(n_1798),
.Y(n_1963)
);

OAI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1963),
.A2(n_1962),
.B(n_1816),
.Y(n_1964)
);

OAI21x1_ASAP7_75t_L g1965 ( 
.A1(n_1964),
.A2(n_1817),
.B(n_1856),
.Y(n_1965)
);

OAI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1965),
.A2(n_1817),
.B(n_1812),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1966),
.A2(n_1805),
.B1(n_1819),
.B2(n_1815),
.Y(n_1967)
);

AOI211xp5_ASAP7_75t_L g1968 ( 
.A1(n_1967),
.A2(n_1812),
.B(n_1819),
.C(n_1815),
.Y(n_1968)
);


endmodule