module fake_jpeg_1904_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_56),
.B(n_58),
.Y(n_63)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_1),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_2),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_61),
.Y(n_62)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_63),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_43),
.B1(n_47),
.B2(n_53),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_70),
.B1(n_52),
.B2(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_58),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_38),
.B1(n_47),
.B2(n_46),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_68),
.A2(n_55),
.B(n_61),
.C(n_60),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_38),
.B1(n_50),
.B2(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_81),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_82),
.Y(n_96)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

AO21x2_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_83),
.B(n_68),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_40),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_39),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_44),
.B1(n_4),
.B2(n_5),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_86),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_17),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_3),
.Y(n_98)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_103),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_71),
.C(n_68),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_101),
.C(n_86),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_16),
.B(n_34),
.C(n_33),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_9),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_36),
.C(n_32),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_4),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_5),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_96),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_106),
.B(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_75),
.B1(n_7),
.B2(n_8),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_110),
.B1(n_121),
.B2(n_92),
.Y(n_129)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_26),
.C(n_25),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_114),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_6),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_22),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_116),
.A2(n_118),
.B(n_119),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_10),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_18),
.C(n_19),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_104),
.A2(n_93),
.B(n_98),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_122),
.A2(n_129),
.B(n_132),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_134),
.C(n_135),
.Y(n_138)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

A2O1A1O1Ixp25_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_108),
.B(n_113),
.C(n_106),
.D(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_124),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_137),
.A2(n_127),
.B(n_124),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_140),
.B(n_129),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_138),
.A2(n_123),
.B(n_132),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_141),
.B(n_142),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_126),
.B(n_128),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_112),
.C(n_119),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_12),
.B(n_13),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_15),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_15),
.Y(n_148)
);


endmodule