module fake_netlist_6_1367_n_728 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_728);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_728;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_449;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_532;
wire n_535;
wire n_691;
wire n_544;
wire n_372;
wire n_468;
wire n_250;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_611;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_692;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_404;
wire n_271;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_681;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_427;
wire n_288;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

INVx2_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_140),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_68),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_13),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_91),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_87),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_184),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_58),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_139),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_47),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_93),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_26),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_3),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_187),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_127),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_83),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_132),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_116),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_161),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_144),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_35),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_27),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_142),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_60),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_64),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_8),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_109),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_112),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_157),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_24),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_17),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_178),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_41),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_30),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_118),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_171),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_44),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_40),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_23),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_19),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_65),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_95),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_155),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_100),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_88),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_121),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_143),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_56),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_101),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_8),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_166),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_148),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_0),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_173),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_131),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_51),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_1),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_183),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_129),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_158),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_43),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_42),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_94),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_81),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_150),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_75),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_119),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_72),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_162),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_82),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_160),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_164),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_70),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_124),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_71),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_92),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_114),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_59),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_181),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_98),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_103),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_50),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_32),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_104),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_2),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_9),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_28),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_137),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_165),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_113),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_49),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_43),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_23),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_61),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_107),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_45),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_152),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_90),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_74),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_32),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_26),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_172),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_105),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_15),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_4),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_57),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_24),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_159),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_69),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_29),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_18),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_46),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_167),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_135),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_108),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_138),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_84),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_79),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_20),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_190),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_204),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_203),
.Y(n_317)
);

INVxp33_ASAP7_75t_SL g318 ( 
.A(n_270),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_196),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_213),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_230),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_214),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_197),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_225),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_194),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_226),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_198),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_232),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_243),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_255),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_208),
.Y(n_331)
);

BUFx6f_ASAP7_75t_SL g332 ( 
.A(n_256),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_279),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_231),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_280),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_200),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_205),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_287),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_206),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_210),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_313),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_196),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_201),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_201),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_193),
.B(n_2),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_212),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_281),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_241),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_295),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_216),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_221),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_285),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_300),
.B(n_5),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_302),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_218),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_224),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_228),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_192),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_202),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_207),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_222),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_209),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_223),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_229),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_211),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_215),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_251),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_236),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_238),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_217),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_244),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_219),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_195),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_241),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_227),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_233),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_268),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_248),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_234),
.B(n_6),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_249),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_252),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_237),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_240),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_242),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_253),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_245),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_254),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_241),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_195),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_257),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_258),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_259),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_277),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_247),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_261),
.Y(n_397)
);

NOR2xp67_ASAP7_75t_L g398 ( 
.A(n_290),
.B(n_7),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_360),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_317),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_320),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_318),
.B(n_220),
.Y(n_402)
);

AND2x2_ASAP7_75t_SL g403 ( 
.A(n_355),
.B(n_191),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_347),
.B(n_235),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_325),
.B(n_235),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_361),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_396),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_362),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_367),
.B(n_262),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_364),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_314),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_319),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_368),
.Y(n_414)
);

OA21x2_ASAP7_75t_L g415 ( 
.A1(n_381),
.A2(n_269),
.B(n_267),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_356),
.B(n_375),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_324),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_375),
.B(n_189),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_326),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_374),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_319),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_328),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_329),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_330),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_333),
.Y(n_425)
);

BUFx8_ASAP7_75t_L g426 ( 
.A(n_332),
.Y(n_426)
);

OA21x2_ASAP7_75t_L g427 ( 
.A1(n_350),
.A2(n_275),
.B(n_272),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_377),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_335),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_372),
.B(n_263),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_336),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_385),
.B(n_264),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_378),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_388),
.B(n_265),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_395),
.B(n_260),
.Y(n_435)
);

OA21x2_ASAP7_75t_L g436 ( 
.A1(n_350),
.A2(n_278),
.B(n_276),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_339),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_384),
.B(n_266),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_386),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_342),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_343),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_376),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_315),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_344),
.Y(n_444)
);

NAND2xp33_ASAP7_75t_L g445 ( 
.A(n_345),
.B(n_191),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_323),
.B(n_273),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_346),
.B(n_274),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_390),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_354),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_327),
.B(n_337),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_338),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_340),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_341),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_348),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_352),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_353),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_403),
.B(n_410),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_413),
.B(n_398),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_448),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_403),
.B(n_358),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_399),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_407),
.B(n_391),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_448),
.Y(n_463)
);

NAND2x1p5_ASAP7_75t_L g464 ( 
.A(n_454),
.B(n_239),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_406),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_413),
.B(n_283),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_448),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_410),
.B(n_359),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_191),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_442),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_435),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_408),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_411),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_421),
.B(n_284),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_199),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_430),
.B(n_370),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_414),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_449),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_421),
.B(n_371),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_412),
.B(n_331),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_449),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_449),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_416),
.B(n_373),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_449),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_419),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_420),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_419),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_454),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_454),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_430),
.B(n_380),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_419),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_450),
.B(n_382),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_418),
.B(n_444),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_431),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_428),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_433),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_431),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_451),
.B(n_383),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_431),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_447),
.B(n_387),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_400),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_439),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_432),
.B(n_389),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_401),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_432),
.B(n_392),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_434),
.B(n_447),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_455),
.B(n_393),
.Y(n_507)
);

NAND2xp33_ASAP7_75t_L g508 ( 
.A(n_434),
.B(n_394),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_409),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_438),
.B(n_397),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_489),
.Y(n_511)
);

AO22x2_ASAP7_75t_L g512 ( 
.A1(n_457),
.A2(n_402),
.B1(n_404),
.B2(n_405),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_480),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_460),
.B(n_456),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_506),
.B(n_446),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_492),
.B(n_468),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_461),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_465),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_472),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_473),
.Y(n_520)
);

NOR2x1p5_ASAP7_75t_L g521 ( 
.A(n_462),
.B(n_426),
.Y(n_521)
);

AO22x2_ASAP7_75t_L g522 ( 
.A1(n_471),
.A2(n_291),
.B1(n_292),
.B2(n_289),
.Y(n_522)
);

AO22x2_ASAP7_75t_L g523 ( 
.A1(n_510),
.A2(n_306),
.B1(n_307),
.B2(n_297),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_477),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_476),
.B(n_415),
.Y(n_525)
);

AO22x2_ASAP7_75t_L g526 ( 
.A1(n_500),
.A2(n_309),
.B1(n_311),
.B2(n_308),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_490),
.B(n_415),
.Y(n_527)
);

AO22x2_ASAP7_75t_L g528 ( 
.A1(n_483),
.A2(n_321),
.B1(n_334),
.B2(n_316),
.Y(n_528)
);

NOR2xp67_ASAP7_75t_L g529 ( 
.A(n_488),
.B(n_498),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_486),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_470),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_495),
.Y(n_532)
);

NAND2x1p5_ASAP7_75t_L g533 ( 
.A(n_479),
.B(n_429),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_503),
.B(n_415),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_501),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_496),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_502),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_504),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_509),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_505),
.B(n_427),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_458),
.B(n_427),
.Y(n_541)
);

AO22x2_ASAP7_75t_L g542 ( 
.A1(n_466),
.A2(n_351),
.B1(n_349),
.B2(n_357),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_466),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_481),
.Y(n_544)
);

AO22x2_ASAP7_75t_L g545 ( 
.A1(n_474),
.A2(n_365),
.B1(n_366),
.B2(n_363),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_507),
.B(n_363),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_481),
.Y(n_547)
);

AO22x2_ASAP7_75t_L g548 ( 
.A1(n_458),
.A2(n_366),
.B1(n_369),
.B2(n_365),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_482),
.Y(n_549)
);

OAI221xp5_ASAP7_75t_L g550 ( 
.A1(n_508),
.A2(n_425),
.B1(n_417),
.B2(n_422),
.C(n_423),
.Y(n_550)
);

OAI221xp5_ASAP7_75t_L g551 ( 
.A1(n_464),
.A2(n_424),
.B1(n_437),
.B2(n_440),
.C(n_299),
.Y(n_551)
);

OAI221xp5_ASAP7_75t_L g552 ( 
.A1(n_499),
.A2(n_440),
.B1(n_294),
.B2(n_298),
.C(n_305),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_499),
.B(n_427),
.Y(n_553)
);

BUFx8_ASAP7_75t_L g554 ( 
.A(n_469),
.Y(n_554)
);

NAND2x1p5_ASAP7_75t_L g555 ( 
.A(n_494),
.B(n_441),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_516),
.B(n_485),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_515),
.B(n_497),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_529),
.B(n_487),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_511),
.B(n_487),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_511),
.B(n_533),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_513),
.B(n_379),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_SL g562 ( 
.A(n_521),
.B(n_282),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_525),
.B(n_491),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_517),
.B(n_518),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_519),
.B(n_484),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_527),
.B(n_491),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_543),
.B(n_478),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_520),
.B(n_478),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_534),
.B(n_459),
.Y(n_569)
);

AND2x2_ASAP7_75t_SL g570 ( 
.A(n_546),
.B(n_199),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_524),
.B(n_443),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_L g572 ( 
.A(n_541),
.B(n_540),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_514),
.B(n_463),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_530),
.B(n_467),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_532),
.B(n_288),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_536),
.B(n_469),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_537),
.B(n_469),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_531),
.B(n_469),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_535),
.B(n_293),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_538),
.B(n_296),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_539),
.B(n_531),
.Y(n_581)
);

NAND2xp33_ASAP7_75t_SL g582 ( 
.A(n_544),
.B(n_303),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_547),
.B(n_310),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_549),
.B(n_312),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_555),
.B(n_246),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_512),
.B(n_475),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_554),
.B(n_271),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_553),
.B(n_271),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_551),
.B(n_241),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_552),
.B(n_250),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_556),
.B(n_522),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_572),
.A2(n_550),
.B(n_436),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_559),
.Y(n_593)
);

O2A1O1Ixp5_ASAP7_75t_L g594 ( 
.A1(n_589),
.A2(n_522),
.B(n_523),
.C(n_526),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_564),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_581),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_563),
.A2(n_436),
.B(n_445),
.Y(n_597)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_569),
.A2(n_250),
.B(n_523),
.Y(n_598)
);

OAI21x1_ASAP7_75t_L g599 ( 
.A1(n_566),
.A2(n_250),
.B(n_526),
.Y(n_599)
);

OAI21x1_ASAP7_75t_L g600 ( 
.A1(n_573),
.A2(n_250),
.B(n_48),
.Y(n_600)
);

AO31x2_ASAP7_75t_L g601 ( 
.A1(n_586),
.A2(n_578),
.A3(n_558),
.B(n_577),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_570),
.B(n_528),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_567),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_576),
.B(n_250),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_574),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_588),
.A2(n_250),
.B(n_53),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_557),
.A2(n_542),
.B(n_545),
.Y(n_607)
);

OAI21x1_ASAP7_75t_L g608 ( 
.A1(n_568),
.A2(n_54),
.B(n_52),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_560),
.B(n_55),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_575),
.B(n_548),
.Y(n_610)
);

AO31x2_ASAP7_75t_L g611 ( 
.A1(n_590),
.A2(n_10),
.A3(n_11),
.B(n_12),
.Y(n_611)
);

NOR2x1_ASAP7_75t_R g612 ( 
.A(n_561),
.B(n_10),
.Y(n_612)
);

AO31x2_ASAP7_75t_L g613 ( 
.A1(n_585),
.A2(n_14),
.A3(n_15),
.B(n_16),
.Y(n_613)
);

OA21x2_ASAP7_75t_L g614 ( 
.A1(n_571),
.A2(n_63),
.B(n_62),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_587),
.Y(n_615)
);

AOI21x1_ASAP7_75t_L g616 ( 
.A1(n_565),
.A2(n_67),
.B(n_66),
.Y(n_616)
);

AO31x2_ASAP7_75t_L g617 ( 
.A1(n_582),
.A2(n_21),
.A3(n_22),
.B(n_25),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_593),
.B(n_603),
.Y(n_618)
);

OAI21x1_ASAP7_75t_L g619 ( 
.A1(n_592),
.A2(n_606),
.B(n_597),
.Y(n_619)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_600),
.A2(n_584),
.B(n_583),
.Y(n_620)
);

OA21x2_ASAP7_75t_L g621 ( 
.A1(n_598),
.A2(n_580),
.B(n_579),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_596),
.Y(n_622)
);

OAI21x1_ASAP7_75t_L g623 ( 
.A1(n_608),
.A2(n_562),
.B(n_73),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_599),
.A2(n_77),
.B(n_76),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_591),
.A2(n_115),
.B(n_188),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_595),
.Y(n_626)
);

OAI21x1_ASAP7_75t_L g627 ( 
.A1(n_616),
.A2(n_117),
.B(n_186),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_605),
.Y(n_628)
);

OA21x2_ASAP7_75t_L g629 ( 
.A1(n_594),
.A2(n_120),
.B(n_185),
.Y(n_629)
);

AND2x6_ASAP7_75t_L g630 ( 
.A(n_609),
.B(n_78),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_L g631 ( 
.A1(n_604),
.A2(n_122),
.B(n_180),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_602),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_632)
);

OAI21x1_ASAP7_75t_L g633 ( 
.A1(n_614),
.A2(n_123),
.B(n_179),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_615),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_610),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_607),
.B(n_36),
.Y(n_636)
);

AO31x2_ASAP7_75t_L g637 ( 
.A1(n_601),
.A2(n_37),
.A3(n_38),
.B(n_39),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_601),
.A2(n_126),
.B(n_177),
.Y(n_638)
);

OAI21x1_ASAP7_75t_L g639 ( 
.A1(n_611),
.A2(n_111),
.B(n_176),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_612),
.A2(n_110),
.B(n_175),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_613),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_612),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_622),
.Y(n_643)
);

OAI21x1_ASAP7_75t_L g644 ( 
.A1(n_619),
.A2(n_617),
.B(n_613),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_618),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_626),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_641),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_628),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_623),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_637),
.Y(n_650)
);

AO21x2_ASAP7_75t_L g651 ( 
.A1(n_638),
.A2(n_130),
.B(n_170),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_639),
.Y(n_652)
);

OAI21x1_ASAP7_75t_L g653 ( 
.A1(n_624),
.A2(n_128),
.B(n_169),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_633),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_627),
.Y(n_655)
);

INVx8_ASAP7_75t_L g656 ( 
.A(n_630),
.Y(n_656)
);

OAI21x1_ASAP7_75t_L g657 ( 
.A1(n_620),
.A2(n_134),
.B(n_168),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_635),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_636),
.B(n_133),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_634),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_629),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_629),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_621),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_621),
.Y(n_664)
);

OR2x6_ASAP7_75t_L g665 ( 
.A(n_656),
.B(n_640),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_646),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_658),
.B(n_642),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_658),
.B(n_630),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_660),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_659),
.B(n_632),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_643),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_645),
.B(n_625),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_645),
.B(n_625),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_648),
.B(n_631),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_647),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_675),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_666),
.B(n_650),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_671),
.B(n_651),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_670),
.B(n_663),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_674),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_674),
.B(n_663),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_667),
.B(n_664),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_665),
.B(n_644),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_672),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_672),
.B(n_664),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_673),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_668),
.B(n_644),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_665),
.B(n_652),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_678),
.B(n_661),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_676),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_685),
.B(n_661),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_688),
.B(n_683),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_682),
.B(n_662),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_682),
.B(n_662),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_684),
.B(n_649),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_686),
.B(n_649),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_679),
.B(n_669),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_686),
.B(n_654),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_690),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_689),
.B(n_680),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_692),
.B(n_687),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_700),
.B(n_697),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_701),
.B(n_695),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_702),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_703),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_704),
.B(n_699),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_706),
.B(n_705),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_707),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_708),
.A2(n_696),
.B1(n_698),
.B2(n_691),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_709),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_710),
.Y(n_711)
);

NAND2xp33_ASAP7_75t_SL g712 ( 
.A(n_711),
.B(n_694),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_R g713 ( 
.A(n_711),
.B(n_80),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_712),
.A2(n_693),
.B1(n_681),
.B2(n_677),
.Y(n_714)
);

INVx5_ASAP7_75t_L g715 ( 
.A(n_713),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_715),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_715),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_716),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_717),
.Y(n_719)
);

AOI31xp33_ASAP7_75t_L g720 ( 
.A1(n_718),
.A2(n_714),
.A3(n_86),
.B(n_89),
.Y(n_720)
);

AOI31xp33_ASAP7_75t_L g721 ( 
.A1(n_719),
.A2(n_85),
.A3(n_96),
.B(n_97),
.Y(n_721)
);

NOR5xp2_ASAP7_75t_L g722 ( 
.A(n_720),
.B(n_99),
.C(n_102),
.D(n_106),
.E(n_136),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_721),
.A2(n_657),
.B(n_653),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_R g724 ( 
.A1(n_722),
.A2(n_141),
.B1(n_145),
.B2(n_146),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_723),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_725),
.Y(n_726)
);

AOI221xp5_ASAP7_75t_L g727 ( 
.A1(n_726),
.A2(n_724),
.B1(n_147),
.B2(n_149),
.C(n_153),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_727),
.A2(n_677),
.B1(n_681),
.B2(n_655),
.Y(n_728)
);


endmodule