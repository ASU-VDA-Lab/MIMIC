module fake_jpeg_2503_n_45 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_4),
.B(n_0),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx3_ASAP7_75t_SL g9 ( 
.A(n_0),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_1),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_5),
.B(n_6),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_20),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_14),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_17),
.A2(n_2),
.B1(n_5),
.B2(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

AO22x1_ASAP7_75t_SL g19 ( 
.A1(n_11),
.A2(n_9),
.B1(n_13),
.B2(n_8),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_11),
.B(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_7),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_21),
.B(n_22),
.Y(n_24)
);

CKINVDCx12_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_29),
.Y(n_35)
);

MAJx2_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_12),
.C(n_9),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_16),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_19),
.A2(n_10),
.B(n_2),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_17),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_36),
.B(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_25),
.B1(n_26),
.B2(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_34),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_35),
.C(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_42),
.Y(n_43)
);

AOI322xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_39),
.A3(n_38),
.B1(n_37),
.B2(n_24),
.C1(n_20),
.C2(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_38),
.Y(n_45)
);


endmodule