module fake_jpeg_3096_n_160 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_30),
.B(n_27),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_64),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_66),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_42),
.B1(n_55),
.B2(n_49),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_70),
.A2(n_59),
.B1(n_47),
.B2(n_52),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_62),
.B(n_41),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_73),
.Y(n_83)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_80),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_49),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_77),
.A2(n_65),
.B1(n_42),
.B2(n_73),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_87),
.B1(n_92),
.B2(n_59),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_53),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_88),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_63),
.B1(n_52),
.B2(n_57),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_69),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_67),
.A2(n_57),
.B1(n_52),
.B2(n_43),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_90),
.B1(n_40),
.B2(n_46),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_74),
.B1(n_68),
.B2(n_72),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_91),
.B(n_41),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_94),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_103),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_72),
.B1(n_68),
.B2(n_71),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_101),
.B1(n_109),
.B2(n_5),
.Y(n_118)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_89),
.B(n_59),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_24),
.B(n_23),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_71),
.B1(n_43),
.B2(n_69),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_54),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_104),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_0),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_106),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_40),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_17),
.C(n_35),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_46),
.B1(n_2),
.B2(n_3),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_6),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_113),
.C(n_123),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_39),
.Y(n_113)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_34),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_126),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_121),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_6),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_122),
.B(n_127),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_103),
.Y(n_123)
);

OAI22x1_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_28),
.B1(n_26),
.B2(n_25),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_18),
.Y(n_135)
);

AO21x1_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_8),
.B(n_9),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_21),
.B(n_19),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_7),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_135),
.B1(n_139),
.B2(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_138),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_11),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_124),
.B1(n_121),
.B2(n_112),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_143),
.B1(n_135),
.B2(n_130),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_113),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_132),
.C(n_133),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_131),
.A2(n_115),
.B(n_123),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_147),
.B(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_144),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_149),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_150),
.A2(n_151),
.B(n_138),
.C(n_136),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_152),
.A2(n_141),
.B(n_145),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_154),
.B(n_145),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_153),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_149),
.Y(n_157)
);

OAI321xp33_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_129),
.A3(n_146),
.B1(n_120),
.B2(n_114),
.C(n_14),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_120),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_15),
.Y(n_160)
);


endmodule