module fake_jpeg_22258_n_301 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_34),
.B(n_38),
.Y(n_57)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_17),
.Y(n_44)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_28),
.B1(n_29),
.B2(n_17),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_56),
.B(n_18),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_46),
.Y(n_63)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx2_ASAP7_75t_SL g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_52),
.Y(n_60)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_55),
.Y(n_74)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_39),
.B(n_36),
.C(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_62),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_69),
.Y(n_103)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx5_ASAP7_75t_SL g89 ( 
.A(n_61),
.Y(n_89)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_66),
.A2(n_67),
.B1(n_55),
.B2(n_52),
.Y(n_90)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_36),
.B(n_34),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_34),
.C(n_39),
.Y(n_92)
);

AND2x4_ASAP7_75t_SL g69 ( 
.A(n_44),
.B(n_36),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_73),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_75),
.Y(n_98)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_40),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_41),
.B1(n_37),
.B2(n_34),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_77),
.A2(n_79),
.B1(n_80),
.B2(n_55),
.Y(n_109)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_81),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_41),
.B1(n_37),
.B2(n_18),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_51),
.A2(n_41),
.B1(n_37),
.B2(n_25),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_25),
.B1(n_41),
.B2(n_20),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_84),
.Y(n_105)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_100),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_90),
.A2(n_16),
.B1(n_23),
.B2(n_27),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_108),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_86),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_40),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_110),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_75),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_107),
.B(n_58),
.Y(n_124)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_115),
.B1(n_78),
.B2(n_49),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_40),
.Y(n_110)
);

AOI22x1_ASAP7_75t_L g111 ( 
.A1(n_69),
.A2(n_54),
.B1(n_52),
.B2(n_47),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_72),
.B1(n_83),
.B2(n_81),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_54),
.C(n_47),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_62),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_69),
.C(n_63),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_103),
.C(n_96),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_117),
.B(n_139),
.Y(n_156)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_69),
.B(n_66),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_133),
.B(n_138),
.Y(n_144)
);

OAI22x1_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_63),
.B1(n_68),
.B2(n_23),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_125),
.B1(n_126),
.B2(n_128),
.Y(n_146)
);

BUFx24_ASAP7_75t_SL g120 ( 
.A(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_122),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_105),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_124),
.B(n_142),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_72),
.B1(n_61),
.B2(n_31),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_84),
.B1(n_73),
.B2(n_67),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_136),
.B1(n_95),
.B2(n_100),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_94),
.A2(n_32),
.B(n_21),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_107),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_143),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_91),
.A2(n_49),
.B1(n_31),
.B2(n_20),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_112),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_49),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_65),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_95),
.B1(n_89),
.B2(n_113),
.Y(n_150)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_21),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_98),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_172),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_106),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_158),
.C(n_166),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_171),
.B1(n_139),
.B2(n_117),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_165),
.B1(n_125),
.B2(n_136),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_92),
.B(n_103),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_153),
.Y(n_198)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_161),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_95),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_159),
.B(n_162),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_103),
.B(n_96),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_88),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_130),
.B(n_108),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_163),
.B(n_164),
.Y(n_190)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_119),
.A2(n_93),
.B1(n_101),
.B2(n_32),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_93),
.C(n_65),
.Y(n_166)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_23),
.Y(n_169)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_173),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_118),
.A2(n_33),
.B1(n_26),
.B2(n_24),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_23),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_116),
.B(n_99),
.C(n_33),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_27),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_176),
.A2(n_192),
.B1(n_196),
.B2(n_199),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_189),
.Y(n_218)
);

BUFx4f_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_157),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_181),
.B(n_203),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_144),
.A2(n_133),
.B(n_118),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_183),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_123),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_186),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_122),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_172),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_187),
.A2(n_197),
.B(n_175),
.Y(n_225)
);

XNOR2x2_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_121),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_188),
.B(n_178),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_26),
.B1(n_24),
.B2(n_22),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_204),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_146),
.A2(n_22),
.B1(n_99),
.B2(n_27),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_9),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_27),
.B1(n_99),
.B2(n_2),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_200)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_10),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_174),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_154),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_166),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_151),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_207),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_160),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_223),
.C(n_202),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_168),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_213),
.B(n_219),
.Y(n_234)
);

OA21x2_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_150),
.B(n_156),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_201),
.B(n_193),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_155),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_186),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_152),
.Y(n_216)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_153),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_222),
.B(n_224),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_147),
.Y(n_223)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_191),
.B(n_168),
.CI(n_170),
.CON(n_224),
.SN(n_224)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_225),
.B(n_200),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_236),
.B1(n_204),
.B2(n_206),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_233),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_231),
.A2(n_214),
.B1(n_218),
.B2(n_222),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_210),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_235),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_179),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_209),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_196),
.B1(n_177),
.B2(n_192),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_239),
.C(n_241),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_187),
.C(n_179),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_197),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_189),
.C(n_195),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_221),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_224),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_244),
.A2(n_256),
.B1(n_239),
.B2(n_224),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_257),
.B1(n_230),
.B2(n_180),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_234),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_252),
.Y(n_266)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_228),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_215),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_211),
.C(n_212),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_251),
.C(n_238),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_237),
.A2(n_240),
.B1(n_214),
.B2(n_208),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_205),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_227),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_227),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_260),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_229),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_261),
.B(n_267),
.Y(n_275)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_233),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_265),
.A2(n_269),
.B(n_270),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_253),
.B1(n_249),
.B2(n_250),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_173),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_279),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_251),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_277),
.B(n_278),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_264),
.A2(n_252),
.B(n_246),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_11),
.B(n_14),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_11),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_260),
.Y(n_281)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_274),
.A2(n_265),
.B(n_263),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_288),
.B(n_271),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_11),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_283),
.B(n_286),
.Y(n_293)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_279),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_275),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_3),
.C(n_6),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_284),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_291),
.A2(n_292),
.B(n_8),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_12),
.B(n_14),
.Y(n_292)
);

OAI321xp33_ASAP7_75t_L g297 ( 
.A1(n_294),
.A2(n_295),
.A3(n_296),
.B1(n_10),
.B2(n_12),
.C(n_13),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_289),
.A2(n_288),
.B(n_293),
.Y(n_295)
);

A2O1A1Ixp33_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_12),
.B(n_15),
.C(n_3),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_15),
.B(n_7),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_7),
.B(n_298),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_300),
.B(n_7),
.Y(n_301)
);


endmodule