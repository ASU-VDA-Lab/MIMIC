module fake_ariane_710_n_864 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_864);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_864;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_779;
wire n_731;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_553;
wire n_446;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_821;
wire n_218;
wire n_839;
wire n_770;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_365;
wire n_238;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_861;
wire n_780;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_747;
wire n_772;
wire n_741;
wire n_847;
wire n_371;
wire n_845;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_8),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_47),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_135),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_72),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_23),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_92),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_129),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_53),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_52),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_42),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_97),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_120),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_117),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_115),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_74),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_3),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_28),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_109),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_151),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_1),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_60),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_67),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_11),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_14),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_107),
.Y(n_217)
);

NOR2xp67_ASAP7_75t_L g218 ( 
.A(n_16),
.B(n_167),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_40),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_37),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_9),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_57),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_122),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_138),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_45),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_25),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_146),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_26),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_101),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_144),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_34),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_73),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_66),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_18),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_181),
.B(n_171),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_14),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_112),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_76),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_12),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_145),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_8),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_125),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_108),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_156),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_71),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_39),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_55),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_153),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_136),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_21),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_49),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_184),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_189),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_224),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_193),
.Y(n_256)
);

OAI21x1_ASAP7_75t_L g257 ( 
.A1(n_188),
.A2(n_89),
.B(n_182),
.Y(n_257)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_193),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_193),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_193),
.Y(n_260)
);

AND2x4_ASAP7_75t_L g261 ( 
.A(n_215),
.B(n_0),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_190),
.Y(n_262)
);

OA22x2_ASAP7_75t_L g263 ( 
.A1(n_221),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_236),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g265 ( 
.A(n_185),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_192),
.B(n_5),
.Y(n_266)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_223),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_194),
.B(n_6),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_195),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_239),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_199),
.B(n_7),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_200),
.Y(n_272)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_223),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_220),
.B(n_7),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_247),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_248),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_207),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_223),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_203),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_204),
.Y(n_280)
);

AND2x4_ASAP7_75t_L g281 ( 
.A(n_208),
.B(n_9),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_226),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_223),
.Y(n_283)
);

BUFx8_ASAP7_75t_SL g284 ( 
.A(n_216),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_241),
.Y(n_285)
);

CKINVDCx6p67_ASAP7_75t_R g286 ( 
.A(n_211),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_186),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_230),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_232),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_233),
.Y(n_291)
);

OA21x2_ASAP7_75t_L g292 ( 
.A1(n_242),
.A2(n_10),
.B(n_11),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_217),
.B(n_10),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_220),
.B(n_12),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_228),
.B(n_13),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_228),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_228),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_228),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_187),
.Y(n_299)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_196),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_197),
.Y(n_301)
);

NOR2xp67_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_235),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_286),
.B(n_191),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_275),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_285),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_276),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_284),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_258),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_284),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_262),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_265),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_265),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_300),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_262),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_264),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_272),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_252),
.B(n_231),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_300),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_300),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_296),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_279),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_300),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_299),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_279),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_L g329 ( 
.A(n_274),
.B(n_198),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_253),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_299),
.Y(n_332)
);

NAND2xp33_ASAP7_75t_R g333 ( 
.A(n_294),
.B(n_201),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_290),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_297),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_256),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_258),
.B(n_202),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_301),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_205),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_253),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_297),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_269),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_256),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_269),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_255),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_252),
.B(n_206),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_291),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_256),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_281),
.B(n_209),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_287),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_270),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_287),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_280),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_282),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_354),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_313),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_306),
.Y(n_358)
);

NOR3xp33_ASAP7_75t_L g359 ( 
.A(n_305),
.B(n_271),
.C(n_268),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_281),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_353),
.B(n_270),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_289),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_340),
.B(n_281),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_308),
.B(n_263),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_312),
.B(n_295),
.Y(n_365)
);

AO221x1_ASAP7_75t_L g366 ( 
.A1(n_333),
.A2(n_263),
.B1(n_277),
.B2(n_261),
.C(n_292),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_303),
.B(n_295),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_313),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_317),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_319),
.Y(n_370)
);

NOR2xp67_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_295),
.Y(n_371)
);

NAND2x1_ASAP7_75t_L g372 ( 
.A(n_320),
.B(n_292),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_342),
.B(n_261),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_328),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_293),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_325),
.B(n_258),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_344),
.B(n_266),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_351),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_266),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_328),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_331),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_350),
.B(n_268),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_333),
.A2(n_246),
.B1(n_213),
.B2(n_214),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_348),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_321),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_334),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_352),
.A2(n_292),
.B1(n_277),
.B2(n_210),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_345),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_258),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_330),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_347),
.B(n_267),
.Y(n_392)
);

AND2x6_ASAP7_75t_SL g393 ( 
.A(n_309),
.B(n_13),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_350),
.B(n_267),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_302),
.B(n_219),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_304),
.B(n_267),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_311),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_304),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_324),
.B(n_267),
.Y(n_399)
);

AO221x1_ASAP7_75t_L g400 ( 
.A1(n_318),
.A2(n_298),
.B1(n_283),
.B2(n_278),
.C(n_260),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_324),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_335),
.B(n_273),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_315),
.B(n_222),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_335),
.Y(n_404)
);

BUFx6f_ASAP7_75t_SL g405 ( 
.A(n_307),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_314),
.B(n_225),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_316),
.B(n_273),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_341),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_322),
.B(n_323),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_341),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_343),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_336),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_326),
.B(n_227),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_343),
.B(n_273),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_349),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_349),
.B(n_273),
.Y(n_416)
);

BUFx5_ASAP7_75t_L g417 ( 
.A(n_310),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_336),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_336),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_337),
.B(n_310),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_352),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_346),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_422),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_361),
.B(n_346),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_357),
.Y(n_426)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_412),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_368),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_397),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_375),
.A2(n_360),
.B1(n_367),
.B2(n_362),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_374),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_378),
.Y(n_432)
);

BUFx8_ASAP7_75t_L g433 ( 
.A(n_405),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_380),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_384),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_360),
.B(n_229),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_390),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_412),
.Y(n_438)
);

CKINVDCx8_ASAP7_75t_R g439 ( 
.A(n_393),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_355),
.B(n_257),
.Y(n_440)
);

NAND3xp33_ASAP7_75t_SL g441 ( 
.A(n_359),
.B(n_318),
.C(n_251),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_365),
.B(n_234),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_398),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_401),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_422),
.Y(n_445)
);

AND2x6_ASAP7_75t_SL g446 ( 
.A(n_379),
.B(n_15),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_365),
.B(n_237),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_412),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_383),
.B(n_238),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_L g450 ( 
.A(n_382),
.B(n_240),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_367),
.B(n_243),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_371),
.B(n_244),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_404),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_418),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_410),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_385),
.B(n_245),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_366),
.B(n_249),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_356),
.Y(n_458)
);

NOR2x1_ASAP7_75t_L g459 ( 
.A(n_406),
.B(n_256),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_R g460 ( 
.A(n_405),
.B(n_250),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_392),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_358),
.B(n_259),
.Y(n_462)
);

INVx5_ASAP7_75t_L g463 ( 
.A(n_411),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_369),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_408),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_370),
.B(n_381),
.Y(n_466)
);

NOR2x1p5_ASAP7_75t_L g467 ( 
.A(n_391),
.B(n_15),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_386),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_388),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_373),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_372),
.A2(n_298),
.B(n_283),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_415),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_376),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_L g474 ( 
.A(n_389),
.B(n_17),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_387),
.B(n_259),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_377),
.B(n_259),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_376),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_419),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_363),
.B(n_259),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_417),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_387),
.B(n_260),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_403),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_420),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_364),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_396),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_396),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_399),
.Y(n_487)
);

INVx5_ASAP7_75t_L g488 ( 
.A(n_400),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_395),
.B(n_260),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_399),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_394),
.A2(n_298),
.B1(n_283),
.B2(n_278),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_402),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_402),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_430),
.A2(n_413),
.B1(n_409),
.B2(n_421),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_425),
.B(n_423),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_442),
.A2(n_407),
.B1(n_416),
.B2(n_414),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_432),
.B(n_414),
.Y(n_497)
);

O2A1O1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_442),
.A2(n_416),
.B(n_16),
.C(n_417),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_424),
.B(n_260),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_451),
.B(n_417),
.Y(n_500)
);

O2A1O1Ixp33_ASAP7_75t_L g501 ( 
.A1(n_447),
.A2(n_417),
.B(n_298),
.C(n_283),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_440),
.A2(n_417),
.B(n_278),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_458),
.B(n_447),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_464),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_440),
.A2(n_278),
.B1(n_20),
.B2(n_22),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_R g506 ( 
.A(n_429),
.B(n_19),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_R g507 ( 
.A(n_433),
.B(n_24),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_445),
.B(n_27),
.Y(n_508)
);

NAND3xp33_ASAP7_75t_L g509 ( 
.A(n_456),
.B(n_450),
.C(n_457),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_482),
.B(n_29),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_471),
.A2(n_30),
.B(n_31),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_427),
.Y(n_512)
);

BUFx8_ASAP7_75t_SL g513 ( 
.A(n_457),
.Y(n_513)
);

O2A1O1Ixp33_ASAP7_75t_L g514 ( 
.A1(n_466),
.A2(n_32),
.B(n_33),
.C(n_35),
.Y(n_514)
);

INVx3_ASAP7_75t_SL g515 ( 
.A(n_470),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_433),
.Y(n_516)
);

INVx5_ASAP7_75t_L g517 ( 
.A(n_438),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_473),
.A2(n_36),
.B(n_38),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_431),
.Y(n_519)
);

O2A1O1Ixp33_ASAP7_75t_L g520 ( 
.A1(n_466),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_468),
.B(n_46),
.Y(n_521)
);

O2A1O1Ixp33_ASAP7_75t_L g522 ( 
.A1(n_436),
.A2(n_48),
.B(n_50),
.C(n_51),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_477),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_460),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_471),
.A2(n_59),
.B(n_61),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_438),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_469),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_461),
.B(n_65),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g529 ( 
.A(n_484),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_426),
.B(n_68),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_485),
.A2(n_69),
.B(n_70),
.Y(n_531)
);

A2O1A1Ixp33_ASAP7_75t_L g532 ( 
.A1(n_487),
.A2(n_75),
.B(n_77),
.C(n_78),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_490),
.A2(n_79),
.B(n_80),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_465),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_428),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_434),
.Y(n_536)
);

NOR3xp33_ASAP7_75t_SL g537 ( 
.A(n_441),
.B(n_449),
.C(n_479),
.Y(n_537)
);

NAND2x1p5_ASAP7_75t_L g538 ( 
.A(n_427),
.B(n_81),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_467),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_439),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_441),
.B(n_82),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_492),
.A2(n_83),
.B(n_84),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_443),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_493),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_480),
.A2(n_88),
.B(n_90),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_452),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_435),
.B(n_95),
.Y(n_547)
);

AND2x2_ASAP7_75t_SL g548 ( 
.A(n_475),
.B(n_96),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_437),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_475),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_486),
.B(n_98),
.Y(n_551)
);

A2O1A1Ixp33_ASAP7_75t_L g552 ( 
.A1(n_483),
.A2(n_99),
.B(n_100),
.C(n_102),
.Y(n_552)
);

OR2x6_ASAP7_75t_L g553 ( 
.A(n_481),
.B(n_103),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_549),
.B(n_427),
.Y(n_554)
);

BUFx12f_ASAP7_75t_L g555 ( 
.A(n_524),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_529),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_504),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_534),
.Y(n_558)
);

AO21x2_ASAP7_75t_L g559 ( 
.A1(n_502),
.A2(n_481),
.B(n_474),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_543),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_535),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_541),
.B(n_476),
.C(n_489),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_526),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_497),
.B(n_427),
.Y(n_564)
);

NAND2x1_ASAP7_75t_L g565 ( 
.A(n_512),
.B(n_448),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_550),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_519),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_516),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_503),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_536),
.Y(n_570)
);

OAI21x1_ASAP7_75t_L g571 ( 
.A1(n_501),
.A2(n_462),
.B(n_454),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_517),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_517),
.Y(n_573)
);

OR2x6_ASAP7_75t_L g574 ( 
.A(n_495),
.B(n_459),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_548),
.A2(n_472),
.B1(n_453),
.B2(n_444),
.Y(n_575)
);

BUFx2_ASAP7_75t_R g576 ( 
.A(n_513),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_517),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_499),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_515),
.Y(n_579)
);

BUFx2_ASAP7_75t_SL g580 ( 
.A(n_540),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_510),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_506),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_521),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_497),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_526),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_547),
.Y(n_586)
);

BUFx12f_ASAP7_75t_L g587 ( 
.A(n_526),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_530),
.A2(n_462),
.B(n_454),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_537),
.B(n_448),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g590 ( 
.A1(n_551),
.A2(n_511),
.B(n_545),
.Y(n_590)
);

BUFx12f_ASAP7_75t_L g591 ( 
.A(n_553),
.Y(n_591)
);

CKINVDCx11_ASAP7_75t_R g592 ( 
.A(n_553),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_498),
.A2(n_480),
.B(n_478),
.Y(n_593)
);

BUFx5_ASAP7_75t_L g594 ( 
.A(n_538),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_528),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_539),
.Y(n_596)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_531),
.A2(n_455),
.B(n_491),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_507),
.Y(n_598)
);

AOI22x1_ASAP7_75t_L g599 ( 
.A1(n_518),
.A2(n_438),
.B1(n_463),
.B2(n_488),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_508),
.A2(n_488),
.B1(n_463),
.B2(n_446),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_494),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_500),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_L g603 ( 
.A1(n_509),
.A2(n_488),
.B(n_463),
.Y(n_603)
);

OA21x2_ASAP7_75t_L g604 ( 
.A1(n_533),
.A2(n_542),
.B(n_505),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_546),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_523),
.A2(n_488),
.B1(n_463),
.B2(n_106),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_569),
.B(n_544),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_SL g608 ( 
.A1(n_591),
.A2(n_527),
.B1(n_496),
.B2(n_525),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_592),
.A2(n_522),
.B1(n_532),
.B2(n_520),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_L g610 ( 
.A1(n_601),
.A2(n_514),
.B(n_552),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_557),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_556),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_569),
.B(n_104),
.Y(n_613)
);

OAI21x1_ASAP7_75t_L g614 ( 
.A1(n_588),
.A2(n_590),
.B(n_571),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_560),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_560),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_582),
.Y(n_617)
);

AOI21x1_ASAP7_75t_L g618 ( 
.A1(n_602),
.A2(n_105),
.B(n_110),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_558),
.Y(n_619)
);

AO21x2_ASAP7_75t_L g620 ( 
.A1(n_559),
.A2(n_113),
.B(n_114),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_566),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_561),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_566),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_603),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_597),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_584),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_605),
.A2(n_119),
.B1(n_121),
.B2(n_123),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_567),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_592),
.A2(n_124),
.B1(n_126),
.B2(n_128),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_587),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_559),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_570),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_578),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_605),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_583),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_587),
.Y(n_636)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_593),
.A2(n_133),
.B(n_134),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_574),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_574),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_591),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_640)
);

BUFx2_ASAP7_75t_R g641 ( 
.A(n_580),
.Y(n_641)
);

INVx6_ASAP7_75t_L g642 ( 
.A(n_577),
.Y(n_642)
);

AO21x2_ASAP7_75t_L g643 ( 
.A1(n_593),
.A2(n_141),
.B(n_142),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_583),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_581),
.A2(n_143),
.B1(n_147),
.B2(n_148),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_L g646 ( 
.A1(n_600),
.A2(n_149),
.B1(n_150),
.B2(n_152),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_568),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_602),
.B(n_154),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_574),
.Y(n_649)
);

BUFx2_ASAP7_75t_SL g650 ( 
.A(n_577),
.Y(n_650)
);

AOI21x1_ASAP7_75t_L g651 ( 
.A1(n_604),
.A2(n_157),
.B(n_158),
.Y(n_651)
);

AOI21x1_ASAP7_75t_L g652 ( 
.A1(n_604),
.A2(n_159),
.B(n_160),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_603),
.Y(n_653)
);

INVxp67_ASAP7_75t_SL g654 ( 
.A(n_648),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_R g655 ( 
.A(n_630),
.B(n_555),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_623),
.B(n_585),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_612),
.B(n_589),
.Y(n_657)
);

NOR3xp33_ASAP7_75t_SL g658 ( 
.A(n_610),
.B(n_576),
.C(n_562),
.Y(n_658)
);

NOR3xp33_ASAP7_75t_SL g659 ( 
.A(n_646),
.B(n_576),
.C(n_555),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_628),
.B(n_596),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_609),
.A2(n_606),
.B1(n_575),
.B2(n_589),
.Y(n_661)
);

AND2x4_ASAP7_75t_SL g662 ( 
.A(n_636),
.B(n_554),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_623),
.Y(n_663)
);

NOR3xp33_ASAP7_75t_SL g664 ( 
.A(n_641),
.B(n_586),
.C(n_579),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_611),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_R g666 ( 
.A(n_630),
.B(n_598),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_R g667 ( 
.A(n_630),
.B(n_572),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_R g668 ( 
.A(n_648),
.B(n_624),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_622),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_617),
.Y(n_670)
);

NOR2x1p5_ASAP7_75t_L g671 ( 
.A(n_636),
.B(n_572),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_638),
.B(n_573),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_635),
.A2(n_595),
.B1(n_575),
.B2(n_606),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_636),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_622),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_619),
.Y(n_676)
);

AOI222xp33_ASAP7_75t_L g677 ( 
.A1(n_633),
.A2(n_596),
.B1(n_554),
.B2(n_564),
.C1(n_573),
.C2(n_595),
.Y(n_677)
);

OR2x6_ASAP7_75t_L g678 ( 
.A(n_639),
.B(n_649),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_632),
.B(n_564),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_R g680 ( 
.A(n_617),
.B(n_585),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_647),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_615),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_621),
.B(n_563),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_615),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_635),
.A2(n_594),
.B1(n_599),
.B2(n_604),
.Y(n_685)
);

CKINVDCx16_ASAP7_75t_R g686 ( 
.A(n_617),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_616),
.B(n_626),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_R g688 ( 
.A(n_624),
.B(n_563),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_626),
.B(n_565),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_613),
.B(n_594),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_SL g691 ( 
.A1(n_608),
.A2(n_629),
.B1(n_640),
.B2(n_653),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_644),
.B(n_594),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_SL g693 ( 
.A(n_607),
.B(n_594),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_642),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_613),
.B(n_594),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_644),
.B(n_594),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_642),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_650),
.B(n_161),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_607),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_616),
.Y(n_700)
);

AOI211xp5_ASAP7_75t_L g701 ( 
.A1(n_627),
.A2(n_634),
.B(n_637),
.C(n_653),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_618),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_618),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_650),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_704)
);

INVx2_ASAP7_75t_R g705 ( 
.A(n_643),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_657),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_666),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_667),
.Y(n_708)
);

OA21x2_ASAP7_75t_L g709 ( 
.A1(n_702),
.A2(n_614),
.B(n_631),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_699),
.B(n_665),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_676),
.B(n_643),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_663),
.B(n_643),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_654),
.B(n_669),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_675),
.B(n_625),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_684),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_687),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_682),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_700),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_678),
.B(n_631),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_656),
.B(n_625),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_703),
.Y(n_721)
);

INVx5_ASAP7_75t_L g722 ( 
.A(n_678),
.Y(n_722)
);

BUFx2_ASAP7_75t_SL g723 ( 
.A(n_671),
.Y(n_723)
);

INVxp67_ASAP7_75t_SL g724 ( 
.A(n_668),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_660),
.B(n_620),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_693),
.B(n_620),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_678),
.Y(n_727)
);

OR2x6_ASAP7_75t_SL g728 ( 
.A(n_661),
.B(n_620),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_693),
.B(n_637),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_658),
.A2(n_645),
.B(n_651),
.C(n_652),
.Y(n_730)
);

NAND2x1_ASAP7_75t_L g731 ( 
.A(n_694),
.B(n_642),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_690),
.B(n_614),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_692),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_686),
.B(n_642),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_695),
.B(n_652),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_680),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_679),
.B(n_651),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_689),
.B(n_166),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_705),
.B(n_168),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_681),
.B(n_169),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_694),
.B(n_172),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_SL g742 ( 
.A1(n_704),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_688),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_697),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_683),
.B(n_176),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_696),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_L g747 ( 
.A(n_701),
.B(n_659),
.C(n_704),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_672),
.B(n_177),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_697),
.B(n_179),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_747),
.B(n_701),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_710),
.B(n_674),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_736),
.B(n_691),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_713),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_732),
.B(n_685),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_744),
.B(n_708),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_713),
.B(n_724),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_722),
.B(n_672),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_707),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_723),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_744),
.B(n_691),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_715),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_715),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_725),
.B(n_697),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_746),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_716),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_706),
.B(n_670),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_717),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_721),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_718),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_721),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_733),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_743),
.B(n_673),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_725),
.B(n_664),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_733),
.B(n_677),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_732),
.B(n_655),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_722),
.B(n_698),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_714),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_744),
.B(n_677),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_714),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_720),
.B(n_662),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_711),
.B(n_183),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_711),
.B(n_745),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_753),
.B(n_712),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_771),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_775),
.B(n_737),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_771),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_764),
.B(n_712),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_751),
.B(n_737),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_782),
.B(n_735),
.Y(n_789)
);

NAND2x1p5_ASAP7_75t_L g790 ( 
.A(n_776),
.B(n_722),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_767),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_753),
.B(n_754),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_761),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_759),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_762),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_763),
.B(n_735),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_750),
.A2(n_728),
.B1(n_742),
.B2(n_730),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_776),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_756),
.B(n_727),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_777),
.B(n_719),
.Y(n_800)
);

NOR2xp67_ASAP7_75t_R g801 ( 
.A(n_750),
.B(n_722),
.Y(n_801)
);

NOR3xp33_ASAP7_75t_L g802 ( 
.A(n_797),
.B(n_752),
.C(n_766),
.Y(n_802)
);

OR2x2_ASAP7_75t_L g803 ( 
.A(n_792),
.B(n_779),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_784),
.Y(n_804)
);

INVxp67_ASAP7_75t_SL g805 ( 
.A(n_787),
.Y(n_805)
);

AOI32xp33_ASAP7_75t_L g806 ( 
.A1(n_797),
.A2(n_752),
.A3(n_760),
.B1(n_773),
.B2(n_754),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_785),
.B(n_755),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_796),
.B(n_755),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_798),
.B(n_759),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_792),
.B(n_765),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_786),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_809),
.Y(n_812)
);

NAND3xp33_ASAP7_75t_L g813 ( 
.A(n_806),
.B(n_760),
.C(n_791),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_802),
.Y(n_814)
);

XOR2x2_ASAP7_75t_L g815 ( 
.A(n_806),
.B(n_794),
.Y(n_815)
);

AOI21xp33_ASAP7_75t_L g816 ( 
.A1(n_805),
.A2(n_772),
.B(n_778),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_810),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_803),
.B(n_787),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_814),
.A2(n_774),
.B1(n_726),
.B2(n_776),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_817),
.Y(n_820)
);

OAI221xp5_ASAP7_75t_L g821 ( 
.A1(n_813),
.A2(n_730),
.B1(n_799),
.B2(n_789),
.C(n_795),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_818),
.B(n_807),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_815),
.A2(n_801),
.B(n_758),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_812),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_824),
.B(n_758),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_820),
.B(n_816),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_823),
.B(n_822),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_821),
.B(n_808),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_826),
.B(n_819),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_825),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_828),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_831),
.A2(n_827),
.B(n_740),
.C(n_781),
.Y(n_832)
);

OAI221xp5_ASAP7_75t_L g833 ( 
.A1(n_829),
.A2(n_830),
.B1(n_769),
.B2(n_726),
.C(n_804),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_829),
.A2(n_738),
.B1(n_745),
.B2(n_811),
.Y(n_834)
);

AOI22x1_ASAP7_75t_SL g835 ( 
.A1(n_832),
.A2(n_798),
.B1(n_801),
.B2(n_734),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_834),
.Y(n_836)
);

NOR2x1_ASAP7_75t_L g837 ( 
.A(n_833),
.B(n_748),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_834),
.B(n_788),
.Y(n_838)
);

AND2x2_ASAP7_75t_SL g839 ( 
.A(n_834),
.B(n_749),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_836),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_837),
.A2(n_749),
.B(n_741),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_839),
.A2(n_738),
.B1(n_729),
.B2(n_793),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_838),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_838),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_835),
.B(n_783),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_840),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_844),
.A2(n_731),
.B(n_741),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_843),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_845),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_841),
.Y(n_850)
);

INVx1_ASAP7_75t_SL g851 ( 
.A(n_846),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_848),
.Y(n_852)
);

XOR2xp5_ASAP7_75t_L g853 ( 
.A(n_849),
.B(n_842),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_850),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_852),
.B(n_849),
.Y(n_855)
);

AOI31xp33_ASAP7_75t_L g856 ( 
.A1(n_851),
.A2(n_847),
.A3(n_790),
.B(n_739),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_854),
.A2(n_728),
.B1(n_790),
.B2(n_800),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_853),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_858),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_859),
.A2(n_855),
.B1(n_857),
.B2(n_856),
.Y(n_860)
);

XNOR2xp5_ASAP7_75t_L g861 ( 
.A(n_860),
.B(n_739),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_861),
.A2(n_770),
.B1(n_768),
.B2(n_729),
.Y(n_862)
);

AOI221xp5_ASAP7_75t_L g863 ( 
.A1(n_862),
.A2(n_768),
.B1(n_770),
.B2(n_780),
.C(n_719),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_863),
.A2(n_709),
.B1(n_757),
.B2(n_719),
.Y(n_864)
);


endmodule