module fake_aes_6586_n_28 (n_1, n_2, n_4, n_3, n_0, n_28);
input n_1;
input n_2;
input n_4;
input n_3;
input n_0;
output n_28;
wire n_20;
wire n_5;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_6;
wire n_7;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g5 ( .A(n_1), .Y(n_5) );
INVxp67_ASAP7_75t_L g6 ( .A(n_2), .Y(n_6) );
BUFx10_ASAP7_75t_L g7 ( .A(n_0), .Y(n_7) );
NAND2xp5_ASAP7_75t_SL g8 ( .A(n_0), .B(n_4), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_4), .Y(n_9) );
AND2x2_ASAP7_75t_L g10 ( .A(n_7), .B(n_0), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_7), .B(n_0), .Y(n_11) );
OAI22xp5_ASAP7_75t_L g12 ( .A1(n_5), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_12) );
AOI221xp5_ASAP7_75t_L g13 ( .A1(n_6), .A2(n_1), .B1(n_2), .B2(n_3), .C(n_4), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_7), .B(n_3), .Y(n_14) );
BUFx3_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
INVx3_ASAP7_75t_L g16 ( .A(n_11), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_13), .B(n_7), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_15), .Y(n_21) );
AOI211x1_ASAP7_75t_SL g22 ( .A1(n_19), .A2(n_12), .B(n_8), .C(n_7), .Y(n_22) );
AOI221xp5_ASAP7_75t_SL g23 ( .A1(n_21), .A2(n_18), .B1(n_16), .B2(n_6), .C(n_12), .Y(n_23) );
NOR2xp33_ASAP7_75t_L g24 ( .A(n_23), .B(n_18), .Y(n_24) );
OAI211xp5_ASAP7_75t_L g25 ( .A1(n_22), .A2(n_17), .B(n_21), .C(n_20), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
AOI22xp5_ASAP7_75t_SL g27 ( .A1(n_24), .A2(n_17), .B1(n_9), .B2(n_22), .Y(n_27) );
OAI221xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_9), .B1(n_15), .B2(n_16), .C(n_26), .Y(n_28) );
endmodule