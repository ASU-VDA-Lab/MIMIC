module fake_jpeg_1616_n_102 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_35),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_41),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_28),
.C(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_46),
.Y(n_57)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_35),
.B(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_52),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_36),
.B1(n_38),
.B2(n_28),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_56),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_41),
.B(n_30),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_58),
.B(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_27),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_32),
.B(n_27),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_57),
.B(n_48),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_60),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

AOI22x1_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_42),
.B1(n_12),
.B2(n_13),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_64),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_42),
.B(n_1),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_26),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_66),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_25),
.C(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_72),
.B(n_73),
.Y(n_79)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_76),
.B(n_0),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_53),
.B1(n_22),
.B2(n_20),
.Y(n_78)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_19),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_77),
.C(n_75),
.Y(n_80)
);

A2O1A1O1Ixp25_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_14),
.B(n_11),
.C(n_7),
.D(n_8),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_53),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_82),
.B(n_84),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_71),
.C(n_78),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_87),
.B1(n_17),
.B2(n_15),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_2),
.B(n_3),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_90),
.Y(n_94)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_87),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_80),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_95),
.Y(n_96)
);

OAI21x1_ASAP7_75t_SL g97 ( 
.A1(n_96),
.A2(n_94),
.B(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_92),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_5),
.B(n_6),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_7),
.B(n_9),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);


endmodule