module fake_jpeg_426_n_208 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_208);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_20),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_7),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_33),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_77),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_0),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_68),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

BUFx8_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_81),
.A2(n_60),
.B1(n_63),
.B2(n_54),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_92),
.B1(n_73),
.B2(n_72),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_67),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_59),
.B1(n_66),
.B2(n_74),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_50),
.B1(n_54),
.B2(n_65),
.Y(n_110)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_52),
.B1(n_59),
.B2(n_66),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_52),
.B1(n_51),
.B2(n_57),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_72),
.B1(n_56),
.B2(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_70),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_100),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_19),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_64),
.B(n_58),
.C(n_63),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_106),
.Y(n_119)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_110),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_53),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_63),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_53),
.Y(n_109)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_21),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_1),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_104),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_116),
.B(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

XNOR2x1_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_83),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_122),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_65),
.C(n_50),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_132),
.Y(n_139)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_1),
.Y(n_130)
);

AND2x4_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_49),
.Y(n_131)
);

FAx1_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_2),
.CI(n_5),
.CON(n_137),
.SN(n_137)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_107),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_127),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_140),
.B1(n_146),
.B2(n_156),
.Y(n_174)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_138),
.C(n_143),
.Y(n_164)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_25),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_127),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_145),
.Y(n_171)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_26),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_123),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_29),
.B1(n_47),
.B2(n_46),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_9),
.B(n_10),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_152),
.B(n_16),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_SL g149 ( 
.A(n_130),
.B(n_11),
.C(n_12),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_31),
.C(n_36),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_14),
.B(n_15),
.Y(n_152)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_117),
.A2(n_32),
.B1(n_45),
.B2(n_38),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_154),
.A2(n_131),
.B(n_18),
.Y(n_163)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_120),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_166),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_131),
.Y(n_160)
);

XNOR2x1_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_169),
.Y(n_178)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_23),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_173),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_28),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_172),
.Y(n_183)
);

NOR2x1_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_37),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_137),
.B1(n_143),
.B2(n_138),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_172),
.A2(n_137),
.B(n_154),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_180),
.B(n_160),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_153),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_168),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_189),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_188),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_161),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_157),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_190),
.B(n_191),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_178),
.B(n_158),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_192),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_186),
.A2(n_181),
.B(n_164),
.Y(n_194)
);

OAI31xp33_ASAP7_75t_L g199 ( 
.A1(n_194),
.A2(n_181),
.A3(n_177),
.B(n_168),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_199),
.B(n_200),
.Y(n_202)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_196),
.A2(n_185),
.B1(n_174),
.B2(n_182),
.Y(n_201)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_201),
.B(n_185),
.CI(n_195),
.CON(n_203),
.SN(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_195),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_204),
.A2(n_202),
.B(n_197),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_164),
.B(n_193),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_203),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_183),
.Y(n_208)
);


endmodule