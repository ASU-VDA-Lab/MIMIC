module real_jpeg_14890_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_381, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_381;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_3),
.B(n_42),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_3),
.B(n_36),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_3),
.B(n_31),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_3),
.B(n_89),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_3),
.B(n_56),
.Y(n_319)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_5),
.B(n_45),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_5),
.B(n_31),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_5),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_5),
.B(n_70),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_5),
.B(n_89),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_5),
.B(n_42),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_6),
.B(n_25),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_6),
.B(n_89),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_6),
.B(n_36),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_6),
.B(n_31),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_6),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_6),
.B(n_56),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_6),
.B(n_42),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_6),
.B(n_45),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_7),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_7),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_7),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_7),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_7),
.B(n_25),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_7),
.B(n_89),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_7),
.B(n_56),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_10),
.B(n_89),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_10),
.B(n_56),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_10),
.B(n_25),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_10),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_10),
.B(n_42),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_12),
.B(n_42),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_12),
.B(n_25),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_12),
.B(n_89),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_12),
.B(n_70),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_12),
.B(n_36),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_13),
.B(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_13),
.B(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_13),
.B(n_31),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_13),
.B(n_36),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_14),
.B(n_42),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_14),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_14),
.B(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_14),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_14),
.B(n_36),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_14),
.B(n_70),
.Y(n_211)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_148),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_147),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_20),
.B(n_123),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_20),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_20),
.B(n_150),
.Y(n_377)
);

FAx1_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_63),
.CI(n_97),
.CON(n_20),
.SN(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_40),
.C(n_49),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_22),
.A2(n_23),
.B1(n_40),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_24),
.B(n_30),
.C(n_34),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_24),
.A2(n_39),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_24),
.B(n_141),
.C(n_313),
.Y(n_341)
);

INVx5_ASAP7_75t_SL g199 ( 
.A(n_25),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_29),
.A2(n_30),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_29),
.A2(n_30),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_30),
.B(n_88),
.C(n_92),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_30),
.B(n_251),
.C(n_253),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_32),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_32),
.B(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_32),
.B(n_58),
.Y(n_317)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_67),
.C(n_75),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_34),
.A2(n_35),
.B1(n_75),
.B2(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_34),
.A2(n_35),
.B1(n_122),
.B2(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_34),
.A2(n_35),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_35),
.B(n_119),
.C(n_122),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_35),
.B(n_211),
.Y(n_265)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_37),
.B(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_37),
.B(n_230),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_40),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_43),
.C(n_48),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_41),
.A2(n_43),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_42),
.Y(n_132)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_73),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_44),
.B(n_58),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_44),
.B(n_230),
.Y(n_301)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_47),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_47),
.B(n_199),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_49),
.A2(n_50),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_62),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_54),
.C(n_59),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_55),
.B(n_187),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_61),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_61),
.B(n_189),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_85),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_77),
.B2(n_78),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_65),
.B(n_78),
.C(n_85),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_67),
.A2(n_68),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.C(n_74),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_69),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_69),
.B(n_120),
.C(n_121),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_69),
.A2(n_112),
.B1(n_120),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_69),
.A2(n_112),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_69),
.B(n_191),
.Y(n_207)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_70),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_71),
.A2(n_72),
.B1(n_92),
.B2(n_93),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_71),
.B(n_92),
.C(n_301),
.Y(n_320)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_74),
.A2(n_110),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_84),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_80),
.B(n_82),
.C(n_83),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_81),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_94),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_95),
.C(n_96),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_87),
.A2(n_88),
.B1(n_106),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_106),
.C(n_107),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_92),
.A2(n_93),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_114),
.C(n_118),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_98),
.A2(n_99),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_105),
.C(n_108),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_100),
.A2(n_101),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_105),
.A2(n_108),
.B1(n_109),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_106),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_107),
.B(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_114),
.B(n_118),
.Y(n_172)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_120),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_120),
.A2(n_163),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_120),
.B(n_258),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_122),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_146),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_144),
.B2(n_145),
.Y(n_124)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_135),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_142),
.B2(n_143),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_140),
.A2(n_141),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_173),
.B(n_377),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_166),
.C(n_170),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_151),
.B(n_370),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_157),
.C(n_160),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_152),
.A2(n_153),
.B1(n_364),
.B2(n_365),
.Y(n_363)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_157),
.B(n_160),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_165),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_161),
.B(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_164),
.A2(n_165),
.B1(n_349),
.B2(n_350),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_164),
.Y(n_350)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_165),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_166),
.B(n_170),
.Y(n_370)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI321xp33_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_357),
.A3(n_367),
.B1(n_371),
.B2(n_376),
.C(n_381),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_304),
.C(n_352),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_275),
.B(n_303),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_245),
.B(n_274),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_214),
.B(n_244),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_193),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_179),
.B(n_193),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.C(n_190),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_196),
.B1(n_197),
.B2(n_205),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_180),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_180),
.B(n_241),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.CI(n_183),
.CON(n_180),
.SN(n_180)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_184),
.A2(n_185),
.B1(n_190),
.B2(n_242),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_186),
.B(n_188),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_189),
.B(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_190),
.Y(n_242)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_206),
.B2(n_213),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_196),
.B(n_205),
.C(n_213),
.Y(n_246)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_198),
.B(n_201),
.C(n_204),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_203),
.Y(n_204)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_207),
.B(n_209),
.C(n_210),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_211),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_211),
.A2(n_212),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_211),
.B(n_325),
.C(n_328),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_238),
.B(n_243),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_227),
.B(n_237),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_222),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_225),
.C(n_226),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_232),
.B(n_236),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_229),
.B(n_231),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_239),
.B(n_240),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_246),
.B(n_247),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_260),
.B2(n_261),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_262),
.C(n_273),
.Y(n_276)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_255),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_256),
.C(n_257),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_272),
.B2(n_273),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_271),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_268),
.C(n_270),
.Y(n_294)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_266),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_267),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_276),
.B(n_277),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_293),
.B2(n_302),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_292),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_280),
.B(n_292),
.C(n_302),
.Y(n_353)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_288),
.B2(n_289),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_283),
.B(n_290),
.C(n_291),
.Y(n_321)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g379 ( 
.A(n_284),
.Y(n_379)
);

FAx1_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_286),
.CI(n_287),
.CON(n_284),
.SN(n_284)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_285),
.B(n_286),
.C(n_287),
.Y(n_330)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_293),
.Y(n_302)
);

BUFx24_ASAP7_75t_SL g380 ( 
.A(n_293),
.Y(n_380)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_295),
.CI(n_299),
.CON(n_293),
.SN(n_293)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_294),
.B(n_295),
.C(n_299),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B(n_298),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_297),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_298),
.A2(n_330),
.B1(n_331),
.B2(n_332),
.Y(n_329)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_298),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

AOI21xp33_ASAP7_75t_L g372 ( 
.A1(n_305),
.A2(n_373),
.B(n_374),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_334),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_306),
.B(n_334),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_322),
.C(n_333),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_307),
.B(n_355),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_321),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_314),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_309),
.B(n_314),
.C(n_321),
.Y(n_351)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_312),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_317),
.B(n_318),
.C(n_320),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_322),
.A2(n_323),
.B1(n_333),
.B2(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_329),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_330),
.C(n_332),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_327),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_330),
.Y(n_331)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_333),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_351),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_343),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_336),
.B(n_343),
.C(n_351),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_340),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_341),
.C(n_342),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_346),
.C(n_347),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_354),
.Y(n_373)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_358),
.A2(n_372),
.B(n_375),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_359),
.B(n_360),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_366),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_363),
.C(n_366),
.Y(n_368)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_368),
.B(n_369),
.Y(n_376)
);


endmodule