module fake_netlist_1_12466_n_40 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
wire n_39;
INVx3_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_2), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_4), .Y(n_18) );
CKINVDCx20_ASAP7_75t_R g19 ( .A(n_7), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_13), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_13), .B(n_0), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_13), .B(n_0), .Y(n_23) );
INVx1_ASAP7_75t_SL g24 ( .A(n_22), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_21), .Y(n_25) );
AOI22xp5_ASAP7_75t_L g26 ( .A1(n_20), .A2(n_19), .B1(n_18), .B2(n_17), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
OAI211xp5_ASAP7_75t_SL g29 ( .A1(n_28), .A2(n_26), .B(n_24), .C(n_23), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
NOR4xp25_ASAP7_75t_SL g32 ( .A(n_29), .B(n_15), .C(n_19), .D(n_27), .Y(n_32) );
AOI22xp5_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_14), .B1(n_2), .B2(n_3), .Y(n_33) );
OAI22xp5_ASAP7_75t_L g34 ( .A1(n_31), .A2(n_1), .B1(n_4), .B2(n_5), .Y(n_34) );
INVx2_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
OR5x1_ASAP7_75t_L g36 ( .A(n_34), .B(n_32), .C(n_6), .D(n_9), .E(n_10), .Y(n_36) );
INVx2_ASAP7_75t_L g37 ( .A(n_36), .Y(n_37) );
INVxp67_ASAP7_75t_L g38 ( .A(n_35), .Y(n_38) );
NAND2xp5_ASAP7_75t_L g39 ( .A(n_38), .B(n_37), .Y(n_39) );
HB1xp67_ASAP7_75t_L g40 ( .A(n_39), .Y(n_40) );
endmodule