module fake_netlist_6_842_n_1229 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_18, n_21, n_193, n_147, n_269, n_258, n_281, n_154, n_191, n_88, n_3, n_209, n_98, n_277, n_260, n_265, n_283, n_113, n_39, n_63, n_223, n_278, n_270, n_73, n_279, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_166, n_28, n_184, n_212, n_268, n_271, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_285, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_286, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_284, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_274, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_289, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_267, n_282, n_58, n_116, n_280, n_211, n_287, n_64, n_220, n_288, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_273, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_272, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_275, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_276, n_51, n_44, n_56, n_221, n_1229);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_18;
input n_21;
input n_193;
input n_147;
input n_269;
input n_258;
input n_281;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_277;
input n_260;
input n_265;
input n_283;
input n_113;
input n_39;
input n_63;
input n_223;
input n_278;
input n_270;
input n_73;
input n_279;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_166;
input n_28;
input n_184;
input n_212;
input n_268;
input n_271;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_285;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_286;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_284;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_274;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_289;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_267;
input n_282;
input n_58;
input n_116;
input n_280;
input n_211;
input n_287;
input n_64;
input n_220;
input n_288;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_273;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_272;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_275;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_276;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1229;

wire n_992;
wire n_801;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1032;
wire n_893;
wire n_1099;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_836;
wire n_375;
wire n_522;
wire n_945;
wire n_1143;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_487;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_530;
wire n_618;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_304;
wire n_694;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_615;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_899;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_292;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1223;
wire n_303;
wire n_511;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_848;
wire n_301;
wire n_1096;
wire n_1091;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_575;
wire n_368;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_1213;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_548;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_652;
wire n_560;
wire n_569;
wire n_737;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_502;
wire n_672;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_300;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_709;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_670;
wire n_1089;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_649;

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_121),
.Y(n_290)
);

HB1xp67_ASAP7_75t_SL g291 ( 
.A(n_30),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_206),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_110),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_131),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_237),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_112),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_0),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_244),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_178),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_182),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_183),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_31),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_282),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_30),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_239),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_119),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_111),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_145),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_196),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_261),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_66),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_10),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_151),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_33),
.Y(n_314)
);

BUFx8_ASAP7_75t_SL g315 ( 
.A(n_138),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_276),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_86),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_67),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_232),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_235),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_181),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_264),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_163),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_249),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_42),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_134),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_16),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_190),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_91),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_100),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_127),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_22),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_142),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_17),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_13),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_95),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_286),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_5),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_260),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_220),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_162),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_184),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_80),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_126),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_169),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_284),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_16),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_204),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_152),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_34),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_255),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_192),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_154),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_189),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_202),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_267),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_24),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_146),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_29),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_247),
.Y(n_360)
);

BUFx8_ASAP7_75t_SL g361 ( 
.A(n_12),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_188),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_106),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_156),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_281),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_274),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_0),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_96),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_140),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_48),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_83),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_268),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_263),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_139),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_31),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_113),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_116),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_222),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_109),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_90),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_92),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_97),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_283),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_19),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_217),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_229),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_285),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_62),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_42),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_270),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_123),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_57),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_287),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_259),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_107),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_170),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_225),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_280),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_230),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_137),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_289),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_233),
.Y(n_402)
);

BUFx10_ASAP7_75t_L g403 ( 
.A(n_279),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_52),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_174),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_41),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_54),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_231),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_155),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_173),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_10),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_47),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_108),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_200),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_214),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_240),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_216),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_165),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_32),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_17),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_28),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_115),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_47),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_221),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_185),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_128),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_177),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_180),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_161),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_124),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_215),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_213),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_179),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_11),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_212),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_87),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_99),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_80),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_83),
.Y(n_439)
);

BUFx10_ASAP7_75t_L g440 ( 
.A(n_198),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_144),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_193),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_25),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_136),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_53),
.Y(n_445)
);

BUFx8_ASAP7_75t_SL g446 ( 
.A(n_194),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_234),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_245),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_262),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_236),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_39),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_20),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_159),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_223),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_241),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_187),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_130),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_266),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_71),
.Y(n_459)
);

BUFx2_ASAP7_75t_R g460 ( 
.A(n_186),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_34),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_224),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_56),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_271),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_238),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_7),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_41),
.Y(n_467)
);

BUFx5_ASAP7_75t_L g468 ( 
.A(n_22),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_251),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_175),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_105),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_278),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_46),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_207),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_21),
.Y(n_475)
);

BUFx5_ASAP7_75t_L g476 ( 
.A(n_39),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_143),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_208),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_375),
.B(n_1),
.Y(n_479)
);

INVx5_ASAP7_75t_L g480 ( 
.A(n_306),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_344),
.B(n_2),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_468),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_336),
.B(n_2),
.Y(n_483)
);

AND2x6_ASAP7_75t_L g484 ( 
.A(n_432),
.B(n_93),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_468),
.B(n_3),
.Y(n_485)
);

BUFx8_ASAP7_75t_L g486 ( 
.A(n_413),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_306),
.Y(n_487)
);

INVx5_ASAP7_75t_L g488 ( 
.A(n_306),
.Y(n_488)
);

INVx5_ASAP7_75t_L g489 ( 
.A(n_306),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_468),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_309),
.Y(n_491)
);

INVx6_ASAP7_75t_L g492 ( 
.A(n_326),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_327),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_309),
.Y(n_494)
);

INVx5_ASAP7_75t_L g495 ( 
.A(n_309),
.Y(n_495)
);

BUFx8_ASAP7_75t_SL g496 ( 
.A(n_361),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_309),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_417),
.Y(n_498)
);

BUFx12f_ASAP7_75t_L g499 ( 
.A(n_326),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_417),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_344),
.B(n_3),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_336),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_410),
.B(n_4),
.Y(n_503)
);

INVx6_ASAP7_75t_L g504 ( 
.A(n_326),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_468),
.B(n_4),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_476),
.Y(n_506)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_417),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_417),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_410),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_476),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_361),
.B(n_6),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_319),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_432),
.B(n_6),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_319),
.B(n_7),
.Y(n_514)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_396),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_318),
.B(n_8),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_348),
.B(n_8),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_476),
.B(n_9),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_459),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_348),
.B(n_12),
.Y(n_520)
);

INVx5_ASAP7_75t_L g521 ( 
.A(n_396),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_387),
.B(n_13),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_313),
.B(n_14),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_365),
.B(n_14),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_302),
.Y(n_525)
);

BUFx8_ASAP7_75t_SL g526 ( 
.A(n_315),
.Y(n_526)
);

NOR2x1_ASAP7_75t_L g527 ( 
.A(n_387),
.B(n_15),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_396),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_314),
.B(n_18),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_405),
.B(n_20),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_405),
.B(n_21),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_401),
.B(n_23),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_304),
.Y(n_533)
);

INVx5_ASAP7_75t_L g534 ( 
.A(n_403),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_327),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_411),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_290),
.Y(n_537)
);

INVx6_ASAP7_75t_L g538 ( 
.A(n_403),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_420),
.B(n_24),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_411),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_430),
.B(n_25),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_403),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_440),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_430),
.B(n_26),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_297),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_299),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_311),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_312),
.Y(n_548)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_440),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_301),
.B(n_358),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_394),
.B(n_26),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_425),
.B(n_427),
.Y(n_552)
);

CKINVDCx11_ASAP7_75t_R g553 ( 
.A(n_407),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_360),
.B(n_27),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_300),
.Y(n_555)
);

BUFx8_ASAP7_75t_SL g556 ( 
.A(n_446),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_408),
.B(n_27),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_292),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_437),
.B(n_28),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_444),
.B(n_29),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_323),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_450),
.B(n_32),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_317),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_308),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_324),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_339),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_338),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_346),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_469),
.B(n_33),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_294),
.B(n_35),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_293),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_351),
.B(n_35),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_320),
.B(n_36),
.Y(n_573)
);

BUFx12f_ASAP7_75t_L g574 ( 
.A(n_325),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_322),
.B(n_37),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_295),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_391),
.B(n_38),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_352),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_353),
.Y(n_579)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_446),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_298),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_354),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_388),
.B(n_40),
.Y(n_583)
);

INVx5_ASAP7_75t_L g584 ( 
.A(n_291),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_395),
.B(n_40),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_404),
.B(n_43),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_372),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_332),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_373),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_423),
.B(n_44),
.Y(n_590)
);

INVx5_ASAP7_75t_L g591 ( 
.A(n_334),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_378),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_434),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_335),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_381),
.B(n_386),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_343),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_399),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_416),
.B(n_44),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_400),
.B(n_45),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_347),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_303),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_443),
.B(n_45),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_350),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_451),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_357),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_461),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_SL g607 ( 
.A(n_460),
.B(n_48),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_418),
.B(n_49),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_424),
.Y(n_609)
);

OAI22xp33_ASAP7_75t_SL g610 ( 
.A1(n_559),
.A2(n_367),
.B1(n_370),
.B2(n_359),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_481),
.B(n_428),
.Y(n_611)
);

NOR2x1p5_ASAP7_75t_L g612 ( 
.A(n_543),
.B(n_371),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_552),
.A2(n_560),
.B1(n_551),
.B2(n_501),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_543),
.B(n_453),
.Y(n_614)
);

NAND2x1p5_ASAP7_75t_L g615 ( 
.A(n_584),
.B(n_433),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_487),
.Y(n_616)
);

BUFx6f_ASAP7_75t_SL g617 ( 
.A(n_515),
.Y(n_617)
);

OAI22xp33_ASAP7_75t_R g618 ( 
.A1(n_570),
.A2(n_463),
.B1(n_467),
.B2(n_466),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_599),
.A2(n_462),
.B1(n_426),
.B2(n_333),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_545),
.B(n_305),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_515),
.B(n_435),
.Y(n_621)
);

AO22x2_ASAP7_75t_L g622 ( 
.A1(n_513),
.A2(n_441),
.B1(n_458),
.B2(n_455),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_487),
.Y(n_623)
);

AO22x2_ASAP7_75t_L g624 ( 
.A1(n_513),
.A2(n_465),
.B1(n_471),
.B2(n_464),
.Y(n_624)
);

OAI22xp33_ASAP7_75t_SL g625 ( 
.A1(n_511),
.A2(n_389),
.B1(n_392),
.B2(n_384),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_548),
.B(n_307),
.Y(n_626)
);

OAI22xp33_ASAP7_75t_L g627 ( 
.A1(n_607),
.A2(n_412),
.B1(n_421),
.B2(n_406),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_570),
.A2(n_340),
.B1(n_393),
.B2(n_296),
.Y(n_628)
);

OAI22xp33_ASAP7_75t_SL g629 ( 
.A1(n_492),
.A2(n_438),
.B1(n_439),
.B2(n_436),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_537),
.B(n_478),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_487),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_494),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_588),
.B(n_310),
.Y(n_633)
);

AO22x2_ASAP7_75t_L g634 ( 
.A1(n_483),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_573),
.A2(n_457),
.B1(n_442),
.B2(n_452),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_528),
.A2(n_445),
.B1(n_475),
.B2(n_473),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_494),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_494),
.Y(n_638)
);

AND2x2_ASAP7_75t_SL g639 ( 
.A(n_479),
.B(n_419),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_576),
.B(n_316),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_563),
.B(n_321),
.Y(n_641)
);

AO22x2_ASAP7_75t_L g642 ( 
.A1(n_483),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_642)
);

OR2x6_ASAP7_75t_L g643 ( 
.A(n_574),
.B(n_419),
.Y(n_643)
);

BUFx6f_ASAP7_75t_SL g644 ( 
.A(n_496),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_502),
.B(n_328),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_SL g646 ( 
.A1(n_492),
.A2(n_538),
.B1(n_504),
.B2(n_557),
.Y(n_646)
);

AO22x2_ASAP7_75t_L g647 ( 
.A1(n_503),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_575),
.A2(n_330),
.B1(n_331),
.B2(n_329),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_521),
.B(n_337),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_577),
.A2(n_342),
.B1(n_345),
.B2(n_341),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_498),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_498),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_585),
.A2(n_355),
.B1(n_356),
.B2(n_349),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_512),
.Y(n_654)
);

AO22x2_ASAP7_75t_L g655 ( 
.A1(n_503),
.A2(n_59),
.B1(n_55),
.B2(n_58),
.Y(n_655)
);

OAI22xp33_ASAP7_75t_SL g656 ( 
.A1(n_504),
.A2(n_363),
.B1(n_364),
.B2(n_362),
.Y(n_656)
);

OAI22xp33_ASAP7_75t_L g657 ( 
.A1(n_557),
.A2(n_368),
.B1(n_369),
.B2(n_366),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_498),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_526),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_500),
.Y(n_660)
);

AO22x2_ASAP7_75t_L g661 ( 
.A1(n_554),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_500),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_SL g663 ( 
.A1(n_538),
.A2(n_376),
.B1(n_377),
.B2(n_374),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_562),
.A2(n_380),
.B1(n_382),
.B2(n_379),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_581),
.B(n_383),
.Y(n_665)
);

OAI22xp33_ASAP7_75t_L g666 ( 
.A1(n_562),
.A2(n_477),
.B1(n_474),
.B2(n_472),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_521),
.B(n_385),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_601),
.B(n_390),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_500),
.Y(n_669)
);

AO22x2_ASAP7_75t_L g670 ( 
.A1(n_554),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_670)
);

AND2x2_ASAP7_75t_SL g671 ( 
.A(n_514),
.B(n_517),
.Y(n_671)
);

OAI22xp33_ASAP7_75t_L g672 ( 
.A1(n_520),
.A2(n_470),
.B1(n_456),
.B2(n_454),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_520),
.A2(n_541),
.B1(n_544),
.B2(n_530),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_SL g674 ( 
.A1(n_541),
.A2(n_449),
.B1(n_448),
.B2(n_447),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_508),
.Y(n_675)
);

AO22x2_ASAP7_75t_L g676 ( 
.A1(n_514),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_676)
);

OR2x6_ASAP7_75t_L g677 ( 
.A(n_499),
.B(n_65),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_512),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_508),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_544),
.A2(n_431),
.B1(n_429),
.B2(n_422),
.Y(n_680)
);

AO22x2_ASAP7_75t_L g681 ( 
.A1(n_517),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_681)
);

AO22x2_ASAP7_75t_L g682 ( 
.A1(n_522),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_508),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_534),
.B(n_397),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_523),
.A2(n_409),
.B1(n_415),
.B2(n_414),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_542),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_509),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_550),
.B(n_398),
.Y(n_688)
);

AO22x2_ASAP7_75t_L g689 ( 
.A1(n_522),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_553),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_482),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_523),
.A2(n_402),
.B1(n_73),
.B2(n_74),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_542),
.B(n_94),
.Y(n_693)
);

AO22x2_ASAP7_75t_L g694 ( 
.A1(n_531),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_490),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_524),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_558),
.B(n_78),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_671),
.B(n_595),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_631),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_631),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_658),
.Y(n_701)
);

INVxp67_ASAP7_75t_SL g702 ( 
.A(n_623),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_614),
.B(n_571),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_691),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_658),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_654),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_673),
.B(n_571),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_617),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_678),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_613),
.B(n_595),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_619),
.B(n_519),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_623),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_651),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_663),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_628),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_616),
.Y(n_716)
);

INVxp67_ASAP7_75t_SL g717 ( 
.A(n_632),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_637),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_687),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_638),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_652),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_660),
.Y(n_722)
);

XOR2xp5_ASAP7_75t_L g723 ( 
.A(n_659),
.B(n_547),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_645),
.B(n_550),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_662),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_611),
.B(n_630),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_695),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_669),
.Y(n_728)
);

OAI21xp5_ASAP7_75t_L g729 ( 
.A1(n_668),
.A2(n_484),
.B(n_485),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_675),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_640),
.A2(n_488),
.B(n_480),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_679),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_683),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_622),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_693),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_672),
.B(n_584),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_622),
.Y(n_737)
);

OAI21xp5_ASAP7_75t_L g738 ( 
.A1(n_641),
.A2(n_484),
.B(n_485),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_624),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_624),
.Y(n_740)
);

OAI21xp5_ASAP7_75t_L g741 ( 
.A1(n_620),
.A2(n_484),
.B(n_505),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_688),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_688),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_626),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_649),
.B(n_480),
.Y(n_745)
);

CKINVDCx20_ASAP7_75t_R g746 ( 
.A(n_635),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_633),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_665),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_612),
.Y(n_749)
);

XOR2xp5_ASAP7_75t_L g750 ( 
.A(n_659),
.B(n_639),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_621),
.B(n_529),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_686),
.B(n_539),
.Y(n_752)
);

INVxp33_ASAP7_75t_L g753 ( 
.A(n_636),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_667),
.B(n_584),
.Y(n_754)
);

AO21x1_ASAP7_75t_L g755 ( 
.A1(n_657),
.A2(n_532),
.B(n_524),
.Y(n_755)
);

XOR2x2_ASAP7_75t_L g756 ( 
.A(n_610),
.B(n_532),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_690),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_684),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_676),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_676),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_681),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_681),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_682),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_682),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_648),
.B(n_516),
.Y(n_765)
);

NAND2xp33_ASAP7_75t_R g766 ( 
.A(n_643),
.B(n_572),
.Y(n_766)
);

XNOR2xp5_ASAP7_75t_L g767 ( 
.A(n_643),
.B(n_556),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_689),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_694),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_634),
.Y(n_770)
);

AND2x6_ASAP7_75t_L g771 ( 
.A(n_696),
.B(n_531),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_615),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_650),
.B(n_549),
.Y(n_773)
);

NAND2x1p5_ASAP7_75t_L g774 ( 
.A(n_697),
.B(n_527),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_634),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_661),
.Y(n_776)
);

NOR2xp67_ASAP7_75t_L g777 ( 
.A(n_653),
.B(n_580),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_732),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_751),
.B(n_685),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_719),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_719),
.B(n_572),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_748),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_704),
.Y(n_783)
);

INVx4_ASAP7_75t_L g784 ( 
.A(n_727),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_735),
.B(n_680),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_711),
.B(n_627),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_735),
.B(n_666),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_732),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_726),
.B(n_664),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_727),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_698),
.B(n_661),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_698),
.B(n_670),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_757),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_753),
.B(n_625),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_699),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_729),
.A2(n_484),
.B(n_674),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_700),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_701),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_705),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_741),
.B(n_646),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_716),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_718),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_738),
.A2(n_518),
.B(n_505),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_724),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_755),
.B(n_656),
.Y(n_805)
);

INVx4_ASAP7_75t_L g806 ( 
.A(n_754),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_720),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_707),
.B(n_629),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_721),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_758),
.B(n_598),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_706),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_752),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_703),
.B(n_608),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_709),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_722),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_710),
.A2(n_518),
.B(n_569),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_749),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_749),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_725),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_710),
.B(n_642),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_744),
.B(n_747),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_757),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_742),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_728),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_743),
.Y(n_825)
);

INVxp67_ASAP7_75t_L g826 ( 
.A(n_723),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_712),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_730),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_733),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_713),
.Y(n_830)
);

INVx1_ASAP7_75t_SL g831 ( 
.A(n_750),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_702),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_774),
.B(n_608),
.Y(n_833)
);

INVx1_ASAP7_75t_SL g834 ( 
.A(n_773),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_774),
.B(n_591),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_717),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_734),
.B(n_527),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_737),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_739),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_760),
.B(n_768),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_740),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_760),
.B(n_525),
.Y(n_842)
);

INVx4_ASAP7_75t_L g843 ( 
.A(n_771),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_772),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_765),
.B(n_692),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_708),
.Y(n_846)
);

OR2x2_ASAP7_75t_SL g847 ( 
.A(n_764),
.B(n_618),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_765),
.B(n_547),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_745),
.B(n_591),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_771),
.B(n_594),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_766),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_768),
.Y(n_852)
);

AND2x6_ASAP7_75t_L g853 ( 
.A(n_759),
.B(n_761),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_771),
.B(n_594),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_776),
.B(n_647),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_764),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_776),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_736),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_762),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_817),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_803),
.B(n_771),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_SL g862 ( 
.A(n_843),
.B(n_714),
.Y(n_862)
);

NOR2xp67_ASAP7_75t_L g863 ( 
.A(n_843),
.B(n_736),
.Y(n_863)
);

BUFx2_ASAP7_75t_L g864 ( 
.A(n_822),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_821),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_817),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_856),
.Y(n_867)
);

NAND2x1p5_ASAP7_75t_L g868 ( 
.A(n_843),
.B(n_763),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_817),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_789),
.B(n_771),
.Y(n_870)
);

OR2x6_ASAP7_75t_L g871 ( 
.A(n_846),
.B(n_647),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_857),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_784),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_823),
.B(n_777),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_848),
.B(n_715),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_800),
.B(n_769),
.Y(n_876)
);

AND2x6_ASAP7_75t_L g877 ( 
.A(n_791),
.B(n_792),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_793),
.B(n_812),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_779),
.B(n_770),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_859),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_857),
.B(n_775),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_857),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_823),
.B(n_714),
.Y(n_883)
);

NAND2x1p5_ASAP7_75t_L g884 ( 
.A(n_806),
.B(n_506),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_786),
.B(n_756),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_817),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_783),
.Y(n_887)
);

AND2x6_ASAP7_75t_L g888 ( 
.A(n_791),
.B(n_655),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_818),
.Y(n_889)
);

BUFx12f_ASAP7_75t_L g890 ( 
.A(n_818),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_818),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_851),
.B(n_746),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_782),
.B(n_533),
.Y(n_893)
);

INVx6_ASAP7_75t_L g894 ( 
.A(n_818),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_780),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_846),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_804),
.B(n_493),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_785),
.B(n_655),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_852),
.Y(n_899)
);

NAND2x1p5_ASAP7_75t_L g900 ( 
.A(n_806),
.B(n_784),
.Y(n_900)
);

OR2x6_ASAP7_75t_L g901 ( 
.A(n_792),
.B(n_677),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_852),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_790),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_778),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_780),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_780),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_795),
.Y(n_907)
);

INVx8_ASAP7_75t_L g908 ( 
.A(n_853),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_858),
.B(n_486),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_841),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_834),
.B(n_493),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_825),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_788),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_830),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_795),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_798),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_SL g917 ( 
.A(n_794),
.B(n_644),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_798),
.Y(n_918)
);

INVx1_ASAP7_75t_SL g919 ( 
.A(n_840),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_787),
.B(n_510),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_799),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_825),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_890),
.Y(n_923)
);

BUFx2_ASAP7_75t_SL g924 ( 
.A(n_860),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_867),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_878),
.Y(n_926)
);

INVx4_ASAP7_75t_L g927 ( 
.A(n_860),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_883),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_883),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_887),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_860),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_896),
.Y(n_932)
);

BUFx6f_ASAP7_75t_SL g933 ( 
.A(n_901),
.Y(n_933)
);

CKINVDCx16_ASAP7_75t_R g934 ( 
.A(n_917),
.Y(n_934)
);

BUFx8_ASAP7_75t_L g935 ( 
.A(n_864),
.Y(n_935)
);

BUFx16f_ASAP7_75t_R g936 ( 
.A(n_874),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_911),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_880),
.Y(n_938)
);

BUFx5_ASAP7_75t_L g939 ( 
.A(n_872),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_869),
.Y(n_940)
);

BUFx8_ASAP7_75t_L g941 ( 
.A(n_892),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_869),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_870),
.B(n_813),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_910),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_875),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_882),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_866),
.B(n_842),
.Y(n_947)
);

CKINVDCx16_ASAP7_75t_R g948 ( 
.A(n_917),
.Y(n_948)
);

BUFx5_ASAP7_75t_L g949 ( 
.A(n_916),
.Y(n_949)
);

BUFx5_ASAP7_75t_L g950 ( 
.A(n_921),
.Y(n_950)
);

INVx5_ASAP7_75t_L g951 ( 
.A(n_869),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_886),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_922),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_919),
.Y(n_954)
);

NAND2x1p5_ASAP7_75t_L g955 ( 
.A(n_912),
.B(n_844),
.Y(n_955)
);

BUFx10_ASAP7_75t_L g956 ( 
.A(n_909),
.Y(n_956)
);

CKINVDCx11_ASAP7_75t_R g957 ( 
.A(n_901),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_886),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_889),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_889),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_914),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_891),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_891),
.Y(n_963)
);

INVxp67_ASAP7_75t_SL g964 ( 
.A(n_873),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_914),
.Y(n_965)
);

INVx6_ASAP7_75t_L g966 ( 
.A(n_894),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_881),
.Y(n_967)
);

NAND2x1p5_ASAP7_75t_L g968 ( 
.A(n_912),
.B(n_922),
.Y(n_968)
);

INVx3_ASAP7_75t_SL g969 ( 
.A(n_901),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_894),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_897),
.B(n_820),
.Y(n_971)
);

BUFx4f_ASAP7_75t_L g972 ( 
.A(n_877),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_881),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_895),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_907),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_919),
.Y(n_976)
);

INVx5_ASAP7_75t_L g977 ( 
.A(n_922),
.Y(n_977)
);

INVx3_ASAP7_75t_SL g978 ( 
.A(n_885),
.Y(n_978)
);

BUFx12f_ASAP7_75t_L g979 ( 
.A(n_871),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_930),
.Y(n_980)
);

INVx4_ASAP7_75t_L g981 ( 
.A(n_977),
.Y(n_981)
);

BUFx12f_ASAP7_75t_L g982 ( 
.A(n_957),
.Y(n_982)
);

AOI21xp33_ASAP7_75t_SL g983 ( 
.A1(n_934),
.A2(n_845),
.B(n_826),
.Y(n_983)
);

BUFx10_ASAP7_75t_L g984 ( 
.A(n_923),
.Y(n_984)
);

OAI22xp33_ASAP7_75t_L g985 ( 
.A1(n_945),
.A2(n_862),
.B1(n_865),
.B2(n_858),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_925),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_930),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_967),
.A2(n_879),
.B1(n_876),
.B2(n_898),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_974),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_946),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_946),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_971),
.A2(n_805),
.B1(n_858),
.B2(n_870),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_938),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_928),
.A2(n_805),
.B1(n_858),
.B2(n_808),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_967),
.B(n_876),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_SL g996 ( 
.A1(n_948),
.A2(n_862),
.B1(n_888),
.B2(n_871),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_973),
.B(n_943),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_937),
.B(n_831),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_975),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_SL g1000 ( 
.A1(n_948),
.A2(n_888),
.B1(n_871),
.B2(n_820),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_929),
.A2(n_808),
.B1(n_816),
.B2(n_893),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_973),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_977),
.Y(n_1003)
);

OAI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_978),
.A2(n_865),
.B1(n_898),
.B2(n_879),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_SL g1005 ( 
.A1(n_941),
.A2(n_888),
.B1(n_796),
.B2(n_861),
.Y(n_1005)
);

OAI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_926),
.A2(n_766),
.B1(n_833),
.B2(n_861),
.Y(n_1006)
);

BUFx8_ASAP7_75t_L g1007 ( 
.A(n_933),
.Y(n_1007)
);

INVx6_ASAP7_75t_L g1008 ( 
.A(n_935),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_961),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_935),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_932),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_965),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_972),
.A2(n_863),
.B1(n_873),
.B2(n_900),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_965),
.Y(n_1014)
);

BUFx5_ASAP7_75t_L g1015 ( 
.A(n_952),
.Y(n_1015)
);

INVx6_ASAP7_75t_L g1016 ( 
.A(n_941),
.Y(n_1016)
);

CKINVDCx11_ASAP7_75t_R g1017 ( 
.A(n_969),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_956),
.Y(n_1018)
);

INVx1_ASAP7_75t_SL g1019 ( 
.A(n_954),
.Y(n_1019)
);

INVx6_ASAP7_75t_L g1020 ( 
.A(n_966),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_944),
.Y(n_1021)
);

INVx6_ASAP7_75t_L g1022 ( 
.A(n_966),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_976),
.Y(n_1023)
);

INVx6_ASAP7_75t_L g1024 ( 
.A(n_979),
.Y(n_1024)
);

INVx6_ASAP7_75t_L g1025 ( 
.A(n_956),
.Y(n_1025)
);

INVxp67_ASAP7_75t_SL g1026 ( 
.A(n_964),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_976),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_970),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_949),
.Y(n_1029)
);

BUFx10_ASAP7_75t_L g1030 ( 
.A(n_947),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_987),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_991),
.Y(n_1032)
);

BUFx8_ASAP7_75t_SL g1033 ( 
.A(n_1010),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_1004),
.A2(n_943),
.B1(n_583),
.B2(n_590),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_980),
.Y(n_1035)
);

OAI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_983),
.A2(n_854),
.B1(n_850),
.B2(n_835),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_995),
.B(n_947),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_996),
.A2(n_868),
.B1(n_847),
.B2(n_955),
.Y(n_1038)
);

OAI222xp33_ASAP7_75t_L g1039 ( 
.A1(n_1005),
.A2(n_602),
.B1(n_590),
.B2(n_586),
.C1(n_920),
.C2(n_903),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_990),
.Y(n_1040)
);

OAI222xp33_ASAP7_75t_L g1041 ( 
.A1(n_1000),
.A2(n_602),
.B1(n_586),
.B2(n_920),
.C1(n_913),
.C2(n_904),
.Y(n_1041)
);

OAI222xp33_ASAP7_75t_L g1042 ( 
.A1(n_1000),
.A2(n_936),
.B1(n_918),
.B2(n_915),
.C1(n_567),
.C2(n_606),
.Y(n_1042)
);

INVx1_ASAP7_75t_SL g1043 ( 
.A(n_1027),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_988),
.A2(n_837),
.B1(n_567),
.B2(n_509),
.Y(n_1044)
);

OAI222xp33_ASAP7_75t_L g1045 ( 
.A1(n_985),
.A2(n_936),
.B1(n_767),
.B2(n_797),
.C1(n_902),
.C2(n_899),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_1020),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_997),
.B(n_855),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_SL g1048 ( 
.A1(n_1016),
.A2(n_950),
.B1(n_949),
.B2(n_908),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1009),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_1006),
.A2(n_811),
.B1(n_814),
.B2(n_810),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_1001),
.A2(n_951),
.B1(n_895),
.B2(n_905),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_SL g1052 ( 
.A1(n_1016),
.A2(n_950),
.B1(n_949),
.B2(n_908),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1012),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_993),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_999),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_994),
.A2(n_1019),
.B1(n_992),
.B2(n_1018),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1002),
.Y(n_1057)
);

OR2x2_ASAP7_75t_SL g1058 ( 
.A(n_1008),
.B(n_824),
.Y(n_1058)
);

AOI21xp33_ASAP7_75t_L g1059 ( 
.A1(n_1023),
.A2(n_802),
.B(n_801),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_1021),
.A2(n_824),
.B1(n_819),
.B2(n_809),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_1022),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1014),
.Y(n_1062)
);

OAI21xp33_ASAP7_75t_L g1063 ( 
.A1(n_998),
.A2(n_829),
.B(n_828),
.Y(n_1063)
);

BUFx8_ASAP7_75t_SL g1064 ( 
.A(n_982),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_1007),
.A2(n_604),
.B1(n_593),
.B2(n_555),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_986),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1026),
.Y(n_1067)
);

OAI21xp33_ASAP7_75t_L g1068 ( 
.A1(n_1011),
.A2(n_781),
.B(n_849),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1015),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1015),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1015),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_1028),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_1017),
.A2(n_1024),
.B1(n_1025),
.B2(n_555),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_1024),
.A2(n_564),
.B1(n_565),
.B2(n_546),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1015),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1015),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_989),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_1025),
.A2(n_564),
.B1(n_565),
.B2(n_546),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1031),
.B(n_1029),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_1036),
.B(n_1013),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1057),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_SL g1082 ( 
.A1(n_1038),
.A2(n_1030),
.B1(n_981),
.B2(n_1003),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1058),
.A2(n_981),
.B1(n_968),
.B2(n_906),
.Y(n_1083)
);

OAI221xp5_ASAP7_75t_L g1084 ( 
.A1(n_1065),
.A2(n_838),
.B1(n_884),
.B2(n_839),
.C(n_836),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_SL g1085 ( 
.A1(n_1056),
.A2(n_939),
.B1(n_924),
.B2(n_984),
.Y(n_1085)
);

NAND3xp33_ASAP7_75t_L g1086 ( 
.A(n_1034),
.B(n_566),
.C(n_565),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1040),
.Y(n_1087)
);

AOI221xp5_ASAP7_75t_L g1088 ( 
.A1(n_1039),
.A2(n_566),
.B1(n_568),
.B2(n_578),
.C(n_579),
.Y(n_1088)
);

AOI222xp33_ASAP7_75t_L g1089 ( 
.A1(n_1042),
.A2(n_781),
.B1(n_535),
.B2(n_536),
.C1(n_540),
.C2(n_603),
.Y(n_1089)
);

OAI22xp33_ASAP7_75t_SL g1090 ( 
.A1(n_1037),
.A2(n_1022),
.B1(n_906),
.B2(n_536),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1032),
.B(n_989),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1068),
.A2(n_827),
.B1(n_807),
.B2(n_815),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1049),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1063),
.A2(n_603),
.B1(n_605),
.B2(n_600),
.Y(n_1094)
);

AND2x2_ASAP7_75t_SL g1095 ( 
.A(n_1044),
.B(n_927),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1032),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1044),
.A2(n_939),
.B1(n_953),
.B2(n_832),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1055),
.B(n_974),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_1050),
.A2(n_582),
.B1(n_589),
.B2(n_597),
.Y(n_1099)
);

NAND3xp33_ASAP7_75t_L g1100 ( 
.A(n_1059),
.B(n_568),
.C(n_566),
.Y(n_1100)
);

OAI221xp5_ASAP7_75t_L g1101 ( 
.A1(n_1073),
.A2(n_540),
.B1(n_535),
.B2(n_603),
.C(n_594),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1050),
.A2(n_587),
.B1(n_589),
.B2(n_597),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1043),
.A2(n_582),
.B1(n_587),
.B2(n_609),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_SL g1104 ( 
.A1(n_1045),
.A2(n_958),
.B1(n_931),
.B2(n_962),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1066),
.A2(n_605),
.B1(n_600),
.B2(n_596),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1054),
.A2(n_579),
.B1(n_592),
.B2(n_578),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1067),
.A2(n_963),
.B1(n_931),
.B2(n_960),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1035),
.B(n_1053),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1072),
.A2(n_960),
.B1(n_959),
.B2(n_958),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1047),
.B(n_974),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1060),
.A2(n_960),
.B1(n_959),
.B2(n_942),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1074),
.A2(n_959),
.B1(n_942),
.B2(n_940),
.Y(n_1112)
);

AOI221xp5_ASAP7_75t_L g1113 ( 
.A1(n_1041),
.A2(n_596),
.B1(n_605),
.B2(n_600),
.C(n_561),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1051),
.A2(n_497),
.B1(n_731),
.B2(n_507),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_SL g1115 ( 
.A1(n_1069),
.A2(n_495),
.B1(n_491),
.B2(n_489),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1078),
.A2(n_489),
.B1(n_488),
.B2(n_82),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1062),
.B(n_79),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1062),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1070),
.Y(n_1119)
);

OAI221xp5_ASAP7_75t_L g1120 ( 
.A1(n_1048),
.A2(n_79),
.B1(n_81),
.B2(n_84),
.C(n_85),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1108),
.B(n_1079),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1108),
.B(n_1071),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_1090),
.B(n_1052),
.Y(n_1123)
);

AOI221xp5_ASAP7_75t_L g1124 ( 
.A1(n_1120),
.A2(n_1077),
.B1(n_1075),
.B2(n_1061),
.C(n_1046),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1081),
.B(n_1076),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_1113),
.B(n_1088),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1087),
.B(n_85),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1104),
.A2(n_1033),
.B1(n_1064),
.B2(n_88),
.Y(n_1128)
);

NOR3xp33_ASAP7_75t_SL g1129 ( 
.A(n_1101),
.B(n_89),
.C(n_98),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1091),
.B(n_288),
.Y(n_1130)
);

OA21x2_ASAP7_75t_L g1131 ( 
.A1(n_1080),
.A2(n_101),
.B(n_102),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1082),
.B(n_103),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1093),
.B(n_104),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_1085),
.B(n_114),
.Y(n_1134)
);

OAI221xp5_ASAP7_75t_L g1135 ( 
.A1(n_1105),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.C(n_122),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1110),
.B(n_125),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1119),
.B(n_129),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1119),
.B(n_132),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_L g1139 ( 
.A(n_1089),
.B(n_133),
.C(n_135),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1096),
.B(n_141),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1118),
.B(n_147),
.Y(n_1141)
);

NAND4xp25_ASAP7_75t_L g1142 ( 
.A(n_1117),
.B(n_148),
.C(n_149),
.D(n_150),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1095),
.B(n_153),
.Y(n_1143)
);

NAND2xp33_ASAP7_75t_SL g1144 ( 
.A(n_1083),
.B(n_157),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1095),
.B(n_158),
.Y(n_1145)
);

OAI221xp5_ASAP7_75t_L g1146 ( 
.A1(n_1103),
.A2(n_160),
.B1(n_164),
.B2(n_166),
.C(n_167),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1098),
.B(n_168),
.Y(n_1147)
);

OAI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1086),
.A2(n_171),
.B1(n_172),
.B2(n_176),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_L g1149 ( 
.A(n_1094),
.B(n_1107),
.C(n_1106),
.Y(n_1149)
);

NOR3xp33_ASAP7_75t_L g1150 ( 
.A(n_1132),
.B(n_1100),
.C(n_1084),
.Y(n_1150)
);

NAND3xp33_ASAP7_75t_L g1151 ( 
.A(n_1129),
.B(n_1116),
.C(n_1109),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1121),
.B(n_1114),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_1122),
.B(n_1111),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_1125),
.Y(n_1154)
);

INVx1_ASAP7_75t_SL g1155 ( 
.A(n_1127),
.Y(n_1155)
);

NAND3xp33_ASAP7_75t_L g1156 ( 
.A(n_1124),
.B(n_1097),
.C(n_1092),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1130),
.B(n_1137),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1131),
.B(n_1137),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1138),
.B(n_1112),
.Y(n_1159)
);

NAND3xp33_ASAP7_75t_L g1160 ( 
.A(n_1139),
.B(n_1115),
.C(n_1099),
.Y(n_1160)
);

NOR2x1_ASAP7_75t_L g1161 ( 
.A(n_1131),
.B(n_1102),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1133),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1126),
.A2(n_191),
.B(n_195),
.Y(n_1163)
);

NAND3xp33_ASAP7_75t_SL g1164 ( 
.A(n_1128),
.B(n_1143),
.C(n_1145),
.Y(n_1164)
);

NAND3xp33_ASAP7_75t_L g1165 ( 
.A(n_1123),
.B(n_197),
.C(n_199),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1145),
.A2(n_201),
.B(n_203),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1136),
.B(n_205),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1155),
.B(n_1140),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1154),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1154),
.B(n_1141),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1158),
.Y(n_1171)
);

XOR2x2_ASAP7_75t_L g1172 ( 
.A(n_1164),
.B(n_1134),
.Y(n_1172)
);

XOR2x2_ASAP7_75t_L g1173 ( 
.A(n_1166),
.B(n_1134),
.Y(n_1173)
);

NAND4xp75_ASAP7_75t_L g1174 ( 
.A(n_1163),
.B(n_1161),
.C(n_1166),
.D(n_1131),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_1162),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_1157),
.Y(n_1176)
);

XNOR2x2_ASAP7_75t_L g1177 ( 
.A(n_1165),
.B(n_1142),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1153),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1150),
.A2(n_1144),
.B1(n_1149),
.B2(n_1135),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_1159),
.Y(n_1180)
);

XOR2x2_ASAP7_75t_L g1181 ( 
.A(n_1172),
.B(n_1151),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1175),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1178),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1176),
.Y(n_1184)
);

XOR2x2_ASAP7_75t_L g1185 ( 
.A(n_1173),
.B(n_1156),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1180),
.B(n_1152),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1169),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1171),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1168),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_1170),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1185),
.A2(n_1181),
.B1(n_1174),
.B2(n_1179),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1183),
.Y(n_1192)
);

XOR2x2_ASAP7_75t_L g1193 ( 
.A(n_1185),
.B(n_1177),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_1186),
.Y(n_1194)
);

XOR2x2_ASAP7_75t_L g1195 ( 
.A(n_1184),
.B(n_1160),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1190),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1188),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1196),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1194),
.Y(n_1199)
);

OAI322xp33_ASAP7_75t_L g1200 ( 
.A1(n_1191),
.A2(n_1189),
.A3(n_1187),
.B1(n_1182),
.B2(n_1148),
.C1(n_1167),
.C2(n_1146),
.Y(n_1200)
);

AO22x1_ASAP7_75t_L g1201 ( 
.A1(n_1193),
.A2(n_1147),
.B1(n_1144),
.B2(n_209),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1192),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_1199),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1202),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1203),
.Y(n_1205)
);

AOI221xp5_ASAP7_75t_L g1206 ( 
.A1(n_1204),
.A2(n_1200),
.B1(n_1198),
.B2(n_1201),
.C(n_1197),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1206),
.B(n_1195),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1205),
.B(n_210),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1207),
.A2(n_211),
.B1(n_218),
.B2(n_219),
.Y(n_1209)
);

BUFx8_ASAP7_75t_L g1210 ( 
.A(n_1208),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1210),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1209),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1211),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_1212),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1213),
.Y(n_1215)
);

AO22x2_ASAP7_75t_L g1216 ( 
.A1(n_1214),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1216),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1215),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1216),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_SL g1220 ( 
.A1(n_1219),
.A2(n_242),
.B1(n_243),
.B2(n_246),
.Y(n_1220)
);

AO22x2_ASAP7_75t_L g1221 ( 
.A1(n_1217),
.A2(n_248),
.B1(n_250),
.B2(n_252),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1221),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1220),
.Y(n_1223)
);

OAI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1223),
.A2(n_1218),
.B1(n_254),
.B2(n_256),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1222),
.A2(n_253),
.B1(n_257),
.B2(n_258),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1224),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1225),
.Y(n_1227)
);

AOI221xp5_ASAP7_75t_L g1228 ( 
.A1(n_1226),
.A2(n_265),
.B1(n_269),
.B2(n_272),
.C(n_273),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1228),
.A2(n_1227),
.B1(n_275),
.B2(n_277),
.Y(n_1229)
);


endmodule