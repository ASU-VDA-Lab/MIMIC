module fake_netlist_5_2311_n_1411 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1411);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1411;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_292;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1314;
wire n_709;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_308;
wire n_297;
wire n_1078;
wire n_775;
wire n_219;
wire n_600;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_196;
wire n_215;
wire n_646;
wire n_436;
wire n_1394;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1322;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_324;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_252;
wire n_624;
wire n_1380;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_256;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1096;
wire n_234;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_733;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_221;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_236;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_229;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_246;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_566;
wire n_565;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g182 ( 
.A(n_85),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_32),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_89),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_101),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_81),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_139),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_8),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_69),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_11),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_6),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_77),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_137),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_13),
.Y(n_198)
);

BUFx2_ASAP7_75t_SL g199 ( 
.A(n_141),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_110),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_37),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_106),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_96),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_9),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_150),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_105),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_118),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_27),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_1),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_32),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_9),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_143),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_180),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_88),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_10),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_18),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_99),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_149),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_25),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_36),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_129),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_79),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_45),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_87),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_131),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_43),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_145),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_114),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_160),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_59),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_90),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_73),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_75),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_174),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_172),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_83),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_127),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_82),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_28),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_108),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_5),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_78),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_37),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_170),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_38),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_102),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_42),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_119),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_152),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_86),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_148),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_69),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_47),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_93),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_176),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_159),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_3),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_138),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_147),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_157),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_66),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_113),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_84),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_104),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_167),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_58),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_61),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_171),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_48),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_120),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_153),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_13),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_133),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_10),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_173),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_128),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_155),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_134),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_161),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_76),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_54),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_20),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_41),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_91),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_181),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_100),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_55),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_42),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_5),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_140),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_156),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_47),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_27),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_56),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_92),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_15),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_158),
.Y(n_301)
);

BUFx2_ASAP7_75t_SL g302 ( 
.A(n_109),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_0),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_51),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_151),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_125),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_7),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_116),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_142),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_57),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_20),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_126),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_130),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_94),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_12),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_31),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_63),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_61),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_121),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_64),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_12),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_220),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_212),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_212),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_223),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_212),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_275),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_243),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_212),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_212),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_208),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_208),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_227),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_203),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_209),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_228),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_214),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_230),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_233),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_209),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_0),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_273),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_279),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_252),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_315),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_232),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_216),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_253),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_238),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_299),
.Y(n_350)
);

INVxp33_ASAP7_75t_L g351 ( 
.A(n_204),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_273),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_205),
.B(n_2),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_239),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_312),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_300),
.Y(n_356)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_184),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_240),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_241),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_251),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_244),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_251),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_246),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_305),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_248),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_205),
.B(n_2),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_310),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_263),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_198),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_201),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_267),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_245),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_247),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_268),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_257),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_278),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_269),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_245),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_272),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_285),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_282),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_283),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_296),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_284),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_307),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_217),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_311),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_276),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_188),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_218),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_221),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_305),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_276),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_188),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_235),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_222),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_235),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_190),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_236),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_245),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_306),
.B(n_3),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_226),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_236),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_182),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_260),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_260),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_323),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_347),
.B(n_306),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_323),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_324),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_405),
.B(n_309),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_324),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_334),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_326),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_356),
.A2(n_298),
.B1(n_304),
.B2(n_256),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_322),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_325),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_333),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_336),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_364),
.B(n_309),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_338),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_328),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_326),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_329),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_329),
.Y(n_428)
);

AND2x6_ASAP7_75t_L g429 ( 
.A(n_347),
.B(n_197),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_396),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_346),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_396),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_398),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_398),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_349),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_400),
.Y(n_436)
);

NOR2xp67_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_183),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_354),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_358),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_361),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_SL g441 ( 
.A(n_351),
.B(n_191),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_404),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_404),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_393),
.B(n_185),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_360),
.B(n_186),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_407),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_407),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_406),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_406),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_390),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_363),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_370),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_365),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_360),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_370),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_353),
.B(n_190),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_331),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_362),
.B(n_187),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_369),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_371),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_375),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_331),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_332),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_378),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_332),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_339),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_387),
.B(n_189),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_371),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_335),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_380),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_383),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_359),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_341),
.B(n_271),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_335),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_340),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_340),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_362),
.B(n_194),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_423),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g479 ( 
.A(n_444),
.B(n_197),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_444),
.B(n_197),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_467),
.B(n_391),
.Y(n_481)
);

AO22x2_ASAP7_75t_L g482 ( 
.A1(n_456),
.A2(n_327),
.B1(n_265),
.B2(n_210),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_473),
.B(n_337),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_426),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_429),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_458),
.B(n_477),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_425),
.B(n_344),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_426),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_426),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_408),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_416),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_427),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_473),
.B(n_348),
.Y(n_493)
);

AND2x2_ASAP7_75t_SL g494 ( 
.A(n_456),
.B(n_197),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_427),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_412),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_458),
.B(n_219),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_423),
.B(n_392),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_419),
.B(n_397),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_408),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_429),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_423),
.B(n_444),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_410),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_445),
.B(n_367),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_458),
.B(n_225),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_412),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_410),
.Y(n_507)
);

AO22x2_ASAP7_75t_L g508 ( 
.A1(n_413),
.A2(n_231),
.B1(n_259),
.B2(n_242),
.Y(n_508)
);

AO22x2_ASAP7_75t_L g509 ( 
.A1(n_413),
.A2(n_264),
.B1(n_274),
.B2(n_266),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_425),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_412),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_445),
.B(n_403),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_441),
.B(n_379),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_420),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_411),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_412),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_427),
.Y(n_517)
);

BUFx10_ASAP7_75t_L g518 ( 
.A(n_421),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_422),
.B(n_345),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_424),
.B(n_372),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_428),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_431),
.B(n_382),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_435),
.B(n_438),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_428),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_411),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_439),
.B(n_385),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_440),
.B(n_395),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_451),
.B(n_453),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_458),
.B(n_277),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_414),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_459),
.B(n_399),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_454),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_461),
.B(n_355),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_428),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_462),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_464),
.B(n_470),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_414),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_417),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_471),
.B(n_373),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_477),
.B(n_401),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_445),
.B(n_366),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_478),
.B(n_472),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_490),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_490),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_494),
.B(n_477),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_500),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_494),
.B(n_478),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_500),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_494),
.B(n_477),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_502),
.B(n_454),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_503),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_481),
.B(n_343),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_498),
.B(n_454),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_541),
.B(n_409),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_512),
.B(n_196),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_499),
.B(n_539),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_483),
.B(n_196),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_488),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_504),
.B(n_452),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_503),
.B(n_507),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_487),
.B(n_350),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_488),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_488),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_532),
.B(n_409),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_489),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_489),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_532),
.B(n_442),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_487),
.B(n_493),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_507),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_482),
.A2(n_402),
.B1(n_321),
.B2(n_418),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_532),
.B(n_442),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_515),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_486),
.B(n_442),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_486),
.B(n_442),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_486),
.B(n_417),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_508),
.A2(n_418),
.B1(n_255),
.B2(n_313),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_489),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_486),
.B(n_200),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_504),
.B(n_452),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_515),
.B(n_465),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_525),
.B(n_530),
.Y(n_581)
);

NAND2x1_ASAP7_75t_L g582 ( 
.A(n_485),
.B(n_429),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_492),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_525),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_530),
.B(n_537),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_492),
.Y(n_586)
);

INVx8_ASAP7_75t_L g587 ( 
.A(n_479),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_492),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_508),
.A2(n_437),
.B1(n_460),
.B2(n_455),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_535),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_537),
.B(n_465),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_538),
.B(n_465),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_538),
.B(n_465),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_508),
.A2(n_199),
.B1(n_302),
.B2(n_281),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_495),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_497),
.A2(n_437),
.B(n_429),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_514),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_508),
.A2(n_294),
.B1(n_295),
.B2(n_280),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_495),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_519),
.B(n_200),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_495),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_535),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_497),
.B(n_474),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_540),
.B(n_513),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_509),
.A2(n_460),
.B1(n_468),
.B2(n_314),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_497),
.B(n_474),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_497),
.B(n_474),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_517),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_482),
.B(n_468),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_485),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_482),
.B(n_367),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_517),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_505),
.B(n_474),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_505),
.B(n_462),
.Y(n_614)
);

NAND2x1_ASAP7_75t_L g615 ( 
.A(n_485),
.B(n_429),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_517),
.Y(n_616)
);

INVxp67_ASAP7_75t_SL g617 ( 
.A(n_535),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_505),
.B(n_462),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_513),
.B(n_450),
.Y(n_619)
);

O2A1O1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_505),
.A2(n_433),
.B(n_436),
.C(n_434),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_510),
.Y(n_621)
);

OR2x6_ASAP7_75t_L g622 ( 
.A(n_509),
.B(n_197),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_529),
.B(n_462),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_521),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_521),
.Y(n_625)
);

A2O1A1Ixp33_ASAP7_75t_L g626 ( 
.A1(n_529),
.A2(n_433),
.B(n_436),
.C(n_434),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_553),
.B(n_529),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_621),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_556),
.B(n_536),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_550),
.B(n_529),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_621),
.Y(n_631)
);

OR2x6_ASAP7_75t_L g632 ( 
.A(n_587),
.B(n_509),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_587),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_559),
.B(n_510),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_559),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_SL g636 ( 
.A1(n_552),
.A2(n_466),
.B1(n_491),
.B2(n_450),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_597),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_595),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_547),
.A2(n_509),
.B1(n_479),
.B2(n_480),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_558),
.Y(n_640)
);

NOR3xp33_ASAP7_75t_SL g641 ( 
.A(n_570),
.B(n_192),
.C(n_191),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_579),
.B(n_485),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_545),
.A2(n_501),
.B(n_480),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_610),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_558),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_622),
.Y(n_646)
);

NOR3xp33_ASAP7_75t_SL g647 ( 
.A(n_570),
.B(n_193),
.C(n_192),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_568),
.B(n_520),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_579),
.B(n_518),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_604),
.B(n_522),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_561),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_622),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_558),
.Y(n_653)
);

BUFx4f_ASAP7_75t_SL g654 ( 
.A(n_542),
.Y(n_654)
);

NAND2x1p5_ASAP7_75t_L g655 ( 
.A(n_610),
.B(n_582),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_562),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_619),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_562),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_595),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_SL g660 ( 
.A1(n_576),
.A2(n_531),
.B1(n_526),
.B2(n_195),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_601),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_543),
.B(n_501),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_562),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_563),
.Y(n_664)
);

BUFx12f_ASAP7_75t_L g665 ( 
.A(n_611),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_601),
.Y(n_666)
);

NOR2xp67_ASAP7_75t_L g667 ( 
.A(n_549),
.B(n_501),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_R g668 ( 
.A(n_622),
.B(n_202),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_616),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_543),
.B(n_544),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_616),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_610),
.B(n_518),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_544),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_624),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_587),
.Y(n_675)
);

INVx5_ASAP7_75t_L g676 ( 
.A(n_610),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_620),
.A2(n_527),
.B(n_528),
.C(n_523),
.Y(n_677)
);

INVxp33_ASAP7_75t_L g678 ( 
.A(n_611),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_573),
.A2(n_501),
.B(n_496),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_605),
.B(n_518),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_624),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_554),
.B(n_479),
.Y(n_682)
);

AND2x6_ASAP7_75t_L g683 ( 
.A(n_589),
.B(n_511),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_563),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_587),
.B(n_533),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_546),
.B(n_479),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_563),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_565),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_565),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_565),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_605),
.B(n_518),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_566),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_622),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_566),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_587),
.Y(n_695)
);

AOI221xp5_ASAP7_75t_SL g696 ( 
.A1(n_609),
.A2(n_389),
.B1(n_394),
.B2(n_368),
.C(n_376),
.Y(n_696)
);

BUFx2_ASAP7_75t_L g697 ( 
.A(n_622),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_546),
.B(n_511),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_566),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_548),
.B(n_368),
.Y(n_700)
);

NOR3xp33_ASAP7_75t_SL g701 ( 
.A(n_555),
.B(n_195),
.C(n_193),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_594),
.A2(n_479),
.B1(n_480),
.B2(n_484),
.Y(n_702)
);

BUFx12f_ASAP7_75t_L g703 ( 
.A(n_609),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_548),
.B(n_479),
.Y(n_704)
);

BUFx4f_ASAP7_75t_L g705 ( 
.A(n_551),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_577),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_577),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_551),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_582),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_577),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_583),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_590),
.Y(n_712)
);

OR2x2_ASAP7_75t_SL g713 ( 
.A(n_576),
.B(n_389),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_583),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_557),
.B(n_357),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_583),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_586),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_569),
.B(n_479),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_600),
.B(n_202),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_569),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_578),
.Y(n_721)
);

OAI21x1_ASAP7_75t_L g722 ( 
.A1(n_679),
.A2(n_602),
.B(n_590),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_629),
.B(n_572),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_650),
.A2(n_560),
.B1(n_584),
.B2(n_572),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_676),
.A2(n_574),
.B(n_615),
.Y(n_725)
);

OAI21x1_ASAP7_75t_L g726 ( 
.A1(n_655),
.A2(n_643),
.B(n_640),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_670),
.Y(n_727)
);

OAI21x1_ASAP7_75t_L g728 ( 
.A1(n_655),
.A2(n_602),
.B(n_590),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_631),
.Y(n_729)
);

AO22x2_ASAP7_75t_L g730 ( 
.A1(n_680),
.A2(n_584),
.B1(n_560),
.B2(n_589),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_634),
.B(n_635),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_705),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_631),
.B(n_581),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_648),
.A2(n_705),
.B(n_670),
.C(n_719),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_657),
.B(n_700),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_676),
.A2(n_615),
.B(n_617),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_700),
.B(n_634),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_676),
.A2(n_618),
.B(n_614),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_705),
.Y(n_739)
);

OAI21x1_ASAP7_75t_L g740 ( 
.A1(n_655),
.A2(n_602),
.B(n_590),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_673),
.B(n_708),
.Y(n_741)
);

OAI21xp5_ASAP7_75t_L g742 ( 
.A1(n_630),
.A2(n_606),
.B(n_603),
.Y(n_742)
);

OAI21x1_ASAP7_75t_L g743 ( 
.A1(n_640),
.A2(n_602),
.B(n_623),
.Y(n_743)
);

AND3x4_ASAP7_75t_L g744 ( 
.A(n_641),
.B(n_588),
.C(n_586),
.Y(n_744)
);

A2O1A1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_720),
.A2(n_585),
.B(n_598),
.C(n_596),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_649),
.B(n_596),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_L g747 ( 
.A1(n_627),
.A2(n_613),
.B(n_607),
.Y(n_747)
);

AOI21x1_ASAP7_75t_L g748 ( 
.A1(n_682),
.A2(n_564),
.B(n_567),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_676),
.A2(n_642),
.B1(n_708),
.B2(n_673),
.Y(n_749)
);

AO31x2_ASAP7_75t_L g750 ( 
.A1(n_638),
.A2(n_626),
.A3(n_591),
.B(n_592),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_638),
.Y(n_751)
);

OAI21x1_ASAP7_75t_L g752 ( 
.A1(n_645),
.A2(n_571),
.B(n_580),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_649),
.B(n_575),
.Y(n_753)
);

AOI21x1_ASAP7_75t_L g754 ( 
.A1(n_659),
.A2(n_593),
.B(n_588),
.Y(n_754)
);

OAI222xp33_ASAP7_75t_L g755 ( 
.A1(n_691),
.A2(n_297),
.B1(n_211),
.B2(n_318),
.C1(n_317),
.C2(n_303),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_676),
.A2(n_506),
.B(n_496),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_L g757 ( 
.A1(n_642),
.A2(n_588),
.B(n_586),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_676),
.A2(n_506),
.B(n_496),
.Y(n_758)
);

OAI21xp5_ASAP7_75t_L g759 ( 
.A1(n_642),
.A2(n_608),
.B(n_599),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_628),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_720),
.B(n_599),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_659),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_645),
.Y(n_763)
);

OAI21xp5_ASAP7_75t_L g764 ( 
.A1(n_642),
.A2(n_608),
.B(n_599),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_653),
.Y(n_765)
);

BUFx12f_ASAP7_75t_L g766 ( 
.A(n_665),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_644),
.A2(n_506),
.B(n_496),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_644),
.A2(n_506),
.B(n_496),
.Y(n_768)
);

AOI21x1_ASAP7_75t_L g769 ( 
.A1(n_661),
.A2(n_625),
.B(n_612),
.Y(n_769)
);

OAI21x1_ASAP7_75t_L g770 ( 
.A1(n_653),
.A2(n_625),
.B(n_612),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_715),
.B(n_612),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_678),
.B(n_625),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_644),
.B(n_511),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_662),
.A2(n_506),
.B(n_496),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_646),
.B(n_394),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_721),
.B(n_480),
.Y(n_776)
);

AO31x2_ASAP7_75t_L g777 ( 
.A1(n_661),
.A2(n_521),
.A3(n_524),
.B(n_484),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_685),
.B(n_446),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_662),
.A2(n_506),
.B(n_511),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_656),
.A2(n_516),
.B(n_524),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_662),
.A2(n_516),
.B(n_534),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_709),
.Y(n_782)
);

AO31x2_ASAP7_75t_L g783 ( 
.A1(n_666),
.A2(n_534),
.A3(n_432),
.B(n_443),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_677),
.B(n_480),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_709),
.Y(n_785)
);

OAI21x1_ASAP7_75t_L g786 ( 
.A1(n_656),
.A2(n_516),
.B(n_443),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_637),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_637),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_662),
.A2(n_516),
.B(n_443),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_658),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_703),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_709),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_667),
.A2(n_432),
.B(n_430),
.Y(n_793)
);

OAI21x1_ASAP7_75t_L g794 ( 
.A1(n_658),
.A2(n_432),
.B(n_446),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_646),
.B(n_447),
.Y(n_795)
);

A2O1A1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_647),
.A2(n_292),
.B(n_211),
.C(n_287),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_703),
.B(n_447),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_698),
.B(n_666),
.Y(n_798)
);

OAI21x1_ASAP7_75t_L g799 ( 
.A1(n_663),
.A2(n_449),
.B(n_457),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_665),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_SL g801 ( 
.A1(n_651),
.A2(n_660),
.B1(n_636),
.B2(n_713),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_669),
.Y(n_802)
);

OAI21x1_ASAP7_75t_SL g803 ( 
.A1(n_686),
.A2(n_449),
.B(n_457),
.Y(n_803)
);

O2A1O1Ixp5_ASAP7_75t_L g804 ( 
.A1(n_672),
.A2(n_704),
.B(n_718),
.C(n_698),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_633),
.Y(n_805)
);

OAI21x1_ASAP7_75t_SL g806 ( 
.A1(n_639),
.A2(n_463),
.B(n_457),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_667),
.A2(n_448),
.B(n_430),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_698),
.B(n_480),
.Y(n_808)
);

AND2x6_ASAP7_75t_SL g809 ( 
.A(n_685),
.B(n_632),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_698),
.B(n_480),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_685),
.B(n_652),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_633),
.B(n_216),
.Y(n_812)
);

INVxp67_ASAP7_75t_SL g813 ( 
.A(n_712),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_811),
.B(n_685),
.Y(n_814)
);

AOI21x1_ASAP7_75t_L g815 ( 
.A1(n_754),
.A2(n_671),
.B(n_669),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_787),
.Y(n_816)
);

AO32x2_ASAP7_75t_L g817 ( 
.A1(n_724),
.A2(n_696),
.A3(n_713),
.B1(n_632),
.B2(n_683),
.Y(n_817)
);

AO21x2_ASAP7_75t_L g818 ( 
.A1(n_734),
.A2(n_674),
.B(n_671),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_769),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_L g820 ( 
.A1(n_734),
.A2(n_702),
.B(n_683),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_811),
.B(n_652),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_731),
.B(n_701),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_731),
.B(n_693),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_742),
.A2(n_747),
.B(n_784),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_782),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_729),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_788),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_753),
.B(n_674),
.Y(n_828)
);

AOI21x1_ASAP7_75t_L g829 ( 
.A1(n_748),
.A2(n_681),
.B(n_684),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_760),
.Y(n_830)
);

OAI21x1_ASAP7_75t_L g831 ( 
.A1(n_743),
.A2(n_681),
.B(n_664),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_763),
.Y(n_832)
);

OAI21x1_ASAP7_75t_L g833 ( 
.A1(n_743),
.A2(n_664),
.B(n_663),
.Y(n_833)
);

OAI21x1_ASAP7_75t_L g834 ( 
.A1(n_794),
.A2(n_692),
.B(n_687),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_788),
.Y(n_835)
);

OA21x2_ASAP7_75t_L g836 ( 
.A1(n_752),
.A2(n_688),
.B(n_684),
.Y(n_836)
);

OAI22xp33_ASAP7_75t_L g837 ( 
.A1(n_737),
.A2(n_654),
.B1(n_668),
.B2(n_632),
.Y(n_837)
);

A2O1A1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_723),
.A2(n_697),
.B(n_693),
.C(n_688),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_735),
.B(n_697),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_811),
.B(n_633),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_763),
.Y(n_841)
);

AO31x2_ASAP7_75t_L g842 ( 
.A1(n_745),
.A2(n_689),
.A3(n_694),
.B(n_690),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_732),
.B(n_739),
.Y(n_843)
);

OAI21x1_ASAP7_75t_L g844 ( 
.A1(n_794),
.A2(n_692),
.B(n_687),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_733),
.B(n_712),
.Y(n_845)
);

NAND3x1_ASAP7_75t_L g846 ( 
.A(n_775),
.B(n_376),
.C(n_374),
.Y(n_846)
);

AOI222xp33_ASAP7_75t_L g847 ( 
.A1(n_801),
.A2(n_303),
.B1(n_297),
.B2(n_317),
.C1(n_318),
.C2(n_293),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_736),
.A2(n_675),
.B(n_633),
.Y(n_848)
);

AO21x2_ASAP7_75t_L g849 ( 
.A1(n_803),
.A2(n_690),
.B(n_689),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_753),
.B(n_683),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_765),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_766),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_733),
.B(n_712),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_775),
.B(n_632),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_766),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_738),
.A2(n_675),
.B(n_633),
.Y(n_856)
);

AO31x2_ASAP7_75t_L g857 ( 
.A1(n_745),
.A2(n_710),
.A3(n_716),
.B(n_714),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_800),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_730),
.A2(n_683),
.B1(n_224),
.B2(n_237),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_730),
.A2(n_683),
.B1(n_224),
.B2(n_237),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_755),
.A2(n_384),
.B(n_388),
.C(n_381),
.Y(n_861)
);

CKINVDCx14_ASAP7_75t_R g862 ( 
.A(n_791),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_727),
.B(n_694),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_741),
.A2(n_675),
.B1(n_695),
.B2(n_709),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_795),
.B(n_271),
.Y(n_865)
);

AOI21x1_ASAP7_75t_L g866 ( 
.A1(n_812),
.A2(n_707),
.B(n_706),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_765),
.Y(n_867)
);

OA21x2_ASAP7_75t_L g868 ( 
.A1(n_752),
.A2(n_707),
.B(n_706),
.Y(n_868)
);

NAND2x1p5_ASAP7_75t_L g869 ( 
.A(n_732),
.B(n_675),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_795),
.Y(n_870)
);

INVx8_ASAP7_75t_L g871 ( 
.A(n_797),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_782),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_746),
.B(n_710),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_790),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_797),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_797),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_751),
.Y(n_877)
);

CKINVDCx6p67_ASAP7_75t_R g878 ( 
.A(n_797),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_772),
.B(n_271),
.Y(n_879)
);

CKINVDCx11_ASAP7_75t_R g880 ( 
.A(n_809),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_782),
.Y(n_881)
);

AO21x1_ASAP7_75t_L g882 ( 
.A1(n_812),
.A2(n_714),
.B(n_711),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_762),
.Y(n_883)
);

AO31x2_ASAP7_75t_L g884 ( 
.A1(n_749),
.A2(n_716),
.A3(n_711),
.B(n_717),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_730),
.A2(n_683),
.B1(n_237),
.B2(n_224),
.Y(n_885)
);

AOI21x1_ASAP7_75t_L g886 ( 
.A1(n_771),
.A2(n_717),
.B(n_699),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_804),
.A2(n_683),
.B(n_699),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_802),
.Y(n_888)
);

CKINVDCx6p67_ASAP7_75t_R g889 ( 
.A(n_805),
.Y(n_889)
);

AO21x2_ASAP7_75t_L g890 ( 
.A1(n_726),
.A2(n_352),
.B(n_342),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_746),
.A2(n_695),
.B1(n_675),
.B2(n_709),
.Y(n_891)
);

OR2x6_ASAP7_75t_L g892 ( 
.A(n_739),
.B(n_695),
.Y(n_892)
);

OR2x6_ASAP7_75t_L g893 ( 
.A(n_778),
.B(n_695),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_725),
.A2(n_695),
.B(n_448),
.Y(n_894)
);

OAI21x1_ASAP7_75t_L g895 ( 
.A1(n_799),
.A2(n_475),
.B(n_463),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_772),
.B(n_463),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_756),
.A2(n_448),
.B(n_430),
.Y(n_897)
);

OAI21x1_ASAP7_75t_SL g898 ( 
.A1(n_806),
.A2(n_476),
.B(n_475),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_758),
.A2(n_448),
.B(n_430),
.Y(n_899)
);

AND2x6_ASAP7_75t_L g900 ( 
.A(n_785),
.B(n_374),
.Y(n_900)
);

OAI21x1_ASAP7_75t_L g901 ( 
.A1(n_799),
.A2(n_476),
.B(n_475),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_790),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_798),
.Y(n_903)
);

NAND2x1p5_ASAP7_75t_L g904 ( 
.A(n_805),
.B(n_476),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_778),
.A2(n_316),
.B1(n_377),
.B2(n_381),
.Y(n_905)
);

OAI21x1_ASAP7_75t_L g906 ( 
.A1(n_728),
.A2(n_352),
.B(n_342),
.Y(n_906)
);

NAND3xp33_ASAP7_75t_L g907 ( 
.A(n_796),
.B(n_234),
.C(n_229),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_778),
.A2(n_744),
.B1(n_776),
.B2(n_316),
.Y(n_908)
);

AOI221xp5_ASAP7_75t_L g909 ( 
.A1(n_796),
.A2(n_287),
.B1(n_291),
.B2(n_292),
.C(n_249),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_757),
.A2(n_429),
.B(n_207),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_805),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_761),
.A2(n_388),
.B1(n_377),
.B2(n_384),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_759),
.A2(n_386),
.B1(n_216),
.B2(n_261),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_783),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_SL g915 ( 
.A1(n_808),
.A2(n_386),
.B(n_216),
.C(n_7),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_805),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_728),
.A2(n_216),
.B(n_412),
.Y(n_917)
);

OR2x6_ASAP7_75t_L g918 ( 
.A(n_871),
.B(n_726),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_870),
.A2(n_764),
.B1(n_792),
.B2(n_785),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_877),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_883),
.Y(n_921)
);

AND2x2_ASAP7_75t_SL g922 ( 
.A(n_859),
.B(n_785),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_823),
.B(n_206),
.Y(n_923)
);

INVx4_ASAP7_75t_L g924 ( 
.A(n_911),
.Y(n_924)
);

BUFx12f_ASAP7_75t_L g925 ( 
.A(n_816),
.Y(n_925)
);

AOI221xp5_ASAP7_75t_L g926 ( 
.A1(n_861),
.A2(n_270),
.B1(n_291),
.B2(n_286),
.C(n_320),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_830),
.B(n_783),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_859),
.A2(n_286),
.B1(n_249),
.B2(n_216),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_903),
.B(n_813),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_888),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_826),
.B(n_750),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_906),
.A2(n_740),
.B(n_786),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_832),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_827),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_816),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_865),
.B(n_213),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_902),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_854),
.B(n_213),
.Y(n_938)
);

OR2x6_ASAP7_75t_L g939 ( 
.A(n_871),
.B(n_740),
.Y(n_939)
);

OAI22xp33_ASAP7_75t_L g940 ( 
.A1(n_820),
.A2(n_792),
.B1(n_810),
.B2(n_215),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_832),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_841),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_837),
.A2(n_215),
.B1(n_301),
.B2(n_290),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_839),
.B(n_792),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_908),
.A2(n_774),
.B1(n_779),
.B2(n_773),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_879),
.B(n_250),
.Y(n_946)
);

NAND2xp33_ASAP7_75t_SL g947 ( 
.A(n_860),
.B(n_773),
.Y(n_947)
);

AO31x2_ASAP7_75t_L g948 ( 
.A1(n_914),
.A2(n_793),
.A3(n_807),
.B(n_767),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_835),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_841),
.Y(n_950)
);

BUFx4f_ASAP7_75t_L g951 ( 
.A(n_889),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_860),
.A2(n_216),
.B1(n_250),
.B2(n_254),
.Y(n_952)
);

OAI221xp5_ASAP7_75t_L g953 ( 
.A1(n_847),
.A2(n_789),
.B1(n_288),
.B2(n_258),
.C(n_254),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_822),
.B(n_258),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_845),
.B(n_750),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_851),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_906),
.A2(n_786),
.B(n_722),
.Y(n_957)
);

NAND2xp33_ASAP7_75t_L g958 ( 
.A(n_885),
.B(n_768),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_821),
.B(n_262),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_851),
.Y(n_960)
);

NAND2xp33_ASAP7_75t_R g961 ( 
.A(n_814),
.B(n_722),
.Y(n_961)
);

AOI21x1_ASAP7_75t_L g962 ( 
.A1(n_815),
.A2(n_780),
.B(n_770),
.Y(n_962)
);

BUFx12f_ASAP7_75t_L g963 ( 
.A(n_858),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_821),
.B(n_777),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_845),
.B(n_750),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_908),
.A2(n_781),
.B1(n_262),
.B2(n_301),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_885),
.A2(n_873),
.B(n_913),
.C(n_824),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_853),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_880),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_909),
.A2(n_216),
.B1(n_288),
.B2(n_289),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_887),
.A2(n_448),
.B(n_430),
.Y(n_971)
);

INVx5_ASAP7_75t_L g972 ( 
.A(n_900),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_856),
.A2(n_448),
.B(n_430),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_814),
.B(n_777),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_867),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_850),
.B(n_777),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_896),
.B(n_289),
.Y(n_977)
);

AO21x2_ASAP7_75t_L g978 ( 
.A1(n_890),
.A2(n_448),
.B(n_430),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_911),
.Y(n_979)
);

BUFx12f_ASAP7_75t_L g980 ( 
.A(n_880),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_853),
.B(n_290),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_896),
.B(n_462),
.Y(n_982)
);

OR2x6_ASAP7_75t_L g983 ( 
.A(n_871),
.B(n_462),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_838),
.A2(n_319),
.B1(n_462),
.B2(n_469),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_814),
.B(n_74),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_873),
.B(n_319),
.Y(n_986)
);

NAND2x1p5_ASAP7_75t_L g987 ( 
.A(n_840),
.B(n_412),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_838),
.A2(n_429),
.B(n_6),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_852),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_896),
.B(n_469),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_848),
.A2(n_415),
.B(n_412),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_905),
.B(n_469),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_905),
.B(n_875),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_874),
.Y(n_994)
);

AOI221xp5_ASAP7_75t_L g995 ( 
.A1(n_915),
.A2(n_469),
.B1(n_415),
.B2(n_11),
.C(n_14),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_913),
.A2(n_4),
.B(n_8),
.C(n_14),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_907),
.A2(n_469),
.B1(n_415),
.B2(n_16),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_891),
.A2(n_415),
.B(n_469),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_863),
.B(n_469),
.Y(n_999)
);

OAI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_878),
.A2(n_4),
.B1(n_15),
.B2(n_16),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_840),
.Y(n_1001)
);

OAI221xp5_ASAP7_75t_L g1002 ( 
.A1(n_953),
.A2(n_876),
.B1(n_912),
.B2(n_855),
.C(n_852),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_934),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_920),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_921),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_1000),
.A2(n_928),
.B1(n_988),
.B2(n_995),
.Y(n_1006)
);

OR2x6_ASAP7_75t_L g1007 ( 
.A(n_918),
.B(n_893),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_930),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_968),
.B(n_828),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_928),
.A2(n_970),
.B1(n_952),
.B2(n_986),
.Y(n_1010)
);

OAI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_1000),
.A2(n_855),
.B1(n_893),
.B2(n_892),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_927),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_937),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_949),
.Y(n_1014)
);

OAI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_943),
.A2(n_893),
.B1(n_892),
.B2(n_828),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_SL g1016 ( 
.A1(n_922),
.A2(n_900),
.B1(n_862),
.B2(n_840),
.Y(n_1016)
);

AOI21xp33_ASAP7_75t_L g1017 ( 
.A1(n_952),
.A2(n_818),
.B(n_846),
.Y(n_1017)
);

OAI221xp5_ASAP7_75t_L g1018 ( 
.A1(n_997),
.A2(n_910),
.B1(n_869),
.B2(n_864),
.C(n_894),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_SL g1019 ( 
.A1(n_922),
.A2(n_900),
.B1(n_843),
.B2(n_846),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_938),
.B(n_843),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_926),
.A2(n_843),
.B1(n_900),
.B2(n_882),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_944),
.Y(n_1022)
);

AOI21xp33_ASAP7_75t_L g1023 ( 
.A1(n_958),
.A2(n_849),
.B(n_898),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_918),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_972),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_935),
.Y(n_1026)
);

AOI221xp5_ASAP7_75t_L g1027 ( 
.A1(n_996),
.A2(n_874),
.B1(n_849),
.B2(n_899),
.C(n_897),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_931),
.B(n_842),
.Y(n_1028)
);

BUFx10_ASAP7_75t_L g1029 ( 
.A(n_985),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_942),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_997),
.A2(n_900),
.B(n_829),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_950),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_979),
.A2(n_904),
.B1(n_825),
.B2(n_881),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_973),
.A2(n_917),
.B(n_886),
.Y(n_1034)
);

BUFx4f_ASAP7_75t_SL g1035 ( 
.A(n_925),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_940),
.A2(n_819),
.B1(n_825),
.B2(n_872),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_924),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_933),
.Y(n_1038)
);

AOI22x1_ASAP7_75t_L g1039 ( 
.A1(n_954),
.A2(n_904),
.B1(n_916),
.B2(n_872),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_940),
.A2(n_819),
.B1(n_872),
.B2(n_881),
.Y(n_1040)
);

AOI221xp5_ASAP7_75t_L g1041 ( 
.A1(n_996),
.A2(n_881),
.B1(n_890),
.B2(n_817),
.C(n_415),
.Y(n_1041)
);

OAI21xp33_ASAP7_75t_L g1042 ( 
.A1(n_981),
.A2(n_866),
.B(n_917),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_947),
.A2(n_868),
.B1(n_836),
.B2(n_831),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_947),
.A2(n_868),
.B1(n_836),
.B2(n_831),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_951),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_967),
.A2(n_836),
.B1(n_868),
.B2(n_817),
.Y(n_1046)
);

AOI221xp5_ASAP7_75t_L g1047 ( 
.A1(n_967),
.A2(n_966),
.B1(n_958),
.B2(n_923),
.C(n_936),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_SL g1048 ( 
.A1(n_969),
.A2(n_817),
.B1(n_18),
.B2(n_19),
.Y(n_1048)
);

NOR3xp33_ASAP7_75t_L g1049 ( 
.A(n_946),
.B(n_901),
.C(n_895),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_SL g1050 ( 
.A(n_969),
.B(n_817),
.C(n_19),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_993),
.A2(n_833),
.B1(n_844),
.B2(n_834),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_933),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_924),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_SL g1054 ( 
.A1(n_985),
.A2(n_833),
.B1(n_844),
.B2(n_834),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_941),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_941),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_980),
.A2(n_415),
.B1(n_21),
.B2(n_22),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_989),
.Y(n_1058)
);

NAND2x1_ASAP7_75t_L g1059 ( 
.A(n_939),
.B(n_842),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_1013),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_1003),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1024),
.B(n_976),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1024),
.B(n_955),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1024),
.B(n_965),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_1059),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1022),
.B(n_842),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_1012),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1046),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1004),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1005),
.B(n_842),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1034),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_1028),
.B(n_857),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1008),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1034),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1038),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_1043),
.B(n_857),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_1030),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1052),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_1007),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1044),
.B(n_857),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1006),
.A2(n_929),
.B1(n_935),
.B2(n_972),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1044),
.B(n_974),
.Y(n_1082)
);

INVx2_ASAP7_75t_SL g1083 ( 
.A(n_1007),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1055),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1051),
.B(n_1041),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1056),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_1032),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1051),
.B(n_974),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1009),
.B(n_956),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_1007),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_1014),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1042),
.Y(n_1092)
);

INVx4_ASAP7_75t_L g1093 ( 
.A(n_1025),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1054),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_1050),
.B(n_948),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_1036),
.B(n_948),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_1037),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_1036),
.B(n_948),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1040),
.B(n_964),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_1040),
.B(n_948),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1019),
.B(n_964),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1016),
.B(n_918),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1023),
.B(n_978),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_1058),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_1006),
.A2(n_977),
.B1(n_945),
.B2(n_959),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1049),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1105),
.A2(n_1010),
.B1(n_1048),
.B2(n_1047),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1060),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1061),
.B(n_1053),
.Y(n_1109)
);

NAND5xp2_ASAP7_75t_SL g1110 ( 
.A(n_1105),
.B(n_1057),
.C(n_1002),
.D(n_1021),
.E(n_1026),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1060),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1082),
.B(n_1020),
.Y(n_1112)
);

OAI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1081),
.A2(n_1011),
.B1(n_1015),
.B2(n_1018),
.Y(n_1113)
);

AOI31xp33_ASAP7_75t_L g1114 ( 
.A1(n_1081),
.A2(n_1057),
.A3(n_1026),
.B(n_1017),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1082),
.B(n_1031),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1060),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1060),
.Y(n_1117)
);

OA21x2_ASAP7_75t_L g1118 ( 
.A1(n_1071),
.A2(n_1074),
.B(n_1106),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1091),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_1068),
.B(n_1033),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1085),
.A2(n_1029),
.B1(n_984),
.B2(n_1045),
.Y(n_1121)
);

OAI221xp5_ASAP7_75t_SL g1122 ( 
.A1(n_1094),
.A2(n_1027),
.B1(n_971),
.B2(n_992),
.C(n_983),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1082),
.B(n_1063),
.Y(n_1123)
);

INVxp67_ASAP7_75t_L g1124 ( 
.A(n_1091),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1069),
.Y(n_1125)
);

OAI31xp33_ASAP7_75t_L g1126 ( 
.A1(n_1094),
.A2(n_1001),
.A3(n_919),
.B(n_990),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1063),
.B(n_939),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_1104),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1061),
.B(n_1039),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1063),
.B(n_939),
.Y(n_1130)
);

OA21x2_ASAP7_75t_L g1131 ( 
.A1(n_1071),
.A2(n_973),
.B(n_991),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_1072),
.B(n_978),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1069),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_1072),
.B(n_884),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_1067),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1085),
.A2(n_1045),
.B1(n_972),
.B2(n_951),
.Y(n_1136)
);

NAND2xp33_ASAP7_75t_R g1137 ( 
.A(n_1104),
.B(n_1035),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1069),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1064),
.B(n_960),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1064),
.B(n_1025),
.Y(n_1140)
);

NAND2xp33_ASAP7_75t_R g1141 ( 
.A(n_1104),
.B(n_17),
.Y(n_1141)
);

OAI221xp5_ASAP7_75t_L g1142 ( 
.A1(n_1106),
.A2(n_1045),
.B1(n_1025),
.B2(n_983),
.C(n_961),
.Y(n_1142)
);

OAI211xp5_ASAP7_75t_L g1143 ( 
.A1(n_1106),
.A2(n_999),
.B(n_998),
.C(n_972),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1071),
.A2(n_962),
.B(n_957),
.Y(n_1144)
);

NAND3xp33_ASAP7_75t_L g1145 ( 
.A(n_1092),
.B(n_961),
.C(n_982),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1083),
.B(n_983),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1073),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1102),
.A2(n_1029),
.B1(n_963),
.B2(n_987),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1073),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_1067),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1073),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_1077),
.Y(n_1152)
);

AOI221xp5_ASAP7_75t_L g1153 ( 
.A1(n_1092),
.A2(n_998),
.B1(n_994),
.B2(n_975),
.C(n_26),
.Y(n_1153)
);

AO21x1_ASAP7_75t_SL g1154 ( 
.A1(n_1095),
.A2(n_1029),
.B(n_884),
.Y(n_1154)
);

OAI211xp5_ASAP7_75t_SL g1155 ( 
.A1(n_1092),
.A2(n_991),
.B(n_975),
.C(n_25),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1077),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1075),
.Y(n_1157)
);

AOI22x1_ASAP7_75t_L g1158 ( 
.A1(n_1095),
.A2(n_987),
.B1(n_24),
.B2(n_26),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1138),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1118),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1108),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1108),
.B(n_1065),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1156),
.B(n_1087),
.Y(n_1163)
);

INVxp67_ASAP7_75t_L g1164 ( 
.A(n_1152),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1118),
.B(n_1135),
.Y(n_1165)
);

NAND4xp25_ASAP7_75t_L g1166 ( 
.A(n_1107),
.B(n_1095),
.C(n_1085),
.D(n_1089),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1156),
.B(n_1087),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1111),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1111),
.B(n_1065),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1123),
.B(n_1088),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1116),
.Y(n_1171)
);

NAND2xp67_ASAP7_75t_L g1172 ( 
.A(n_1129),
.B(n_1102),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1123),
.B(n_1088),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1116),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1115),
.B(n_1088),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1150),
.B(n_1064),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1118),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1115),
.B(n_1062),
.Y(n_1178)
);

NAND4xp25_ASAP7_75t_SL g1179 ( 
.A(n_1141),
.B(n_1085),
.C(n_1102),
.D(n_1101),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1140),
.B(n_1062),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1117),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1118),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1140),
.B(n_1127),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1119),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1127),
.B(n_1062),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1124),
.B(n_1076),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1130),
.B(n_1080),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1125),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1138),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1130),
.B(n_1080),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1160),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1179),
.A2(n_1110),
.B1(n_1113),
.B2(n_1158),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1188),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1175),
.B(n_1112),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1188),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1186),
.B(n_1128),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1175),
.B(n_1109),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1160),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1161),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1175),
.B(n_1120),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1161),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1162),
.B(n_1065),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1168),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1172),
.B(n_1120),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1168),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1171),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1170),
.B(n_1154),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1171),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1162),
.B(n_1147),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1170),
.B(n_1154),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1174),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1173),
.B(n_1079),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1184),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1160),
.Y(n_1214)
);

OAI22xp33_ASAP7_75t_SL g1215 ( 
.A1(n_1172),
.A2(n_1122),
.B1(n_1158),
.B2(n_1142),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1172),
.B(n_1139),
.Y(n_1216)
);

OR2x2_ASAP7_75t_L g1217 ( 
.A(n_1186),
.B(n_1132),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1179),
.B(n_1136),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1207),
.B(n_1173),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1204),
.B(n_1178),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1193),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1193),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1200),
.B(n_1186),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1216),
.B(n_1178),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1218),
.B(n_1178),
.Y(n_1225)
);

AOI32xp33_ASAP7_75t_L g1226 ( 
.A1(n_1192),
.A2(n_1173),
.A3(n_1190),
.B1(n_1187),
.B2(n_1155),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1196),
.B(n_1184),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1207),
.B(n_1187),
.Y(n_1228)
);

NOR3xp33_ASAP7_75t_L g1229 ( 
.A(n_1215),
.B(n_1166),
.C(n_1114),
.Y(n_1229)
);

INVx1_ASAP7_75t_SL g1230 ( 
.A(n_1213),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1209),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1197),
.B(n_1185),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_1196),
.B(n_1176),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1195),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1210),
.B(n_1190),
.Y(n_1235)
);

AO21x2_ASAP7_75t_L g1236 ( 
.A1(n_1191),
.A2(n_1177),
.B(n_1160),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1202),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1194),
.B(n_1185),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1212),
.B(n_1180),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1209),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_SL g1241 ( 
.A(n_1202),
.B(n_1110),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1199),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1199),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1201),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1201),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1212),
.B(n_1180),
.Y(n_1246)
);

AOI221xp5_ASAP7_75t_L g1247 ( 
.A1(n_1203),
.A2(n_1164),
.B1(n_1153),
.B2(n_1145),
.C(n_1163),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1222),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1219),
.Y(n_1249)
);

OAI21xp33_ASAP7_75t_SL g1250 ( 
.A1(n_1226),
.A2(n_1183),
.B(n_1217),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1222),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1219),
.B(n_1237),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1229),
.A2(n_1164),
.B(n_1165),
.C(n_1143),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1228),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1228),
.B(n_1183),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1225),
.A2(n_1148),
.B1(n_1121),
.B2(n_1083),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1241),
.B(n_1190),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1247),
.A2(n_1167),
.B(n_1163),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_SL g1259 ( 
.A1(n_1230),
.A2(n_1137),
.B(n_1165),
.C(n_1159),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1220),
.A2(n_1167),
.B(n_1202),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1227),
.A2(n_1121),
.B(n_1202),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_1227),
.Y(n_1262)
);

NOR3xp33_ASAP7_75t_L g1263 ( 
.A(n_1234),
.B(n_1177),
.C(n_1191),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1232),
.A2(n_1126),
.B(n_1101),
.C(n_1165),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1224),
.A2(n_1206),
.B(n_1205),
.Y(n_1265)
);

INVxp67_ASAP7_75t_L g1266 ( 
.A(n_1221),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1238),
.B(n_1180),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1233),
.A2(n_1090),
.B1(n_1146),
.B2(n_1079),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1235),
.A2(n_1090),
.B1(n_1079),
.B2(n_1146),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1262),
.B(n_1233),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1252),
.B(n_1231),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1254),
.B(n_1240),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1250),
.B(n_1223),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1249),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1257),
.B(n_1223),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1254),
.B(n_1240),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1256),
.A2(n_1242),
.B1(n_1245),
.B2(n_1244),
.Y(n_1277)
);

OR2x2_ASAP7_75t_L g1278 ( 
.A(n_1249),
.B(n_1243),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1255),
.B(n_1239),
.Y(n_1279)
);

NOR3xp33_ASAP7_75t_SL g1280 ( 
.A(n_1264),
.B(n_1244),
.C(n_1243),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1258),
.B(n_1246),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1248),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1251),
.Y(n_1283)
);

NAND3xp33_ASAP7_75t_L g1284 ( 
.A(n_1253),
.B(n_1245),
.C(n_1198),
.Y(n_1284)
);

OAI321xp33_ASAP7_75t_L g1285 ( 
.A1(n_1261),
.A2(n_1214),
.A3(n_1198),
.B1(n_1191),
.B2(n_1066),
.C(n_1211),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1267),
.B(n_1206),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1264),
.A2(n_1208),
.B(n_1169),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1266),
.B(n_1265),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1263),
.Y(n_1289)
);

OAI21xp33_ASAP7_75t_L g1290 ( 
.A1(n_1260),
.A2(n_1169),
.B(n_1162),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1268),
.B(n_1183),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1263),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1259),
.A2(n_1169),
.B(n_1162),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1274),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1271),
.B(n_1269),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1274),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_R g1297 ( 
.A(n_1288),
.B(n_23),
.Y(n_1297)
);

AOI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1280),
.A2(n_1259),
.B1(n_1169),
.B2(n_1097),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1271),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1278),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1278),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1283),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1282),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1279),
.B(n_1214),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1275),
.B(n_1214),
.Y(n_1305)
);

XNOR2xp5_ASAP7_75t_L g1306 ( 
.A(n_1277),
.B(n_1099),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1277),
.A2(n_1281),
.B1(n_1273),
.B2(n_1288),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1270),
.Y(n_1308)
);

NAND2x1_ASAP7_75t_L g1309 ( 
.A(n_1293),
.B(n_1159),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1287),
.B(n_1097),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1272),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1272),
.B(n_1236),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_R g1313 ( 
.A(n_1289),
.B(n_28),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1292),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1276),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1286),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1284),
.Y(n_1317)
);

INVxp67_ASAP7_75t_L g1318 ( 
.A(n_1291),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1290),
.B(n_1236),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1299),
.B(n_1236),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_SL g1321 ( 
.A(n_1308),
.B(n_1097),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1307),
.A2(n_1285),
.B(n_1182),
.C(n_1096),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_SL g1323 ( 
.A(n_1299),
.B(n_1317),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1311),
.B(n_1295),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1311),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1315),
.B(n_1294),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1296),
.B(n_1181),
.Y(n_1327)
);

NOR2x1_ASAP7_75t_L g1328 ( 
.A(n_1303),
.B(n_1189),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1318),
.B(n_1159),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1300),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1297),
.B(n_1298),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1313),
.B(n_1093),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1300),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_1301),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1314),
.B(n_1133),
.Y(n_1335)
);

OAI211xp5_ASAP7_75t_L g1336 ( 
.A1(n_1313),
.A2(n_1093),
.B(n_1100),
.C(n_1098),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1316),
.B(n_1151),
.Y(n_1337)
);

AND4x1_ASAP7_75t_L g1338 ( 
.A(n_1302),
.B(n_29),
.C(n_30),
.D(n_31),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1303),
.B(n_30),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1309),
.A2(n_1093),
.B1(n_1100),
.B2(n_1096),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1301),
.Y(n_1341)
);

OAI211xp5_ASAP7_75t_SL g1342 ( 
.A1(n_1310),
.A2(n_1096),
.B(n_34),
.C(n_35),
.Y(n_1342)
);

XNOR2x2_ASAP7_75t_L g1343 ( 
.A(n_1306),
.B(n_33),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1304),
.B(n_1305),
.Y(n_1344)
);

OAI21xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1331),
.A2(n_1319),
.B(n_1312),
.Y(n_1345)
);

AOI21xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1331),
.A2(n_33),
.B(n_34),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1334),
.B(n_1149),
.Y(n_1347)
);

OAI21xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1332),
.A2(n_1333),
.B(n_1330),
.Y(n_1348)
);

AOI221x1_ASAP7_75t_L g1349 ( 
.A1(n_1339),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.C(n_39),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1323),
.A2(n_1103),
.B1(n_1157),
.B2(n_1086),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1342),
.A2(n_1157),
.B1(n_1086),
.B2(n_1084),
.Y(n_1351)
);

AOI21xp33_ASAP7_75t_L g1352 ( 
.A1(n_1321),
.A2(n_40),
.B(n_44),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1324),
.A2(n_1084),
.B1(n_1075),
.B2(n_1078),
.Y(n_1353)
);

AO221x1_ASAP7_75t_L g1354 ( 
.A1(n_1340),
.A2(n_1325),
.B1(n_1341),
.B2(n_1343),
.C(n_1336),
.Y(n_1354)
);

AOI221xp5_ASAP7_75t_L g1355 ( 
.A1(n_1322),
.A2(n_1078),
.B1(n_1086),
.B2(n_1084),
.C(n_1070),
.Y(n_1355)
);

AOI221xp5_ASAP7_75t_L g1356 ( 
.A1(n_1326),
.A2(n_1078),
.B1(n_1070),
.B2(n_1074),
.C(n_1071),
.Y(n_1356)
);

AOI211x1_ASAP7_75t_SL g1357 ( 
.A1(n_1341),
.A2(n_45),
.B(n_46),
.C(n_48),
.Y(n_1357)
);

NAND4xp25_ASAP7_75t_SL g1358 ( 
.A(n_1324),
.B(n_1134),
.C(n_1072),
.D(n_1076),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1339),
.A2(n_46),
.B(n_49),
.C(n_50),
.Y(n_1359)
);

AOI211x1_ASAP7_75t_SL g1360 ( 
.A1(n_1329),
.A2(n_1327),
.B(n_1335),
.C(n_1337),
.Y(n_1360)
);

OAI211xp5_ASAP7_75t_L g1361 ( 
.A1(n_1328),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_1361)
);

NOR2x1_ASAP7_75t_L g1362 ( 
.A(n_1344),
.B(n_52),
.Y(n_1362)
);

NOR2x1_ASAP7_75t_L g1363 ( 
.A(n_1320),
.B(n_53),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1338),
.A2(n_1144),
.B(n_1074),
.Y(n_1364)
);

OAI221xp5_ASAP7_75t_SL g1365 ( 
.A1(n_1345),
.A2(n_60),
.B1(n_62),
.B2(n_64),
.C(n_65),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1362),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1363),
.Y(n_1367)
);

NOR2x1_ASAP7_75t_L g1368 ( 
.A(n_1361),
.B(n_67),
.Y(n_1368)
);

AOI21xp33_ASAP7_75t_SL g1369 ( 
.A1(n_1352),
.A2(n_68),
.B(n_70),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1348),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_R g1371 ( 
.A(n_1346),
.B(n_70),
.Y(n_1371)
);

OAI211xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1360),
.A2(n_71),
.B(n_72),
.C(n_80),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1359),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1364),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1357),
.B(n_71),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1349),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1354),
.B(n_72),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1347),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1347),
.Y(n_1379)
);

NAND4xp75_ASAP7_75t_L g1380 ( 
.A(n_1377),
.B(n_1355),
.C(n_1350),
.D(n_1351),
.Y(n_1380)
);

NAND3xp33_ASAP7_75t_L g1381 ( 
.A(n_1370),
.B(n_1356),
.C(n_1353),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1366),
.B(n_1367),
.Y(n_1382)
);

NOR2xp67_ASAP7_75t_L g1383 ( 
.A(n_1366),
.B(n_1378),
.Y(n_1383)
);

INVxp67_ASAP7_75t_SL g1384 ( 
.A(n_1368),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1371),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1372),
.A2(n_1358),
.B(n_1131),
.Y(n_1386)
);

NOR3xp33_ASAP7_75t_SL g1387 ( 
.A(n_1365),
.B(n_95),
.C(n_97),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1371),
.Y(n_1388)
);

AOI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1374),
.A2(n_932),
.B1(n_429),
.B2(n_111),
.Y(n_1389)
);

NAND4xp75_ASAP7_75t_L g1390 ( 
.A(n_1376),
.B(n_103),
.C(n_107),
.D(n_112),
.Y(n_1390)
);

NOR2x1p5_ASAP7_75t_L g1391 ( 
.A(n_1373),
.B(n_115),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1379),
.Y(n_1392)
);

O2A1O1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1384),
.A2(n_1375),
.B(n_1369),
.C(n_1374),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1392),
.Y(n_1394)
);

NAND3xp33_ASAP7_75t_L g1395 ( 
.A(n_1383),
.B(n_1385),
.C(n_1388),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1382),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1381),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1380),
.A2(n_429),
.B1(n_135),
.B2(n_136),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1395),
.A2(n_1391),
.B1(n_1387),
.B2(n_1390),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1396),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1394),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_SL g1402 ( 
.A1(n_1399),
.A2(n_1393),
.B(n_1398),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1400),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1401),
.B(n_1397),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1403),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_SL g1406 ( 
.A1(n_1405),
.A2(n_1402),
.B1(n_1404),
.B2(n_1389),
.Y(n_1406)
);

XNOR2xp5_ASAP7_75t_L g1407 ( 
.A(n_1406),
.B(n_1386),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1407),
.A2(n_144),
.B(n_146),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1408),
.Y(n_1409)
);

OAI221xp5_ASAP7_75t_L g1410 ( 
.A1(n_1409),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.C(n_168),
.Y(n_1410)
);

AOI211xp5_ASAP7_75t_L g1411 ( 
.A1(n_1410),
.A2(n_177),
.B(n_178),
.C(n_179),
.Y(n_1411)
);


endmodule