module fake_aes_11740_n_40 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
wire n_39;
OAI22xp5_ASAP7_75t_SL g12 ( .A1(n_0), .A2(n_7), .B1(n_6), .B2(n_2), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_1), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_11), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_7), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_10), .B(n_11), .Y(n_17) );
AOI22xp33_ASAP7_75t_L g18 ( .A1(n_14), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_16), .B(n_3), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_16), .B(n_3), .Y(n_20) );
NAND2xp5_ASAP7_75t_SL g21 ( .A(n_16), .B(n_4), .Y(n_21) );
OAI21xp5_ASAP7_75t_L g22 ( .A1(n_19), .A2(n_14), .B(n_17), .Y(n_22) );
A2O1A1Ixp33_ASAP7_75t_L g23 ( .A1(n_19), .A2(n_13), .B(n_15), .C(n_12), .Y(n_23) );
BUFx2_ASAP7_75t_L g24 ( .A(n_19), .Y(n_24) );
AOI221xp5_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_12), .B1(n_19), .B2(n_20), .C(n_18), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
OAI21xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_22), .B(n_24), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_19), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
OAI22xp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_18), .B1(n_20), .B2(n_21), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
OAI322xp33_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_13), .A3(n_20), .B1(n_6), .B2(n_8), .C1(n_9), .C2(n_5), .Y(n_32) );
AOI22xp5_ASAP7_75t_L g33 ( .A1(n_29), .A2(n_27), .B1(n_20), .B2(n_13), .Y(n_33) );
INVx2_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
AOI221xp5_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_27), .B1(n_13), .B2(n_8), .C(n_9), .Y(n_35) );
INVx1_ASAP7_75t_SL g36 ( .A(n_33), .Y(n_36) );
INVx3_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
OAI21xp5_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_13), .B(n_4), .Y(n_38) );
AOI21xp33_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_36), .B(n_13), .Y(n_39) );
AOI22xp33_ASAP7_75t_L g40 ( .A1(n_39), .A2(n_5), .B1(n_37), .B2(n_36), .Y(n_40) );
endmodule