module fake_jpeg_17235_n_344 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_48),
.Y(n_53)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_42),
.B(n_24),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_18),
.B(n_0),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_31),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_33),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_21),
.B1(n_24),
.B2(n_31),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_66),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_27),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_27),
.B(n_28),
.C(n_19),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_72),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_93),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_47),
.B1(n_46),
.B2(n_40),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_77),
.A2(n_81),
.B1(n_91),
.B2(n_94),
.Y(n_118)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_43),
.B1(n_26),
.B2(n_29),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_87),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_31),
.B(n_30),
.C(n_21),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_96),
.B(n_0),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_41),
.C(n_32),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_63),
.C(n_50),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_30),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_30),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_104),
.Y(n_113)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_53),
.A2(n_26),
.B1(n_33),
.B2(n_24),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_92),
.A2(n_100),
.B1(n_106),
.B2(n_110),
.Y(n_123)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_26),
.B1(n_21),
.B2(n_33),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_66),
.A2(n_19),
.B1(n_28),
.B2(n_22),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_97),
.B(n_55),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_67),
.A2(n_23),
.B1(n_22),
.B2(n_19),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_58),
.B1(n_49),
.B2(n_50),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_65),
.A2(n_71),
.B1(n_68),
.B2(n_57),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_111),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_66),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_102),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_0),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_35),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_41),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_52),
.A2(n_23),
.B1(n_28),
.B2(n_34),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_60),
.B(n_17),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_17),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_17),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_55),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_57),
.A2(n_16),
.B1(n_32),
.B2(n_35),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_114),
.A2(n_130),
.B1(n_79),
.B2(n_78),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_16),
.B(n_32),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_127),
.B1(n_103),
.B2(n_101),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_116),
.A2(n_1),
.B(n_2),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_100),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_132),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_128),
.C(n_74),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_126),
.A2(n_135),
.B1(n_86),
.B2(n_76),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_50),
.B1(n_63),
.B2(n_58),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_89),
.C(n_87),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_73),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g131 ( 
.A1(n_88),
.A2(n_63),
.B1(n_16),
.B2(n_72),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_75),
.B1(n_35),
.B2(n_5),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_75),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_136),
.B(n_132),
.CI(n_140),
.CON(n_174),
.SN(n_174)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_99),
.A2(n_55),
.B1(n_35),
.B2(n_3),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_137),
.A2(n_92),
.B1(n_102),
.B2(n_86),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_95),
.B(n_15),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_138),
.B(n_15),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_140),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_97),
.B(n_55),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_1),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_136),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_121),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_150),
.Y(n_178)
);

AO21x1_ASAP7_75t_L g208 ( 
.A1(n_143),
.A2(n_145),
.B(n_142),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_172),
.B1(n_127),
.B2(n_134),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_103),
.B1(n_95),
.B2(n_83),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_147),
.A2(n_153),
.B1(n_154),
.B2(n_166),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_105),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_156),
.C(n_171),
.Y(n_183)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_109),
.B1(n_108),
.B2(n_107),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_111),
.B1(n_93),
.B2(n_90),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_158),
.Y(n_197)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_115),
.A2(n_82),
.B1(n_84),
.B2(n_80),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_161),
.Y(n_203)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_162),
.B(n_164),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_167),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_134),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_123),
.A2(n_78),
.B1(n_84),
.B2(n_3),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_112),
.B(n_84),
.C(n_2),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_113),
.B(n_138),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_1),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_133),
.Y(n_189)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_35),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_120),
.B(n_35),
.C(n_4),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_3),
.C(n_5),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_174),
.B(n_122),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_113),
.A3(n_112),
.B1(n_129),
.B2(n_141),
.C1(n_139),
.C2(n_116),
.Y(n_175)
);

A2O1A1O1Ixp25_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_184),
.B(n_206),
.C(n_159),
.D(n_171),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_155),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_176),
.B(n_190),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_179),
.A2(n_182),
.B(n_188),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_199),
.B1(n_201),
.B2(n_145),
.Y(n_212)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_120),
.Y(n_184)
);

AO22x1_ASAP7_75t_SL g186 ( 
.A1(n_152),
.A2(n_118),
.B1(n_137),
.B2(n_117),
.Y(n_186)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_136),
.C(n_137),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_205),
.C(n_193),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_135),
.B(n_122),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_189),
.B(n_180),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_149),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_202),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_151),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_194),
.B(n_195),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_125),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_166),
.A2(n_114),
.B1(n_4),
.B2(n_5),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_154),
.A2(n_114),
.B1(n_5),
.B2(n_6),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_200),
.A2(n_160),
.B1(n_157),
.B2(n_146),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_153),
.A2(n_163),
.B1(n_146),
.B2(n_173),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_161),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_7),
.Y(n_221)
);

XNOR2x2_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_6),
.Y(n_205)
);

AO21x1_ASAP7_75t_L g219 ( 
.A1(n_205),
.A2(n_208),
.B(n_14),
.Y(n_219)
);

AND2x6_ASAP7_75t_L g206 ( 
.A(n_148),
.B(n_7),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_211),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_212),
.A2(n_213),
.B1(n_232),
.B2(n_180),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_144),
.B1(n_152),
.B2(n_169),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_196),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_214),
.B(n_215),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_185),
.A2(n_158),
.B1(n_170),
.B2(n_10),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_218),
.A2(n_233),
.B1(n_234),
.B2(n_182),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_219),
.B(n_227),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_220),
.A2(n_229),
.B1(n_202),
.B2(n_207),
.Y(n_249)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_7),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_225),
.C(n_230),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_226),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_8),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_228),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_178),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_10),
.C(n_13),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_177),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_231),
.B(n_204),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_13),
.B1(n_14),
.B2(n_194),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_186),
.A2(n_13),
.B1(n_14),
.B2(n_208),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_186),
.A2(n_14),
.B1(n_208),
.B2(n_198),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_191),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_187),
.B(n_198),
.C(n_189),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_188),
.C(n_192),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_240),
.A2(n_255),
.B1(n_259),
.B2(n_258),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_243),
.B(n_249),
.Y(n_275)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_244),
.C(n_250),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_217),
.A2(n_206),
.B1(n_191),
.B2(n_195),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_247),
.A2(n_252),
.B1(n_255),
.B2(n_210),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_209),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_253),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_192),
.C(n_176),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_216),
.C(n_211),
.Y(n_269)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_217),
.A2(n_230),
.B1(n_236),
.B2(n_223),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_177),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_235),
.A2(n_179),
.B1(n_200),
.B2(n_177),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_233),
.Y(n_258)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_234),
.B(n_220),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_218),
.B(n_231),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_237),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_239),
.B(n_249),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_224),
.Y(n_261)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_261),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_245),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_270),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_265),
.B(n_282),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_260),
.B(n_257),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_216),
.Y(n_267)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_271),
.C(n_276),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_262),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_238),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_278),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_244),
.C(n_254),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_252),
.C(n_261),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_260),
.C(n_242),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_239),
.B(n_262),
.Y(n_281)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_272),
.B(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_285),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_274),
.A2(n_243),
.B1(n_247),
.B2(n_257),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_286),
.A2(n_297),
.B1(n_280),
.B2(n_283),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_287),
.A2(n_279),
.B(n_274),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g292 ( 
.A(n_267),
.B(n_265),
.CI(n_277),
.CON(n_292),
.SN(n_292)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_270),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_298),
.C(n_299),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_SL g297 ( 
.A1(n_282),
.A2(n_241),
.B(n_281),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_276),
.C(n_269),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_269),
.C(n_264),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_275),
.B(n_283),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_268),
.Y(n_313)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_301),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_268),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_307),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_289),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_305),
.B(n_308),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_284),
.B(n_272),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_306),
.B(n_296),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_292),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_275),
.C(n_264),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_263),
.C(n_266),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_290),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_294),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_287),
.Y(n_323)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_315),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_302),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_317),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_319),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_324),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_312),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_309),
.A2(n_295),
.B1(n_290),
.B2(n_300),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_292),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_288),
.C(n_298),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_330),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_310),
.C(n_311),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_331),
.A2(n_319),
.B(n_322),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_310),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_332),
.A2(n_320),
.B(n_325),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_336),
.C(n_337),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_329),
.A2(n_326),
.B(n_331),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_327),
.A2(n_316),
.B1(n_304),
.B2(n_318),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_333),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_339),
.B(n_335),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_340),
.C(n_333),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_318),
.Y(n_343)
);

BUFx24_ASAP7_75t_SL g344 ( 
.A(n_343),
.Y(n_344)
);


endmodule