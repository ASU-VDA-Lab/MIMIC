module fake_aes_5398_n_517 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_517);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_517;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_141;
wire n_119;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_493;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx3_ASAP7_75t_L g76 ( .A(n_59), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_75), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_73), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_31), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_58), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_57), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_22), .Y(n_82) );
INVxp67_ASAP7_75t_L g83 ( .A(n_45), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_29), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_27), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_5), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_68), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_36), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_72), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_0), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_19), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_2), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_24), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_33), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_28), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_21), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_0), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_2), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_53), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_39), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_11), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_54), .Y(n_102) );
INVxp33_ASAP7_75t_SL g103 ( .A(n_56), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_18), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_41), .Y(n_105) );
INVxp33_ASAP7_75t_SL g106 ( .A(n_1), .Y(n_106) );
BUFx5_ASAP7_75t_L g107 ( .A(n_4), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_60), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_23), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_42), .Y(n_110) );
AND2x4_ASAP7_75t_L g111 ( .A(n_98), .B(n_1), .Y(n_111) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_81), .A2(n_38), .B(n_71), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_107), .Y(n_113) );
AND3x1_ASAP7_75t_L g114 ( .A(n_98), .B(n_3), .C(n_4), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_76), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_107), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_107), .Y(n_117) );
OAI21x1_ASAP7_75t_L g118 ( .A1(n_102), .A2(n_37), .B(n_70), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_107), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_107), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_107), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_86), .B(n_3), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_107), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_107), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_81), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_82), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_102), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_76), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_85), .Y(n_129) );
BUFx3_ASAP7_75t_L g130 ( .A(n_85), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_108), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_108), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_77), .Y(n_133) );
BUFx3_ASAP7_75t_L g134 ( .A(n_115), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_120), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_118), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_120), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_118), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_126), .B(n_110), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_120), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_111), .B(n_101), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_118), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_111), .B(n_101), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_111), .Y(n_144) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_126), .A2(n_106), .B1(n_103), .B2(n_92), .Y(n_145) );
AND2x2_ASAP7_75t_SL g146 ( .A(n_111), .B(n_93), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_125), .B(n_83), .Y(n_147) );
CKINVDCx14_ASAP7_75t_R g148 ( .A(n_111), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_125), .B(n_86), .Y(n_149) );
INVx4_ASAP7_75t_L g150 ( .A(n_120), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_131), .B(n_97), .Y(n_151) );
AND2x6_ASAP7_75t_L g152 ( .A(n_130), .B(n_94), .Y(n_152) );
INVx4_ASAP7_75t_L g153 ( .A(n_120), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_131), .B(n_109), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_128), .Y(n_155) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_130), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_133), .B(n_103), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_115), .Y(n_158) );
INVx5_ASAP7_75t_L g159 ( .A(n_150), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_136), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_144), .Y(n_161) );
INVxp67_ASAP7_75t_SL g162 ( .A(n_156), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_136), .Y(n_163) );
AO22x1_ASAP7_75t_L g164 ( .A1(n_141), .A2(n_106), .B1(n_88), .B2(n_84), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_134), .Y(n_165) );
OR2x4_ASAP7_75t_L g166 ( .A(n_157), .B(n_122), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_151), .B(n_114), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_146), .B(n_87), .Y(n_168) );
NOR2xp33_ASAP7_75t_R g169 ( .A(n_148), .B(n_89), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_144), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_144), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_154), .B(n_130), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_134), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_146), .B(n_87), .Y(n_174) );
NOR2x1p5_ASAP7_75t_L g175 ( .A(n_139), .B(n_122), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_151), .B(n_130), .Y(n_176) );
INVx2_ASAP7_75t_SL g177 ( .A(n_146), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_144), .Y(n_178) );
NOR2x1p5_ASAP7_75t_L g179 ( .A(n_139), .B(n_91), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_149), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_136), .Y(n_181) );
NAND2x1p5_ASAP7_75t_L g182 ( .A(n_149), .B(n_114), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_134), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_141), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_145), .A2(n_105), .B1(n_133), .B2(n_129), .Y(n_185) );
BUFx2_ASAP7_75t_L g186 ( .A(n_152), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_151), .B(n_133), .Y(n_187) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_151), .Y(n_188) );
INVx4_ASAP7_75t_L g189 ( .A(n_150), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_149), .B(n_133), .Y(n_190) );
BUFx4f_ASAP7_75t_L g191 ( .A(n_152), .Y(n_191) );
NAND3xp33_ASAP7_75t_L g192 ( .A(n_164), .B(n_147), .C(n_153), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_161), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_166), .B(n_141), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_189), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_161), .Y(n_196) );
NOR2xp67_ASAP7_75t_L g197 ( .A(n_167), .B(n_141), .Y(n_197) );
BUFx2_ASAP7_75t_L g198 ( .A(n_189), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_166), .B(n_149), .Y(n_199) );
BUFx6f_ASAP7_75t_SL g200 ( .A(n_167), .Y(n_200) );
INVx2_ASAP7_75t_SL g201 ( .A(n_159), .Y(n_201) );
CKINVDCx16_ASAP7_75t_R g202 ( .A(n_169), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_175), .B(n_143), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_170), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_180), .A2(n_143), .B(n_133), .C(n_129), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_159), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_189), .Y(n_207) );
BUFx2_ASAP7_75t_L g208 ( .A(n_180), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_161), .Y(n_209) );
NOR2xp67_ASAP7_75t_L g210 ( .A(n_170), .B(n_143), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_159), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_185), .B(n_143), .Y(n_212) );
OAI21x1_ASAP7_75t_L g213 ( .A1(n_165), .A2(n_112), .B(n_155), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_177), .A2(n_152), .B1(n_90), .B2(n_153), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_177), .A2(n_152), .B1(n_153), .B2(n_150), .Y(n_215) );
INVx2_ASAP7_75t_SL g216 ( .A(n_159), .Y(n_216) );
INVx6_ASAP7_75t_L g217 ( .A(n_159), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_166), .B(n_152), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_171), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_171), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_160), .Y(n_221) );
OAI21xp33_ASAP7_75t_L g222 ( .A1(n_167), .A2(n_135), .B(n_137), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_191), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_203), .A2(n_168), .B1(n_174), .B2(n_179), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_221), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_212), .A2(n_190), .B1(n_162), .B2(n_176), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_220), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_203), .B(n_188), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_220), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_204), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_202), .Y(n_231) );
NAND3xp33_ASAP7_75t_L g232 ( .A(n_192), .B(n_164), .C(n_172), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_197), .B(n_182), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_212), .B(n_182), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_194), .B(n_184), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_204), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_200), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_210), .A2(n_178), .B(n_187), .C(n_184), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_219), .Y(n_239) );
NOR2xp67_ASAP7_75t_L g240 ( .A(n_214), .B(n_5), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_203), .B(n_179), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_219), .Y(n_242) );
OAI221xp5_ASAP7_75t_L g243 ( .A1(n_199), .A2(n_182), .B1(n_178), .B2(n_191), .C(n_186), .Y(n_243) );
OAI21x1_ASAP7_75t_SL g244 ( .A1(n_201), .A2(n_206), .B(n_216), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_193), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_221), .Y(n_246) );
AOI22xp33_ASAP7_75t_SL g247 ( .A1(n_200), .A2(n_186), .B1(n_191), .B2(n_136), .Y(n_247) );
OR2x6_ASAP7_75t_L g248 ( .A(n_195), .B(n_160), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_195), .B(n_129), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_234), .B(n_198), .Y(n_250) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_227), .Y(n_251) );
OAI211xp5_ASAP7_75t_L g252 ( .A1(n_224), .A2(n_222), .B(n_205), .C(n_218), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_226), .A2(n_200), .B1(n_210), .B2(n_208), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_240), .A2(n_208), .B1(n_198), .B2(n_202), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_234), .A2(n_207), .B1(n_209), .B2(n_193), .Y(n_255) );
NOR2xp67_ASAP7_75t_L g256 ( .A(n_227), .B(n_201), .Y(n_256) );
OAI22xp33_ASAP7_75t_L g257 ( .A1(n_243), .A2(n_207), .B1(n_206), .B2(n_216), .Y(n_257) );
OAI221xp5_ASAP7_75t_L g258 ( .A1(n_241), .A2(n_132), .B1(n_215), .B2(n_209), .C(n_196), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_228), .A2(n_207), .B1(n_196), .B2(n_152), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_248), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_229), .Y(n_261) );
OR2x2_ASAP7_75t_L g262 ( .A(n_236), .B(n_211), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_233), .A2(n_152), .B1(n_211), .B2(n_217), .Y(n_263) );
AOI22xp33_ASAP7_75t_SL g264 ( .A1(n_233), .A2(n_217), .B1(n_138), .B2(n_136), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g265 ( .A1(n_232), .A2(n_213), .B(n_165), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_244), .Y(n_266) );
OR2x6_ASAP7_75t_L g267 ( .A(n_248), .B(n_217), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_248), .Y(n_268) );
BUFx12f_ASAP7_75t_L g269 ( .A(n_231), .Y(n_269) );
NAND3xp33_ASAP7_75t_L g270 ( .A(n_238), .B(n_128), .C(n_136), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_254), .A2(n_235), .B1(n_230), .B2(n_237), .Y(n_271) );
OAI211xp5_ASAP7_75t_SL g272 ( .A1(n_253), .A2(n_100), .B(n_79), .C(n_80), .Y(n_272) );
AO21x2_ASAP7_75t_L g273 ( .A1(n_265), .A2(n_213), .B(n_244), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_253), .A2(n_239), .B1(n_242), .B2(n_236), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_266), .A2(n_242), .B(n_239), .C(n_229), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_260), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_251), .A2(n_230), .B1(n_248), .B2(n_247), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_250), .B(n_245), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_266), .B(n_245), .Y(n_279) );
AOI211xp5_ASAP7_75t_L g280 ( .A1(n_257), .A2(n_231), .B(n_95), .C(n_78), .Y(n_280) );
OAI211xp5_ASAP7_75t_L g281 ( .A1(n_252), .A2(n_256), .B(n_255), .C(n_260), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_268), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_250), .B(n_249), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_268), .B(n_249), .Y(n_284) );
OAI22xp33_ASAP7_75t_L g285 ( .A1(n_267), .A2(n_217), .B1(n_99), .B2(n_109), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_261), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_262), .Y(n_287) );
NAND3xp33_ASAP7_75t_SL g288 ( .A(n_262), .B(n_91), .C(n_99), .Y(n_288) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_264), .A2(n_246), .B1(n_225), .B2(n_160), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_258), .A2(n_246), .B1(n_225), .B2(n_160), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_256), .B(n_132), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_272), .A2(n_268), .B1(n_267), .B2(n_269), .Y(n_292) );
AND2x2_ASAP7_75t_SL g293 ( .A(n_276), .B(n_225), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_286), .B(n_267), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_278), .B(n_265), .Y(n_295) );
OAI21xp5_ASAP7_75t_L g296 ( .A1(n_288), .A2(n_270), .B(n_259), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_278), .B(n_267), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_279), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_276), .B(n_267), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_283), .B(n_112), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_283), .B(n_112), .Y(n_301) );
OAI31xp33_ASAP7_75t_L g302 ( .A1(n_281), .A2(n_270), .A3(n_96), .B(n_104), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_273), .Y(n_303) );
AND2x4_ASAP7_75t_SL g304 ( .A(n_279), .B(n_225), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_273), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_282), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_273), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_279), .B(n_269), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_275), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_275), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_287), .B(n_132), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_284), .B(n_225), .Y(n_313) );
AOI21xp5_ASAP7_75t_SL g314 ( .A1(n_277), .A2(n_246), .B(n_221), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_284), .B(n_246), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_274), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_284), .B(n_112), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_291), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g319 ( .A1(n_271), .A2(n_263), .B1(n_127), .B2(n_112), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_289), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_290), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_295), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_295), .B(n_128), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_298), .B(n_128), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_297), .B(n_280), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_294), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_294), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_297), .A2(n_285), .B1(n_127), .B2(n_128), .Y(n_328) );
OAI21xp5_ASAP7_75t_SL g329 ( .A1(n_309), .A2(n_127), .B(n_128), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_306), .Y(n_330) );
OAI21xp33_ASAP7_75t_L g331 ( .A1(n_316), .A2(n_115), .B(n_128), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_306), .B(n_6), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_304), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_313), .B(n_246), .Y(n_334) );
OAI31xp33_ASAP7_75t_L g335 ( .A1(n_302), .A2(n_115), .A3(n_119), .B(n_116), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_313), .B(n_62), .Y(n_336) );
OAI21xp5_ASAP7_75t_L g337 ( .A1(n_296), .A2(n_113), .B(n_117), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_307), .B(n_6), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_307), .B(n_7), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_310), .B(n_7), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_310), .B(n_8), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_318), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_318), .B(n_8), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_300), .B(n_9), .Y(n_344) );
INVxp67_ASAP7_75t_SL g345 ( .A(n_299), .Y(n_345) );
INVx3_ASAP7_75t_SL g346 ( .A(n_304), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_299), .B(n_9), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_303), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_303), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_311), .B(n_10), .Y(n_350) );
NAND2x1p5_ASAP7_75t_L g351 ( .A(n_293), .B(n_221), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_312), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_305), .Y(n_353) );
INVx3_ASAP7_75t_L g354 ( .A(n_304), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_311), .B(n_10), .Y(n_355) );
NAND3x1_ASAP7_75t_SL g356 ( .A(n_300), .B(n_11), .C(n_12), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_301), .B(n_12), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_305), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_305), .B(n_13), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_292), .A2(n_121), .B1(n_116), .B2(n_124), .C(n_119), .Y(n_360) );
OAI21xp5_ASAP7_75t_L g361 ( .A1(n_319), .A2(n_113), .B(n_117), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_308), .B(n_13), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_312), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_308), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_317), .B(n_14), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_322), .B(n_301), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_322), .B(n_315), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_330), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_345), .B(n_293), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_330), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_326), .B(n_293), .Y(n_371) );
NAND3xp33_ASAP7_75t_L g372 ( .A(n_329), .B(n_317), .C(n_319), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_342), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_323), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_323), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_346), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_327), .B(n_320), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_359), .B(n_315), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_347), .B(n_315), .Y(n_379) );
OAI211xp5_ASAP7_75t_SL g380 ( .A1(n_347), .A2(n_314), .B(n_121), .C(n_124), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_359), .B(n_320), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_325), .B(n_14), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_338), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_354), .B(n_315), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_338), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_362), .B(n_313), .Y(n_386) );
INVx3_ASAP7_75t_SL g387 ( .A(n_346), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_362), .B(n_313), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_354), .B(n_320), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_352), .B(n_314), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_363), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_343), .B(n_15), .Y(n_392) );
NAND3xp33_ASAP7_75t_SL g393 ( .A(n_335), .B(n_321), .C(n_15), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_353), .B(n_321), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_333), .B(n_123), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_353), .B(n_123), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_365), .B(n_123), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_332), .Y(n_398) );
AOI32xp33_ASAP7_75t_L g399 ( .A1(n_332), .A2(n_117), .A3(n_113), .B1(n_155), .B2(n_223), .Y(n_399) );
INVx1_ASAP7_75t_SL g400 ( .A(n_339), .Y(n_400) );
NOR3xp33_ASAP7_75t_SL g401 ( .A(n_344), .B(n_16), .C(n_17), .Y(n_401) );
INVxp67_ASAP7_75t_L g402 ( .A(n_324), .Y(n_402) );
INVx1_ASAP7_75t_SL g403 ( .A(n_339), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_340), .Y(n_404) );
OAI21xp33_ASAP7_75t_SL g405 ( .A1(n_365), .A2(n_223), .B(n_25), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_340), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_354), .B(n_20), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_357), .B(n_26), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_358), .B(n_142), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_358), .B(n_30), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_334), .B(n_32), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_364), .B(n_142), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_334), .B(n_34), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_383), .B(n_341), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_373), .Y(n_415) );
NOR2xp33_ASAP7_75t_SL g416 ( .A(n_387), .B(n_331), .Y(n_416) );
AOI211xp5_ASAP7_75t_L g417 ( .A1(n_405), .A2(n_355), .B(n_350), .C(n_341), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_391), .B(n_349), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_382), .A2(n_355), .B1(n_350), .B2(n_324), .Y(n_419) );
INVx2_ASAP7_75t_SL g420 ( .A(n_376), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_400), .B(n_324), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_380), .A2(n_336), .B(n_351), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_392), .A2(n_360), .B1(n_328), .B2(n_348), .C(n_349), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_368), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_375), .Y(n_425) );
AOI32xp33_ASAP7_75t_L g426 ( .A1(n_403), .A2(n_336), .A3(n_356), .B1(n_334), .B2(n_351), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_376), .B(n_336), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_366), .B(n_351), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_370), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_390), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_384), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_393), .A2(n_337), .B1(n_356), .B2(n_361), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_402), .B(n_221), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_366), .B(n_35), .Y(n_434) );
NAND3xp33_ASAP7_75t_L g435 ( .A(n_402), .B(n_138), .C(n_142), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_367), .Y(n_436) );
OR3x2_ASAP7_75t_L g437 ( .A(n_379), .B(n_40), .C(n_43), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_386), .B(n_44), .Y(n_438) );
NOR3xp33_ASAP7_75t_L g439 ( .A(n_393), .B(n_183), .C(n_173), .Y(n_439) );
A2O1A1Ixp33_ASAP7_75t_L g440 ( .A1(n_401), .A2(n_142), .B(n_138), .C(n_160), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_388), .B(n_46), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_385), .B(n_47), .Y(n_442) );
BUFx3_ASAP7_75t_L g443 ( .A(n_384), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_374), .A2(n_138), .B1(n_142), .B2(n_181), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_377), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_377), .B(n_138), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_372), .B(n_138), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_374), .B(n_48), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_398), .B(n_49), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_404), .B(n_50), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_394), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_394), .B(n_51), .Y(n_452) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_389), .A2(n_152), .B(n_173), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_406), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_381), .Y(n_455) );
INVxp33_ASAP7_75t_L g456 ( .A(n_407), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_381), .B(n_52), .Y(n_457) );
XNOR2x1_ASAP7_75t_L g458 ( .A(n_378), .B(n_55), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_397), .Y(n_459) );
XOR2x2_ASAP7_75t_L g460 ( .A(n_369), .B(n_61), .Y(n_460) );
XNOR2xp5_ASAP7_75t_L g461 ( .A(n_371), .B(n_63), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_408), .A2(n_181), .B1(n_163), .B2(n_183), .Y(n_462) );
XOR2x2_ASAP7_75t_L g463 ( .A(n_411), .B(n_64), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_399), .A2(n_158), .B1(n_181), .B2(n_163), .C(n_69), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_396), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_396), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_409), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_409), .B(n_65), .Y(n_468) );
AOI221x1_ASAP7_75t_SL g469 ( .A1(n_412), .A2(n_66), .B1(n_67), .B2(n_74), .C(n_135), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_410), .A2(n_158), .B(n_140), .C(n_137), .Y(n_470) );
INVx3_ASAP7_75t_L g471 ( .A(n_395), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_413), .B(n_163), .Y(n_472) );
XOR2xp5_ASAP7_75t_L g473 ( .A(n_375), .B(n_140), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_375), .B(n_150), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_373), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_375), .Y(n_476) );
OAI321xp33_ASAP7_75t_L g477 ( .A1(n_402), .A2(n_153), .A3(n_393), .B1(n_390), .B2(n_374), .C(n_380), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_420), .A2(n_473), .B1(n_417), .B2(n_431), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g479 ( .A1(n_477), .A2(n_422), .B(n_440), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_430), .B(n_443), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_456), .A2(n_427), .B1(n_425), .B2(n_426), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_459), .B(n_430), .Y(n_482) );
NOR3xp33_ASAP7_75t_L g483 ( .A(n_439), .B(n_464), .C(n_457), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_451), .Y(n_484) );
NAND3xp33_ASAP7_75t_SL g485 ( .A(n_416), .B(n_464), .C(n_432), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_456), .A2(n_427), .B1(n_437), .B2(n_419), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_421), .A2(n_455), .B1(n_436), .B2(n_445), .Y(n_487) );
INVxp33_ASAP7_75t_SL g488 ( .A(n_461), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_447), .A2(n_470), .B(n_416), .C(n_453), .Y(n_489) );
XNOR2x1_ASAP7_75t_L g490 ( .A(n_460), .B(n_463), .Y(n_490) );
OAI22xp33_ASAP7_75t_L g491 ( .A1(n_471), .A2(n_428), .B1(n_476), .B2(n_448), .Y(n_491) );
NAND4xp25_ASAP7_75t_L g492 ( .A(n_469), .B(n_423), .C(n_442), .D(n_449), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_475), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_SL g494 ( .A1(n_433), .A2(n_428), .B(n_434), .C(n_471), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_493), .Y(n_495) );
NOR2x1_ASAP7_75t_L g496 ( .A(n_485), .B(n_458), .Y(n_496) );
OAI221xp5_ASAP7_75t_L g497 ( .A1(n_478), .A2(n_454), .B1(n_415), .B2(n_414), .C(n_424), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_484), .Y(n_498) );
AOI211x1_ASAP7_75t_L g499 ( .A1(n_481), .A2(n_418), .B(n_429), .C(n_457), .Y(n_499) );
OAI311xp33_ASAP7_75t_L g500 ( .A1(n_492), .A2(n_462), .A3(n_450), .B1(n_452), .C1(n_444), .Y(n_500) );
NAND5xp2_ASAP7_75t_L g501 ( .A(n_479), .B(n_470), .C(n_462), .D(n_441), .E(n_438), .Y(n_501) );
OAI22xp33_ASAP7_75t_L g502 ( .A1(n_486), .A2(n_482), .B1(n_491), .B2(n_488), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_480), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_502), .A2(n_494), .B1(n_483), .B2(n_489), .C(n_487), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_503), .Y(n_505) );
NAND5xp2_ASAP7_75t_L g506 ( .A(n_497), .B(n_489), .C(n_490), .D(n_452), .E(n_472), .Y(n_506) );
NOR3xp33_ASAP7_75t_L g507 ( .A(n_502), .B(n_468), .C(n_474), .Y(n_507) );
AND4x1_ASAP7_75t_L g508 ( .A(n_496), .B(n_435), .C(n_468), .D(n_466), .Y(n_508) );
NOR2x1_ASAP7_75t_L g509 ( .A(n_506), .B(n_505), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_507), .Y(n_510) );
OAI321xp33_ASAP7_75t_L g511 ( .A1(n_504), .A2(n_498), .A3(n_500), .B1(n_495), .B2(n_499), .C(n_501), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_509), .A2(n_508), .B1(n_465), .B2(n_467), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_510), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_513), .B(n_511), .Y(n_514) );
BUFx2_ASAP7_75t_L g515 ( .A(n_514), .Y(n_515) );
INVxp67_ASAP7_75t_L g516 ( .A(n_515), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_516), .A2(n_512), .B(n_446), .Y(n_517) );
endmodule