module fake_netlist_5_385_n_1976 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1976);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1976;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1726;
wire n_665;
wire n_1835;
wire n_1584;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

BUFx3_ASAP7_75t_L g204 ( 
.A(n_117),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_148),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_194),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_7),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_50),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_115),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_3),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_88),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_120),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_166),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_132),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_119),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_52),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_91),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_34),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_14),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_122),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_197),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_93),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_165),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_0),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_27),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_201),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_161),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_158),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_125),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_159),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_7),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_109),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_68),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_189),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_112),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_59),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_66),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_21),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_118),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_172),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_196),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_195),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_106),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_20),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_137),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_46),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_199),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_123),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_191),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_72),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_19),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_121),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_176),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_21),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_99),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_186),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_144),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_41),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_58),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_43),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_34),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_111),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_96),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_62),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_0),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_170),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_181),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_75),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_10),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_130),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_31),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_9),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_131),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_26),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_178),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_155),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_2),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_10),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_20),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_60),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_61),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_53),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_152),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_37),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_76),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_84),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_129),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_153),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_16),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_61),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_97),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_70),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_48),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_198),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_173),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_80),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_135),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_67),
.Y(n_299)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_101),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_127),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_36),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_107),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_52),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_98),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_3),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_33),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_14),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_177),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_69),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_59),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_157),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_85),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_182),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_150),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_63),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_203),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_39),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_11),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_77),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_9),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_151),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_33),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_92),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_162),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_39),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_2),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_23),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_42),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_89),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_134),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_54),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_1),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_44),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_12),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_32),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_35),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_11),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_36),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_27),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_100),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_163),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_67),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_1),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g345 ( 
.A(n_17),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_16),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_50),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_17),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_74),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_113),
.Y(n_350)
);

BUFx10_ASAP7_75t_L g351 ( 
.A(n_81),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_87),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_133),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_147),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_8),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_45),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_41),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_108),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_73),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_18),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_180),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_28),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_47),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_164),
.Y(n_364)
);

BUFx10_ASAP7_75t_L g365 ( 
.A(n_174),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_136),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_175),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_102),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_143),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_128),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_35),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_179),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_95),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_56),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_145),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_83),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_40),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_31),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_58),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_60),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_57),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_124),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_22),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_154),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_29),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_18),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_202),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_43),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_139),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_44),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_5),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_5),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_183),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_13),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_187),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_25),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_65),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_19),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_169),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_56),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_24),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_55),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_94),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_25),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_15),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_114),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_290),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_290),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_220),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_290),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_290),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_290),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_290),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_388),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_290),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_290),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_308),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_208),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_262),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_245),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_306),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_262),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_314),
.B(n_4),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_343),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_282),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_282),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_311),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_252),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_311),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_255),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_318),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_317),
.B(n_4),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_268),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_259),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_260),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_261),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_293),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_266),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_318),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_319),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_345),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_319),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_344),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_207),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_373),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_308),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_360),
.Y(n_447)
);

NOR2xp67_ASAP7_75t_L g448 ( 
.A(n_228),
.B(n_6),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_270),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_360),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_216),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_273),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_218),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_279),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_237),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_207),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_280),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_210),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_247),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_210),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_265),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_272),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_246),
.B(n_6),
.Y(n_463)
);

BUFx10_ASAP7_75t_L g464 ( 
.A(n_246),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_379),
.B(n_8),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_325),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_228),
.B(n_12),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_278),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_344),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_219),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_283),
.Y(n_471)
);

NOR2xp67_ASAP7_75t_L g472 ( 
.A(n_228),
.B(n_13),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_285),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_213),
.B(n_15),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_323),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_336),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_377),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_390),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_391),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_291),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_398),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_294),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_345),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_386),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_204),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_404),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_404),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_405),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_204),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_324),
.B(n_22),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_331),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_213),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_287),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_249),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_288),
.B(n_23),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_299),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_250),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_287),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_366),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_251),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_302),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_254),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_366),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_288),
.B(n_26),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_304),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_384),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_384),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_303),
.Y(n_508)
);

BUFx6f_ASAP7_75t_SL g509 ( 
.A(n_227),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_303),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_359),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_264),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_408),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_469),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_408),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_469),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_421),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_494),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_467),
.B(n_205),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_497),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_407),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_411),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_500),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_486),
.Y(n_524)
);

XNOR2x2_ASAP7_75t_L g525 ( 
.A(n_465),
.B(n_337),
.Y(n_525)
);

NAND2xp33_ASAP7_75t_R g526 ( 
.A(n_428),
.B(n_205),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_490),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_412),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_445),
.B(n_222),
.Y(n_529)
);

AND2x6_ASAP7_75t_L g530 ( 
.A(n_490),
.B(n_263),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_417),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_413),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_486),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_502),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_415),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_410),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_410),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_493),
.B(n_206),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_420),
.B(n_227),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_512),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_409),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_428),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_416),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_430),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_430),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_492),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_492),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_433),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_420),
.B(n_206),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_434),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_508),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_508),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_444),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_491),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_510),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_510),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_511),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_498),
.B(n_209),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_435),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_511),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_499),
.B(n_209),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_435),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_503),
.B(n_211),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_436),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_419),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_488),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_419),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_422),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_422),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_425),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_436),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_488),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_446),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_466),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_438),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_447),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_425),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_426),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_426),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_438),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_449),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_506),
.B(n_211),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_427),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_449),
.Y(n_584)
);

NAND2x1_ASAP7_75t_L g585 ( 
.A(n_448),
.B(n_263),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_418),
.B(n_424),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_452),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_427),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_464),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_429),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_429),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_431),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_431),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_439),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_527),
.B(n_485),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_536),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_536),
.Y(n_597)
);

NOR3xp33_ASAP7_75t_L g598 ( 
.A(n_529),
.B(n_432),
.C(n_423),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_553),
.B(n_460),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_527),
.B(n_472),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_553),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_513),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_519),
.B(n_452),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_537),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_537),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_531),
.B(n_489),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_513),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_532),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_531),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_519),
.A2(n_474),
.B1(n_504),
.B2(n_495),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_527),
.B(n_454),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_531),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_589),
.B(n_454),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_573),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_573),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_543),
.B(n_437),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_573),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_576),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_589),
.B(n_275),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_517),
.Y(n_620)
);

BUFx4f_ASAP7_75t_L g621 ( 
.A(n_562),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_576),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_538),
.B(n_460),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_576),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_589),
.B(n_359),
.Y(n_625)
);

INVx4_ASAP7_75t_SL g626 ( 
.A(n_530),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_525),
.A2(n_463),
.B1(n_403),
.B2(n_376),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_538),
.B(n_457),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_558),
.B(n_457),
.Y(n_629)
);

NOR2x1p5_ASAP7_75t_L g630 ( 
.A(n_589),
.B(n_473),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_543),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_587),
.Y(n_632)
);

INVx4_ASAP7_75t_SL g633 ( 
.A(n_530),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_532),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_558),
.B(n_376),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_561),
.B(n_403),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_543),
.B(n_473),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_561),
.B(n_480),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_563),
.B(n_480),
.Y(n_639)
);

OR2x6_ASAP7_75t_L g640 ( 
.A(n_586),
.B(n_441),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_532),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_530),
.B(n_482),
.Y(n_642)
);

OAI21xp33_ASAP7_75t_SL g643 ( 
.A1(n_539),
.A2(n_507),
.B(n_440),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_513),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_L g645 ( 
.A(n_530),
.B(n_263),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_563),
.B(n_263),
.Y(n_646)
);

OAI22xp33_ASAP7_75t_L g647 ( 
.A1(n_582),
.A2(n_362),
.B1(n_346),
.B2(n_414),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_515),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_521),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_518),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_521),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_530),
.B(n_496),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_521),
.Y(n_653)
);

AO22x2_ASAP7_75t_L g654 ( 
.A1(n_525),
.A2(n_235),
.B1(n_244),
.B2(n_214),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_522),
.Y(n_655)
);

AND2x6_ASAP7_75t_L g656 ( 
.A(n_522),
.B(n_263),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_582),
.B(n_358),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_530),
.B(n_522),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_532),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_515),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_530),
.B(n_496),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_549),
.B(n_501),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_528),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_566),
.B(n_451),
.Y(n_664)
);

BUFx4f_ASAP7_75t_L g665 ( 
.A(n_562),
.Y(n_665)
);

AND3x2_ASAP7_75t_L g666 ( 
.A(n_564),
.B(n_328),
.C(n_239),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_528),
.Y(n_667)
);

AND2x6_ASAP7_75t_L g668 ( 
.A(n_528),
.B(n_358),
.Y(n_668)
);

BUFx10_ASAP7_75t_L g669 ( 
.A(n_542),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_535),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_544),
.B(n_501),
.Y(n_671)
);

OR2x6_ASAP7_75t_L g672 ( 
.A(n_566),
.B(n_483),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_585),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_535),
.B(n_505),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_554),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_535),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_545),
.B(n_505),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_532),
.B(n_464),
.Y(n_678)
);

AO22x2_ASAP7_75t_L g679 ( 
.A1(n_585),
.A2(n_253),
.B1(n_256),
.B2(n_248),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_570),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_532),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_570),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_552),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_550),
.B(n_358),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_572),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_547),
.B(n_464),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_572),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_555),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_570),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_559),
.B(n_358),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_555),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_552),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_556),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_556),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_560),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_552),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_570),
.Y(n_697)
);

INVxp67_ASAP7_75t_SL g698 ( 
.A(n_552),
.Y(n_698)
);

NAND3xp33_ASAP7_75t_L g699 ( 
.A(n_526),
.B(n_458),
.C(n_456),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_552),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_552),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_571),
.A2(n_509),
.B1(n_470),
.B2(n_215),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_570),
.Y(n_703)
);

INVx8_ASAP7_75t_L g704 ( 
.A(n_575),
.Y(n_704)
);

OR2x2_ASAP7_75t_SL g705 ( 
.A(n_579),
.B(n_450),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_547),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_L g707 ( 
.A(n_570),
.B(n_358),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_560),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_577),
.Y(n_709)
);

AND2x6_ASAP7_75t_L g710 ( 
.A(n_547),
.B(n_368),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_547),
.B(n_267),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_580),
.B(n_368),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_577),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_579),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_581),
.B(n_368),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_591),
.B(n_509),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_554),
.B(n_453),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_577),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_577),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_591),
.B(n_269),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_591),
.B(n_274),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_583),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_584),
.B(n_455),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_583),
.Y(n_724)
);

NAND2xp33_ASAP7_75t_SL g725 ( 
.A(n_588),
.B(n_281),
.Y(n_725)
);

AO22x2_ASAP7_75t_L g726 ( 
.A1(n_588),
.A2(n_298),
.B1(n_257),
.B2(n_258),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_577),
.B(n_368),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_577),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_590),
.B(n_459),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_590),
.B(n_461),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_546),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_591),
.B(n_277),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_592),
.B(n_462),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_546),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_593),
.Y(n_735)
);

INVxp33_ASAP7_75t_L g736 ( 
.A(n_514),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_514),
.B(n_468),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_546),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_516),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_516),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_603),
.B(n_368),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_685),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_603),
.B(n_551),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_628),
.B(n_369),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_628),
.B(n_369),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_629),
.B(n_551),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_717),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_644),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_629),
.B(n_551),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_644),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_SL g751 ( 
.A(n_619),
.B(n_520),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_638),
.B(n_639),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_627),
.A2(n_338),
.B1(n_340),
.B2(n_327),
.Y(n_753)
);

AND2x6_ASAP7_75t_SL g754 ( 
.A(n_640),
.B(n_471),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_627),
.A2(n_378),
.B1(n_385),
.B2(n_369),
.Y(n_755)
);

BUFx6f_ASAP7_75t_SL g756 ( 
.A(n_669),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_638),
.B(n_557),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_639),
.B(n_369),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_598),
.A2(n_369),
.B1(n_271),
.B2(n_276),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_601),
.Y(n_760)
);

A2O1A1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_610),
.A2(n_611),
.B(n_596),
.C(n_604),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_685),
.Y(n_762)
);

AND2x4_ASAP7_75t_SL g763 ( 
.A(n_669),
.B(n_541),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_602),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_623),
.B(n_212),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_723),
.B(n_523),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_610),
.A2(n_349),
.B1(n_315),
.B2(n_305),
.Y(n_767)
);

BUFx8_ASAP7_75t_L g768 ( 
.A(n_632),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_607),
.Y(n_769)
);

OAI22xp33_ASAP7_75t_L g770 ( 
.A1(n_595),
.A2(n_307),
.B1(n_238),
.B2(n_234),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_597),
.B(n_557),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_706),
.B(n_606),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_704),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_687),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_706),
.B(n_295),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_605),
.B(n_606),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_606),
.B(n_557),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_611),
.B(n_212),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_607),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_674),
.B(n_215),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_706),
.B(n_309),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_614),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_637),
.A2(n_567),
.B(n_565),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_616),
.B(n_310),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_615),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_622),
.B(n_313),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_SL g787 ( 
.A1(n_654),
.A2(n_509),
.B1(n_534),
.B2(n_540),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_688),
.B(n_341),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_729),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_R g790 ( 
.A(n_650),
.B(n_548),
.Y(n_790)
);

INVx8_ASAP7_75t_L g791 ( 
.A(n_704),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_671),
.B(n_345),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_691),
.B(n_354),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_677),
.B(n_475),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_730),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_SL g796 ( 
.A1(n_654),
.A2(n_665),
.B1(n_621),
.B2(n_662),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_693),
.B(n_375),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_662),
.B(n_217),
.Y(n_798)
);

NAND2x1_ASAP7_75t_L g799 ( 
.A(n_734),
.B(n_565),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_600),
.A2(n_286),
.B1(n_284),
.B2(n_289),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_694),
.B(n_382),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_642),
.B(n_387),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_652),
.B(n_406),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_699),
.B(n_217),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_733),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_739),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_739),
.Y(n_807)
);

AND2x6_ASAP7_75t_SL g808 ( 
.A(n_640),
.B(n_672),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_661),
.B(n_292),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_658),
.B(n_673),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_609),
.Y(n_811)
);

A2O1A1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_695),
.A2(n_594),
.B(n_578),
.C(n_569),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_672),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_708),
.B(n_565),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_714),
.B(n_567),
.Y(n_815)
);

NAND2xp33_ASAP7_75t_L g816 ( 
.A(n_613),
.B(n_296),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_722),
.B(n_567),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_736),
.B(n_221),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_724),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_704),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_599),
.B(n_476),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_672),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_650),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_673),
.B(n_297),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_654),
.A2(n_371),
.B1(n_224),
.B2(n_225),
.Y(n_825)
);

OAI221xp5_ASAP7_75t_L g826 ( 
.A1(n_635),
.A2(n_481),
.B1(n_477),
.B2(n_478),
.C(n_479),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_735),
.B(n_568),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_621),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_600),
.B(n_569),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_734),
.B(n_569),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_736),
.B(n_221),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_737),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_643),
.A2(n_350),
.B1(n_301),
.B2(n_320),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_664),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_734),
.B(n_678),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_631),
.B(n_578),
.Y(n_836)
);

INVx4_ASAP7_75t_L g837 ( 
.A(n_634),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_620),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_664),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_664),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_686),
.B(n_578),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_684),
.B(n_223),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_626),
.B(n_322),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_711),
.B(n_594),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_720),
.B(n_594),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_675),
.B(n_219),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_648),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_705),
.B(n_224),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_721),
.B(n_524),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_740),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_609),
.Y(n_851)
);

A2O1A1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_716),
.A2(n_533),
.B(n_353),
.C(n_361),
.Y(n_852)
);

NOR3xp33_ASAP7_75t_L g853 ( 
.A(n_647),
.B(n_725),
.C(n_690),
.Y(n_853)
);

NOR2x1p5_ASAP7_75t_L g854 ( 
.A(n_612),
.B(n_225),
.Y(n_854)
);

OR2x6_ASAP7_75t_L g855 ( 
.A(n_640),
.B(n_574),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_732),
.B(n_330),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_716),
.B(n_342),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_636),
.B(n_352),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_612),
.Y(n_859)
);

AO22x1_ASAP7_75t_L g860 ( 
.A1(n_617),
.A2(n_392),
.B1(n_232),
.B2(n_234),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_684),
.B(n_223),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_636),
.B(n_364),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_617),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_625),
.B(n_367),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_625),
.B(n_618),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_660),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_618),
.B(n_226),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_624),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_SL g869 ( 
.A(n_665),
.B(n_227),
.Y(n_869)
);

INVx4_ASAP7_75t_L g870 ( 
.A(n_634),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_624),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_626),
.B(n_226),
.Y(n_872)
);

INVx8_ASAP7_75t_L g873 ( 
.A(n_710),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_690),
.B(n_231),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_626),
.B(n_231),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_712),
.B(n_715),
.Y(n_876)
);

INVx4_ASAP7_75t_L g877 ( 
.A(n_634),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_731),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_669),
.B(n_439),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_663),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_646),
.A2(n_241),
.B(n_370),
.C(n_312),
.Y(n_881)
);

NOR2xp67_ASAP7_75t_L g882 ( 
.A(n_702),
.B(n_233),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_731),
.Y(n_883)
);

INVx8_ASAP7_75t_L g884 ( 
.A(n_710),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_698),
.A2(n_241),
.B(n_370),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_646),
.B(n_233),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_726),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_712),
.B(n_236),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_715),
.B(n_236),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_657),
.B(n_240),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_657),
.B(n_681),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_SL g892 ( 
.A1(n_726),
.A2(n_229),
.B1(n_230),
.B2(n_365),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_727),
.A2(n_487),
.B(n_484),
.C(n_443),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_725),
.B(n_240),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_676),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_738),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_633),
.B(n_242),
.Y(n_897)
);

O2A1O1Ixp33_ASAP7_75t_SL g898 ( 
.A1(n_741),
.A2(n_727),
.B(n_670),
.C(n_667),
.Y(n_898)
);

BUFx8_ASAP7_75t_L g899 ( 
.A(n_756),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_752),
.A2(n_630),
.B(n_649),
.C(n_651),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_746),
.B(n_653),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_772),
.A2(n_645),
.B(n_608),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_772),
.A2(n_835),
.B(n_777),
.Y(n_903)
);

AOI21x1_ASAP7_75t_L g904 ( 
.A1(n_810),
.A2(n_655),
.B(n_680),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_749),
.B(n_738),
.Y(n_905)
);

INVx11_ASAP7_75t_L g906 ( 
.A(n_768),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_757),
.B(n_738),
.Y(n_907)
);

AOI21x1_ASAP7_75t_L g908 ( 
.A1(n_810),
.A2(n_682),
.B(n_680),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_747),
.B(n_798),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_776),
.A2(n_645),
.B(n_608),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_774),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_743),
.B(n_778),
.Y(n_912)
);

AO21x1_ASAP7_75t_L g913 ( 
.A1(n_741),
.A2(n_707),
.B(n_689),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_830),
.A2(n_659),
.B(n_608),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_798),
.B(n_633),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_879),
.B(n_633),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_778),
.B(n_738),
.Y(n_917)
);

AND2x6_ASAP7_75t_L g918 ( 
.A(n_876),
.B(n_682),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_811),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_819),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_761),
.A2(n_697),
.B(n_689),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_844),
.A2(n_659),
.B(n_683),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_876),
.A2(n_728),
.B(n_697),
.C(n_719),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_794),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_845),
.A2(n_783),
.B(n_802),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_838),
.B(n_666),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_850),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_841),
.A2(n_659),
.B(n_701),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_780),
.B(n_718),
.Y(n_929)
);

OAI21xp33_ASAP7_75t_L g930 ( 
.A1(n_755),
.A2(n_374),
.B(n_238),
.Y(n_930)
);

CKINVDCx10_ASAP7_75t_R g931 ( 
.A(n_756),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_849),
.A2(n_683),
.B(n_696),
.Y(n_932)
);

BUFx4f_ASAP7_75t_L g933 ( 
.A(n_791),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_782),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_780),
.B(n_718),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_818),
.B(n_703),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_765),
.B(n_726),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_811),
.Y(n_938)
);

BUFx2_ASAP7_75t_SL g939 ( 
.A(n_773),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_853),
.A2(n_679),
.B1(n_713),
.B2(n_703),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_811),
.B(n_828),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_818),
.B(n_713),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_831),
.B(n_709),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_821),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_831),
.B(n_709),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_865),
.A2(n_696),
.B(n_683),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_869),
.B(n_641),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_829),
.A2(n_803),
.B(n_802),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_759),
.A2(n_679),
.B1(n_728),
.B2(n_719),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_803),
.A2(n_701),
.B(n_696),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_891),
.A2(n_701),
.B(n_641),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_771),
.A2(n_641),
.B(n_707),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_785),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_744),
.A2(n_710),
.B(n_656),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_868),
.B(n_679),
.Y(n_955)
);

O2A1O1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_744),
.A2(n_484),
.B(n_442),
.C(n_443),
.Y(n_956)
);

AOI21xp33_ASAP7_75t_L g957 ( 
.A1(n_804),
.A2(n_316),
.B(n_321),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_765),
.B(n_692),
.Y(n_958)
);

AO21x1_ASAP7_75t_L g959 ( 
.A1(n_745),
.A2(n_440),
.B(n_487),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_790),
.Y(n_960)
);

O2A1O1Ixp5_ASAP7_75t_L g961 ( 
.A1(n_745),
.A2(n_442),
.B(n_710),
.C(n_668),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_760),
.B(n_894),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_791),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_758),
.A2(n_710),
.B(n_656),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_789),
.B(n_692),
.Y(n_965)
);

BUFx4f_ASAP7_75t_L g966 ( 
.A(n_791),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_758),
.A2(n_656),
.B(n_668),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_795),
.B(n_692),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_894),
.B(n_242),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_814),
.A2(n_817),
.B(n_815),
.Y(n_970)
);

BUFx4f_ASAP7_75t_L g971 ( 
.A(n_763),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_759),
.A2(n_656),
.B(n_668),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_834),
.B(n_700),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_896),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_827),
.A2(n_312),
.B(n_243),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_805),
.B(n_243),
.Y(n_976)
);

NAND2xp33_ASAP7_75t_L g977 ( 
.A(n_873),
.B(n_372),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_742),
.B(n_372),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_836),
.A2(n_389),
.B(n_393),
.Y(n_979)
);

NAND2x1p5_ASAP7_75t_L g980 ( 
.A(n_820),
.B(n_71),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_842),
.A2(n_888),
.B(n_861),
.C(n_874),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_764),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_839),
.B(n_393),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_762),
.B(n_395),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_755),
.A2(n_402),
.B1(n_401),
.B2(n_400),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_837),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_R g987 ( 
.A(n_823),
.B(n_395),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_840),
.A2(n_399),
.B1(n_326),
.B2(n_329),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_842),
.B(n_399),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_804),
.B(n_332),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_769),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_851),
.B(n_78),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_861),
.B(n_333),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_874),
.A2(n_357),
.B(n_334),
.C(n_335),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_888),
.B(n_339),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_799),
.A2(n_347),
.B(n_348),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_895),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_784),
.A2(n_355),
.B(n_356),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_806),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_792),
.B(n_232),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_R g1001 ( 
.A(n_816),
.B(n_307),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_779),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_807),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_878),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_768),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_809),
.A2(n_781),
.B(n_775),
.Y(n_1006)
);

INVx4_ASAP7_75t_L g1007 ( 
.A(n_837),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_796),
.B(n_229),
.Y(n_1008)
);

INVx4_ASAP7_75t_L g1009 ( 
.A(n_870),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_766),
.B(n_363),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_881),
.A2(n_229),
.B(n_230),
.C(n_300),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_889),
.A2(n_402),
.B1(n_401),
.B2(n_400),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_852),
.A2(n_397),
.B(n_396),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_889),
.A2(n_397),
.B(n_396),
.C(n_394),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_767),
.A2(n_394),
.B(n_392),
.C(n_383),
.Y(n_1015)
);

BUFx24_ASAP7_75t_L g1016 ( 
.A(n_790),
.Y(n_1016)
);

NAND3xp33_ASAP7_75t_L g1017 ( 
.A(n_753),
.B(n_383),
.C(n_381),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_SL g1018 ( 
.A(n_855),
.B(n_365),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_883),
.A2(n_380),
.B(n_374),
.Y(n_1019)
);

OAI321xp33_ASAP7_75t_L g1020 ( 
.A1(n_825),
.A2(n_381),
.A3(n_380),
.B1(n_371),
.B2(n_351),
.C(n_300),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_859),
.B(n_300),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_873),
.Y(n_1022)
);

NOR2x1_ASAP7_75t_L g1023 ( 
.A(n_824),
.B(n_351),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_824),
.A2(n_862),
.B(n_858),
.C(n_890),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_863),
.B(n_351),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_775),
.A2(n_86),
.B(n_193),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_880),
.A2(n_82),
.B(n_192),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_871),
.B(n_28),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_843),
.A2(n_90),
.B(n_190),
.Y(n_1029)
);

AO21x1_ASAP7_75t_L g1030 ( 
.A1(n_781),
.A2(n_29),
.B(n_30),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_843),
.A2(n_866),
.B(n_847),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_786),
.A2(n_79),
.B(n_188),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_812),
.A2(n_200),
.B(n_185),
.Y(n_1033)
);

NAND2x1p5_ASAP7_75t_L g1034 ( 
.A(n_870),
.B(n_184),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_857),
.B(n_30),
.Y(n_1035)
);

AND2x6_ASAP7_75t_SL g1036 ( 
.A(n_855),
.B(n_32),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_887),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_867),
.B(n_168),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_884),
.Y(n_1039)
);

AOI21x1_ASAP7_75t_L g1040 ( 
.A1(n_856),
.A2(n_167),
.B(n_160),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_832),
.B(n_37),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_846),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_748),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_750),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_886),
.A2(n_156),
.B1(n_149),
.B2(n_146),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_753),
.B(n_38),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_813),
.B(n_38),
.Y(n_1047)
);

AOI21x1_ASAP7_75t_L g1048 ( 
.A1(n_864),
.A2(n_142),
.B(n_141),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_877),
.B(n_140),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_848),
.B(n_40),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_788),
.B(n_42),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_860),
.B(n_45),
.Y(n_1052)
);

BUFx2_ASAP7_75t_SL g1053 ( 
.A(n_854),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_793),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_877),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_797),
.B(n_801),
.Y(n_1056)
);

NOR2xp67_ASAP7_75t_L g1057 ( 
.A(n_800),
.B(n_826),
.Y(n_1057)
);

AO21x1_ASAP7_75t_L g1058 ( 
.A1(n_872),
.A2(n_46),
.B(n_47),
.Y(n_1058)
);

BUFx12f_ASAP7_75t_L g1059 ( 
.A(n_754),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_887),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_884),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_808),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_833),
.B(n_892),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_882),
.A2(n_48),
.B(n_49),
.C(n_51),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_885),
.B(n_770),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_893),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_872),
.A2(n_138),
.B(n_126),
.Y(n_1067)
);

AOI21x1_ASAP7_75t_L g1068 ( 
.A1(n_875),
.A2(n_116),
.B(n_110),
.Y(n_1068)
);

AOI33xp33_ASAP7_75t_L g1069 ( 
.A1(n_825),
.A2(n_49),
.A3(n_51),
.B1(n_53),
.B2(n_54),
.B3(n_55),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_822),
.B(n_57),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_963),
.B(n_822),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_981),
.A2(n_897),
.B(n_875),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_963),
.B(n_855),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_912),
.B(n_770),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1054),
.B(n_787),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_908),
.A2(n_897),
.B(n_105),
.Y(n_1076)
);

NOR2x1_ASAP7_75t_SL g1077 ( 
.A(n_1022),
.B(n_104),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_990),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_903),
.A2(n_103),
.B(n_65),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_944),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1056),
.B(n_901),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1000),
.B(n_924),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_904),
.A2(n_951),
.B(n_921),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_913),
.A2(n_923),
.A3(n_959),
.B(n_949),
.Y(n_1084)
);

NOR2xp67_ASAP7_75t_L g1085 ( 
.A(n_1042),
.B(n_962),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_951),
.A2(n_946),
.B(n_914),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_903),
.A2(n_970),
.B(n_948),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_911),
.Y(n_1088)
);

AOI21x1_ASAP7_75t_L g1089 ( 
.A1(n_943),
.A2(n_945),
.B(n_935),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_905),
.B(n_907),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_970),
.A2(n_948),
.B(n_925),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_950),
.A2(n_1055),
.B(n_986),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_1070),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_SL g1094 ( 
.A1(n_1024),
.A2(n_1033),
.B(n_1022),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_937),
.B(n_918),
.Y(n_1095)
);

BUFx4f_ASAP7_75t_L g1096 ( 
.A(n_963),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_920),
.B(n_927),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_909),
.B(n_1042),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_918),
.B(n_929),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1006),
.A2(n_922),
.B(n_932),
.Y(n_1100)
);

AO21x2_ASAP7_75t_L g1101 ( 
.A1(n_1006),
.A2(n_900),
.B(n_958),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_969),
.B(n_993),
.Y(n_1102)
);

NAND2x1_ASAP7_75t_SL g1103 ( 
.A(n_1046),
.B(n_1023),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_1010),
.B(n_995),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_922),
.A2(n_932),
.B(n_928),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_989),
.B(n_934),
.Y(n_1106)
);

AOI21x1_ASAP7_75t_L g1107 ( 
.A1(n_915),
.A2(n_946),
.B(n_928),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1037),
.Y(n_1108)
);

AOI21x1_ASAP7_75t_SL g1109 ( 
.A1(n_1065),
.A2(n_1035),
.B(n_955),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_940),
.A2(n_902),
.B(n_910),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1031),
.A2(n_952),
.B(n_1061),
.Y(n_1111)
);

OAI21xp33_ASAP7_75t_L g1112 ( 
.A1(n_985),
.A2(n_930),
.B(n_957),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1041),
.B(n_1050),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1017),
.A2(n_985),
.B1(n_1063),
.B2(n_1008),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_999),
.B(n_1003),
.Y(n_1115)
);

AOI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_1019),
.A2(n_1013),
.B(n_1011),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_952),
.A2(n_1061),
.B(n_1067),
.Y(n_1117)
);

INVx3_ASAP7_75t_SL g1118 ( 
.A(n_1005),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1037),
.B(n_983),
.Y(n_1119)
);

AO21x1_ASAP7_75t_L g1120 ( 
.A1(n_1027),
.A2(n_1038),
.B(n_1029),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_982),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_953),
.B(n_965),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_992),
.B(n_919),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_938),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_968),
.B(n_919),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_997),
.B(n_1004),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_983),
.B(n_960),
.Y(n_1127)
);

NAND2x1_ASAP7_75t_L g1128 ( 
.A(n_1007),
.B(n_1009),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_918),
.B(n_991),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1057),
.A2(n_1015),
.B(n_994),
.C(n_1014),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_974),
.A2(n_1068),
.B(n_1048),
.Y(n_1131)
);

AO21x1_ASAP7_75t_L g1132 ( 
.A1(n_1011),
.A2(n_1045),
.B(n_1032),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_976),
.B(n_1052),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1009),
.A2(n_916),
.B(n_973),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_1020),
.A2(n_1064),
.B(n_1028),
.C(n_1051),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_918),
.B(n_1002),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_938),
.Y(n_1137)
);

AND3x2_ASAP7_75t_L g1138 ( 
.A(n_1018),
.B(n_926),
.C(n_1047),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_978),
.B(n_984),
.Y(n_1139)
);

BUFx10_ASAP7_75t_L g1140 ( 
.A(n_992),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_973),
.A2(n_898),
.B(n_941),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_938),
.B(n_1022),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_972),
.A2(n_1066),
.B1(n_947),
.B2(n_966),
.Y(n_1143)
);

OA21x2_ASAP7_75t_L g1144 ( 
.A1(n_954),
.A2(n_964),
.B(n_967),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_987),
.B(n_1016),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1043),
.A2(n_1044),
.B(n_1040),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1053),
.B(n_1012),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1069),
.B(n_998),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_961),
.A2(n_998),
.B(n_975),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_961),
.A2(n_975),
.B(n_979),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1022),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_979),
.A2(n_996),
.B(n_1025),
.C(n_1021),
.Y(n_1152)
);

BUFx4f_ASAP7_75t_L g1153 ( 
.A(n_980),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_977),
.A2(n_996),
.B1(n_1058),
.B2(n_988),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1034),
.A2(n_1049),
.B(n_1026),
.Y(n_1155)
);

AOI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1026),
.A2(n_1030),
.B(n_956),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_933),
.A2(n_966),
.B(n_1039),
.Y(n_1157)
);

CKINVDCx8_ASAP7_75t_R g1158 ( 
.A(n_931),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_939),
.B(n_1001),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1039),
.B(n_1049),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_933),
.A2(n_1039),
.B(n_1034),
.Y(n_1161)
);

AOI21xp33_ASAP7_75t_L g1162 ( 
.A1(n_956),
.A2(n_980),
.B(n_971),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1039),
.B(n_1062),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_971),
.A2(n_1062),
.B(n_1036),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_1059),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_906),
.A2(n_899),
.B(n_981),
.C(n_752),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1000),
.B(n_747),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_903),
.A2(n_835),
.B(n_917),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_963),
.B(n_1060),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_912),
.B(n_752),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_912),
.B(n_752),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_1037),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_912),
.B(n_752),
.Y(n_1173)
);

INVx4_ASAP7_75t_SL g1174 ( 
.A(n_918),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_944),
.Y(n_1175)
);

NAND2x1_ASAP7_75t_SL g1176 ( 
.A(n_1046),
.B(n_969),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_963),
.Y(n_1177)
);

AOI21x1_ASAP7_75t_L g1178 ( 
.A1(n_917),
.A2(n_942),
.B(n_936),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_SL g1179 ( 
.A1(n_981),
.A2(n_1024),
.B(n_917),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_912),
.B(n_752),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_938),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1037),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_912),
.B(n_752),
.Y(n_1183)
);

INVxp67_ASAP7_75t_L g1184 ( 
.A(n_944),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_908),
.A2(n_904),
.B(n_951),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_981),
.A2(n_903),
.B(n_921),
.Y(n_1186)
);

AO21x2_ASAP7_75t_L g1187 ( 
.A1(n_981),
.A2(n_921),
.B(n_925),
.Y(n_1187)
);

AND2x6_ASAP7_75t_L g1188 ( 
.A(n_1022),
.B(n_1039),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_912),
.B(n_752),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_938),
.Y(n_1190)
);

AO21x2_ASAP7_75t_L g1191 ( 
.A1(n_981),
.A2(n_921),
.B(n_925),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_903),
.A2(n_835),
.B(n_917),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_981),
.A2(n_903),
.B(n_921),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_962),
.B(n_752),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1037),
.Y(n_1195)
);

AOI21x1_ASAP7_75t_L g1196 ( 
.A1(n_917),
.A2(n_942),
.B(n_936),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_903),
.A2(n_835),
.B(n_917),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_963),
.Y(n_1198)
);

AOI221x1_ASAP7_75t_L g1199 ( 
.A1(n_981),
.A2(n_752),
.B1(n_853),
.B2(n_598),
.C(n_969),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_903),
.A2(n_835),
.B(n_917),
.Y(n_1200)
);

AOI221xp5_ASAP7_75t_L g1201 ( 
.A1(n_985),
.A2(n_753),
.B1(n_1017),
.B2(n_755),
.C(n_1046),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1016),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_981),
.A2(n_752),
.B(n_990),
.C(n_969),
.Y(n_1203)
);

AOI21xp33_ASAP7_75t_L g1204 ( 
.A1(n_990),
.A2(n_752),
.B(n_981),
.Y(n_1204)
);

AND2x6_ASAP7_75t_SL g1205 ( 
.A(n_926),
.B(n_855),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_912),
.B(n_752),
.Y(n_1206)
);

AO31x2_ASAP7_75t_L g1207 ( 
.A1(n_913),
.A2(n_981),
.A3(n_923),
.B(n_959),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_908),
.A2(n_904),
.B(n_951),
.Y(n_1208)
);

INVx6_ASAP7_75t_L g1209 ( 
.A(n_963),
.Y(n_1209)
);

AO21x2_ASAP7_75t_L g1210 ( 
.A1(n_981),
.A2(n_921),
.B(n_925),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_981),
.A2(n_903),
.B(n_921),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_963),
.B(n_1060),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_908),
.A2(n_904),
.B(n_951),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_912),
.B(n_752),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_962),
.B(n_752),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_962),
.B(n_752),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1182),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1096),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_1175),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1170),
.B(n_1171),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1113),
.B(n_1167),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1215),
.A2(n_1170),
.B1(n_1171),
.B2(n_1173),
.Y(n_1222)
);

OR2x6_ASAP7_75t_L g1223 ( 
.A(n_1157),
.B(n_1073),
.Y(n_1223)
);

OA22x2_ASAP7_75t_L g1224 ( 
.A1(n_1075),
.A2(n_1138),
.B1(n_1112),
.B2(n_1199),
.Y(n_1224)
);

CKINVDCx11_ASAP7_75t_R g1225 ( 
.A(n_1158),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1133),
.B(n_1119),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1088),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1173),
.B(n_1180),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1180),
.A2(n_1183),
.B1(n_1206),
.B2(n_1214),
.Y(n_1229)
);

NAND2xp33_ASAP7_75t_L g1230 ( 
.A(n_1203),
.B(n_1102),
.Y(n_1230)
);

AND2x2_ASAP7_75t_SL g1231 ( 
.A(n_1201),
.B(n_1153),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1126),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1096),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1082),
.B(n_1127),
.Y(n_1234)
);

OR2x2_ASAP7_75t_L g1235 ( 
.A(n_1074),
.B(n_1194),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1192),
.A2(n_1200),
.B(n_1197),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_1195),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1071),
.B(n_1123),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1093),
.B(n_1104),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1142),
.B(n_1128),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1183),
.A2(n_1214),
.B1(n_1206),
.B2(n_1189),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_1202),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1081),
.A2(n_1092),
.B(n_1091),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1091),
.A2(n_1087),
.B(n_1211),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1087),
.A2(n_1186),
.B(n_1193),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1080),
.Y(n_1246)
);

CKINVDCx8_ASAP7_75t_R g1247 ( 
.A(n_1205),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1198),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1071),
.B(n_1123),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1169),
.B(n_1212),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1118),
.Y(n_1251)
);

INVx8_ASAP7_75t_L g1252 ( 
.A(n_1188),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1085),
.B(n_1098),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1186),
.A2(n_1193),
.B(n_1211),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1081),
.B(n_1216),
.Y(n_1255)
);

CKINVDCx11_ASAP7_75t_R g1256 ( 
.A(n_1073),
.Y(n_1256)
);

NOR2x1_ASAP7_75t_SL g1257 ( 
.A(n_1160),
.B(n_1143),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1204),
.A2(n_1114),
.B1(n_1148),
.B2(n_1116),
.Y(n_1258)
);

INVxp67_ASAP7_75t_SL g1259 ( 
.A(n_1184),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1100),
.A2(n_1090),
.B(n_1105),
.Y(n_1260)
);

INVxp67_ASAP7_75t_SL g1261 ( 
.A(n_1172),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1114),
.A2(n_1139),
.B1(n_1147),
.B2(n_1106),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1097),
.B(n_1108),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1177),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1204),
.A2(n_1148),
.B1(n_1116),
.B2(n_1122),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1177),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1165),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1209),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1095),
.B(n_1097),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1095),
.A2(n_1130),
.B1(n_1153),
.B2(n_1166),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_SL g1271 ( 
.A1(n_1164),
.A2(n_1163),
.B1(n_1165),
.B2(n_1154),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1124),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1135),
.A2(n_1176),
.B(n_1072),
.C(n_1103),
.Y(n_1273)
);

BUFx12f_ASAP7_75t_L g1274 ( 
.A(n_1209),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1121),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1115),
.B(n_1159),
.Y(n_1276)
);

OA22x2_ASAP7_75t_L g1277 ( 
.A1(n_1164),
.A2(n_1115),
.B1(n_1163),
.B2(n_1072),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1145),
.A2(n_1120),
.B1(n_1143),
.B2(n_1169),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1090),
.B(n_1187),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1212),
.B(n_1142),
.Y(n_1280)
);

INVxp67_ASAP7_75t_SL g1281 ( 
.A(n_1124),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1187),
.B(n_1210),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1188),
.Y(n_1283)
);

INVx5_ASAP7_75t_L g1284 ( 
.A(n_1188),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1174),
.B(n_1151),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1124),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1132),
.A2(n_1210),
.B1(n_1191),
.B2(n_1140),
.Y(n_1287)
);

AND2x6_ASAP7_75t_L g1288 ( 
.A(n_1151),
.B(n_1160),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_1140),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1152),
.B(n_1129),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1191),
.A2(n_1110),
.B(n_1086),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1174),
.B(n_1137),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1137),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1078),
.B(n_1190),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1188),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1099),
.B(n_1125),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1099),
.B(n_1110),
.Y(n_1297)
);

INVx5_ASAP7_75t_L g1298 ( 
.A(n_1181),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1136),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1136),
.Y(n_1300)
);

OR2x6_ASAP7_75t_L g1301 ( 
.A(n_1161),
.B(n_1134),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1101),
.A2(n_1083),
.B(n_1111),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1155),
.A2(n_1141),
.B(n_1149),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1174),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1146),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1162),
.A2(n_1150),
.B1(n_1079),
.B2(n_1144),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1077),
.B(n_1207),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1207),
.Y(n_1308)
);

OA21x2_ASAP7_75t_L g1309 ( 
.A1(n_1185),
.A2(n_1213),
.B(n_1208),
.Y(n_1309)
);

CKINVDCx6p67_ASAP7_75t_R g1310 ( 
.A(n_1109),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1084),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1076),
.B(n_1117),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1089),
.B(n_1196),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1084),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1084),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1107),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1178),
.B(n_1144),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1131),
.A2(n_1201),
.B1(n_990),
.B2(n_1112),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1156),
.B(n_1170),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1088),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1071),
.B(n_1123),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1170),
.B(n_1171),
.Y(n_1322)
);

AO21x1_ASAP7_75t_L g1323 ( 
.A1(n_1204),
.A2(n_1116),
.B(n_1102),
.Y(n_1323)
);

BUFx12f_ASAP7_75t_L g1324 ( 
.A(n_1202),
.Y(n_1324)
);

CKINVDCx16_ASAP7_75t_R g1325 ( 
.A(n_1145),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1182),
.Y(n_1326)
);

BUFx4f_ASAP7_75t_SL g1327 ( 
.A(n_1198),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1182),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1074),
.B(n_747),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1104),
.A2(n_990),
.B1(n_752),
.B2(n_969),
.Y(n_1330)
);

INVx4_ASAP7_75t_L g1331 ( 
.A(n_1096),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1170),
.B(n_1171),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1158),
.Y(n_1333)
);

OAI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1102),
.A2(n_752),
.B1(n_619),
.B2(n_751),
.Y(n_1334)
);

BUFx8_ASAP7_75t_L g1335 ( 
.A(n_1145),
.Y(n_1335)
);

A2O1A1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1104),
.A2(n_1203),
.B(n_981),
.C(n_752),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1179),
.A2(n_1094),
.B(n_1203),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1170),
.B(n_1171),
.Y(n_1338)
);

O2A1O1Ixp5_ASAP7_75t_L g1339 ( 
.A1(n_1203),
.A2(n_752),
.B(n_969),
.C(n_1104),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1096),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1071),
.B(n_1123),
.Y(n_1341)
);

INVx2_ASAP7_75t_SL g1342 ( 
.A(n_1175),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1088),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1071),
.B(n_1123),
.Y(n_1344)
);

NOR2x1_ASAP7_75t_R g1345 ( 
.A(n_1202),
.B(n_823),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1170),
.B(n_1171),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1203),
.A2(n_752),
.B(n_981),
.C(n_990),
.Y(n_1347)
);

CKINVDCx20_ASAP7_75t_R g1348 ( 
.A(n_1158),
.Y(n_1348)
);

INVx2_ASAP7_75t_SL g1349 ( 
.A(n_1175),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1170),
.B(n_1171),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1104),
.A2(n_1203),
.B(n_981),
.C(n_752),
.Y(n_1351)
);

INVx4_ASAP7_75t_L g1352 ( 
.A(n_1096),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_1096),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_SL g1354 ( 
.A(n_1203),
.B(n_751),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1113),
.B(n_1167),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1188),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1094),
.A2(n_1179),
.B(n_1168),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1113),
.B(n_1167),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1201),
.A2(n_990),
.B1(n_1112),
.B2(n_969),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1096),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1252),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1330),
.B(n_1334),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1359),
.A2(n_1350),
.B1(n_1346),
.B2(n_1332),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_SL g1364 ( 
.A1(n_1354),
.A2(n_1231),
.B1(n_1224),
.B2(n_1271),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1222),
.B(n_1220),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1224),
.A2(n_1230),
.B1(n_1354),
.B2(n_1262),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1343),
.Y(n_1367)
);

INVx4_ASAP7_75t_L g1368 ( 
.A(n_1233),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_1328),
.Y(n_1369)
);

NAND2x1p5_ASAP7_75t_L g1370 ( 
.A(n_1284),
.B(n_1331),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1328),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1302),
.A2(n_1303),
.B(n_1260),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1274),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1227),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1327),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1233),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1253),
.A2(n_1276),
.B1(n_1226),
.B2(n_1358),
.Y(n_1377)
);

INVx4_ASAP7_75t_L g1378 ( 
.A(n_1233),
.Y(n_1378)
);

NAND2x1p5_ASAP7_75t_L g1379 ( 
.A(n_1284),
.B(n_1331),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1221),
.A2(n_1355),
.B1(n_1223),
.B2(n_1222),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1234),
.B(n_1239),
.Y(n_1381)
);

AOI21xp33_ASAP7_75t_L g1382 ( 
.A1(n_1347),
.A2(n_1339),
.B(n_1258),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1246),
.Y(n_1383)
);

BUFx12f_ASAP7_75t_L g1384 ( 
.A(n_1225),
.Y(n_1384)
);

NAND2x1p5_ASAP7_75t_L g1385 ( 
.A(n_1284),
.B(n_1352),
.Y(n_1385)
);

NAND2x1p5_ASAP7_75t_L g1386 ( 
.A(n_1284),
.B(n_1352),
.Y(n_1386)
);

INVxp67_ASAP7_75t_SL g1387 ( 
.A(n_1244),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1232),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1275),
.Y(n_1389)
);

BUFx12f_ASAP7_75t_L g1390 ( 
.A(n_1333),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_SL g1391 ( 
.A1(n_1337),
.A2(n_1258),
.B1(n_1270),
.B2(n_1277),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1360),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1223),
.A2(n_1270),
.B1(n_1241),
.B2(n_1229),
.Y(n_1393)
);

CKINVDCx6p67_ASAP7_75t_R g1394 ( 
.A(n_1348),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1337),
.A2(n_1277),
.B1(n_1241),
.B2(n_1357),
.Y(n_1395)
);

CKINVDCx6p67_ASAP7_75t_R g1396 ( 
.A(n_1251),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1252),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1220),
.A2(n_1322),
.B1(n_1346),
.B2(n_1350),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_1248),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1254),
.A2(n_1235),
.B1(n_1229),
.B2(n_1245),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1329),
.B(n_1269),
.Y(n_1401)
);

OAI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1228),
.A2(n_1338),
.B1(n_1332),
.B2(n_1322),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1252),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1299),
.Y(n_1404)
);

AO21x1_ASAP7_75t_SL g1405 ( 
.A1(n_1319),
.A2(n_1278),
.B(n_1279),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1263),
.B(n_1238),
.Y(n_1406)
);

CKINVDCx6p67_ASAP7_75t_R g1407 ( 
.A(n_1218),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1340),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1317),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1228),
.A2(n_1338),
.B1(n_1336),
.B2(n_1351),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1313),
.A2(n_1243),
.B(n_1323),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1326),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1300),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1255),
.A2(n_1259),
.B1(n_1318),
.B2(n_1273),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1279),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1305),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1255),
.Y(n_1417)
);

AOI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1313),
.A2(n_1265),
.B(n_1319),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1340),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_1335),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1217),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1325),
.A2(n_1257),
.B1(n_1223),
.B2(n_1265),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1296),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1282),
.Y(n_1424)
);

OR2x6_ASAP7_75t_L g1425 ( 
.A(n_1301),
.B(n_1294),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1290),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1315),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1238),
.A2(n_1341),
.B1(n_1321),
.B2(n_1249),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1296),
.B(n_1249),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1321),
.B(n_1341),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1344),
.B(n_1250),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1261),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1344),
.B(n_1250),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1310),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1297),
.A2(n_1237),
.B1(n_1256),
.B2(n_1308),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1286),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1297),
.B(n_1280),
.Y(n_1437)
);

INVxp67_ASAP7_75t_L g1438 ( 
.A(n_1219),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1340),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1316),
.A2(n_1306),
.B(n_1309),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1282),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1311),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1280),
.B(n_1349),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1292),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1314),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1281),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1353),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1307),
.Y(n_1448)
);

OR2x6_ASAP7_75t_L g1449 ( 
.A(n_1301),
.B(n_1240),
.Y(n_1449)
);

INVx5_ASAP7_75t_L g1450 ( 
.A(n_1353),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1288),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1287),
.A2(n_1301),
.B1(n_1288),
.B2(n_1335),
.Y(n_1452)
);

CKINVDCx11_ASAP7_75t_R g1453 ( 
.A(n_1247),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1288),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1288),
.Y(n_1455)
);

BUFx8_ASAP7_75t_L g1456 ( 
.A(n_1353),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1360),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1298),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1285),
.B(n_1292),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1298),
.Y(n_1460)
);

NAND2x1p5_ASAP7_75t_L g1461 ( 
.A(n_1304),
.B(n_1298),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1267),
.A2(n_1289),
.B1(n_1242),
.B2(n_1324),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1312),
.A2(n_1309),
.B(n_1304),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1272),
.Y(n_1464)
);

INVx4_ASAP7_75t_L g1465 ( 
.A(n_1360),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1342),
.B(n_1293),
.Y(n_1466)
);

INVxp67_ASAP7_75t_SL g1467 ( 
.A(n_1283),
.Y(n_1467)
);

OAI21xp33_ASAP7_75t_L g1468 ( 
.A1(n_1268),
.A2(n_1266),
.B(n_1240),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1295),
.A2(n_1356),
.B(n_1272),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1264),
.B(n_1345),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1330),
.A2(n_752),
.B1(n_1215),
.B2(n_1104),
.Y(n_1471)
);

INVx4_ASAP7_75t_L g1472 ( 
.A(n_1233),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1300),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1225),
.Y(n_1474)
);

AO21x1_ASAP7_75t_L g1475 ( 
.A1(n_1354),
.A2(n_1116),
.B(n_1330),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1330),
.B(n_1215),
.Y(n_1476)
);

NAND2x1p5_ASAP7_75t_L g1477 ( 
.A(n_1284),
.B(n_1331),
.Y(n_1477)
);

INVx8_ASAP7_75t_L g1478 ( 
.A(n_1252),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1320),
.Y(n_1479)
);

CKINVDCx6p67_ASAP7_75t_R g1480 ( 
.A(n_1225),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1223),
.B(n_1337),
.Y(n_1481)
);

INVx1_ASAP7_75t_SL g1482 ( 
.A(n_1328),
.Y(n_1482)
);

INVx6_ASAP7_75t_L g1483 ( 
.A(n_1233),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1320),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1225),
.Y(n_1485)
);

INVx4_ASAP7_75t_L g1486 ( 
.A(n_1233),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1260),
.A2(n_1291),
.B(n_1236),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1320),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1330),
.A2(n_752),
.B1(n_1215),
.B2(n_1104),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1221),
.B(n_1355),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1252),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1320),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1300),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1300),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1300),
.Y(n_1495)
);

AO21x2_ASAP7_75t_L g1496 ( 
.A1(n_1382),
.A2(n_1475),
.B(n_1372),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1426),
.B(n_1409),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1424),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1403),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1383),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1485),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1441),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1448),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1473),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1415),
.B(n_1426),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1415),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1442),
.Y(n_1507)
);

INVx3_ASAP7_75t_SL g1508 ( 
.A(n_1480),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1409),
.B(n_1448),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1432),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1445),
.Y(n_1511)
);

NOR2x1_ASAP7_75t_R g1512 ( 
.A(n_1384),
.B(n_1474),
.Y(n_1512)
);

BUFx4f_ASAP7_75t_SL g1513 ( 
.A(n_1384),
.Y(n_1513)
);

INVxp67_ASAP7_75t_SL g1514 ( 
.A(n_1493),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1391),
.B(n_1400),
.Y(n_1515)
);

INVxp67_ASAP7_75t_L g1516 ( 
.A(n_1381),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1476),
.B(n_1471),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1387),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1400),
.B(n_1387),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1418),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1489),
.A2(n_1362),
.B(n_1366),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1425),
.B(n_1449),
.Y(n_1522)
);

CKINVDCx6p67_ASAP7_75t_R g1523 ( 
.A(n_1480),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1425),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1423),
.B(n_1429),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1398),
.B(n_1417),
.Y(n_1526)
);

INVx6_ASAP7_75t_L g1527 ( 
.A(n_1456),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1490),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1427),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1463),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1494),
.Y(n_1531)
);

INVx2_ASAP7_75t_SL g1532 ( 
.A(n_1495),
.Y(n_1532)
);

BUFx12f_ASAP7_75t_L g1533 ( 
.A(n_1474),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1413),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1374),
.Y(n_1535)
);

AO21x2_ASAP7_75t_L g1536 ( 
.A1(n_1440),
.A2(n_1393),
.B(n_1365),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1401),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1405),
.B(n_1437),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1411),
.Y(n_1539)
);

AO21x2_ASAP7_75t_L g1540 ( 
.A1(n_1402),
.A2(n_1362),
.B(n_1451),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1425),
.B(n_1364),
.Y(n_1541)
);

OA21x2_ASAP7_75t_L g1542 ( 
.A1(n_1366),
.A2(n_1452),
.B(n_1455),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1404),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1449),
.B(n_1454),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1481),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1449),
.B(n_1481),
.Y(n_1546)
);

OAI21xp33_ASAP7_75t_SL g1547 ( 
.A1(n_1452),
.A2(n_1388),
.B(n_1481),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1456),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1403),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1395),
.B(n_1380),
.Y(n_1550)
);

INVxp67_ASAP7_75t_L g1551 ( 
.A(n_1421),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_1369),
.Y(n_1552)
);

INVx2_ASAP7_75t_SL g1553 ( 
.A(n_1416),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1371),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1487),
.A2(n_1410),
.B(n_1414),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1363),
.B(n_1402),
.Y(n_1556)
);

BUFx3_ASAP7_75t_L g1557 ( 
.A(n_1456),
.Y(n_1557)
);

OAI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1422),
.A2(n_1377),
.B(n_1435),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1482),
.B(n_1412),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1492),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_SL g1561 ( 
.A(n_1375),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1367),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1479),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1435),
.A2(n_1434),
.B1(n_1468),
.B2(n_1406),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1484),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1488),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1446),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1436),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1389),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1467),
.Y(n_1570)
);

CKINVDCx12_ASAP7_75t_R g1571 ( 
.A(n_1443),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1467),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1431),
.B(n_1461),
.Y(n_1573)
);

OAI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1438),
.A2(n_1466),
.B(n_1385),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1461),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1458),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1460),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1361),
.B(n_1491),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1469),
.Y(n_1579)
);

OAI21x1_ASAP7_75t_L g1580 ( 
.A1(n_1397),
.A2(n_1491),
.B(n_1469),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1397),
.A2(n_1477),
.B(n_1370),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1376),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1428),
.B(n_1464),
.Y(n_1583)
);

INVx4_ASAP7_75t_L g1584 ( 
.A(n_1478),
.Y(n_1584)
);

OA21x2_ASAP7_75t_L g1585 ( 
.A1(n_1459),
.A2(n_1433),
.B(n_1430),
.Y(n_1585)
);

AO21x1_ASAP7_75t_SL g1586 ( 
.A1(n_1462),
.A2(n_1478),
.B(n_1370),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1379),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1505),
.B(n_1396),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1524),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1519),
.B(n_1509),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1526),
.B(n_1450),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_1524),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1500),
.B(n_1394),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1505),
.B(n_1506),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1503),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1579),
.Y(n_1596)
);

BUFx2_ASAP7_75t_SL g1597 ( 
.A(n_1561),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1579),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1546),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1517),
.B(n_1450),
.Y(n_1600)
);

OAI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1521),
.A2(n_1420),
.B1(n_1396),
.B2(n_1386),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1504),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1585),
.B(n_1444),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1536),
.B(n_1399),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1585),
.B(n_1444),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1550),
.A2(n_1453),
.B1(n_1470),
.B2(n_1459),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1530),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1585),
.B(n_1497),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1530),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1544),
.Y(n_1610)
);

OAI221xp5_ASAP7_75t_L g1611 ( 
.A1(n_1558),
.A2(n_1477),
.B1(n_1386),
.B2(n_1385),
.C(n_1379),
.Y(n_1611)
);

OAI211xp5_ASAP7_75t_SL g1612 ( 
.A1(n_1564),
.A2(n_1453),
.B(n_1439),
.C(n_1419),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1556),
.B(n_1450),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1536),
.B(n_1470),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1546),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1536),
.B(n_1403),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1544),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1532),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1532),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1540),
.B(n_1403),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1540),
.B(n_1470),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1544),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1522),
.Y(n_1623)
);

AO21x2_ASAP7_75t_L g1624 ( 
.A1(n_1539),
.A2(n_1478),
.B(n_1447),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1520),
.B(n_1373),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1546),
.B(n_1545),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1540),
.B(n_1447),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1518),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1515),
.B(n_1447),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1515),
.B(n_1447),
.Y(n_1630)
);

INVxp67_ASAP7_75t_SL g1631 ( 
.A(n_1570),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1518),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1550),
.A2(n_1390),
.B1(n_1373),
.B2(n_1420),
.Y(n_1633)
);

INVxp67_ASAP7_75t_L g1634 ( 
.A(n_1537),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1538),
.B(n_1457),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_1559),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1510),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1538),
.B(n_1457),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1520),
.B(n_1392),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1522),
.Y(n_1640)
);

INVxp67_ASAP7_75t_L g1641 ( 
.A(n_1552),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1555),
.A2(n_1486),
.B(n_1368),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1498),
.B(n_1368),
.Y(n_1643)
);

INVx3_ASAP7_75t_L g1644 ( 
.A(n_1580),
.Y(n_1644)
);

NAND4xp25_ASAP7_75t_SL g1645 ( 
.A(n_1633),
.B(n_1547),
.C(n_1606),
.D(n_1621),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1608),
.B(n_1545),
.Y(n_1646)
);

OAI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1611),
.A2(n_1574),
.B1(n_1528),
.B2(n_1525),
.C(n_1516),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1608),
.B(n_1545),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1590),
.B(n_1603),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1607),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1601),
.B(n_1522),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1590),
.B(n_1496),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1603),
.B(n_1496),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1605),
.B(n_1496),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1634),
.B(n_1514),
.Y(n_1655)
);

NAND4xp25_ASAP7_75t_L g1656 ( 
.A(n_1636),
.B(n_1554),
.C(n_1551),
.D(n_1534),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1641),
.A2(n_1541),
.B1(n_1527),
.B2(n_1583),
.Y(n_1657)
);

AND2x2_ASAP7_75t_SL g1658 ( 
.A(n_1621),
.B(n_1541),
.Y(n_1658)
);

OAI221xp5_ASAP7_75t_SL g1659 ( 
.A1(n_1611),
.A2(n_1583),
.B1(n_1573),
.B2(n_1523),
.C(n_1548),
.Y(n_1659)
);

OAI221xp5_ASAP7_75t_SL g1660 ( 
.A1(n_1614),
.A2(n_1573),
.B1(n_1523),
.B2(n_1548),
.C(n_1557),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1602),
.B(n_1531),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1596),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1594),
.B(n_1502),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1600),
.B(n_1501),
.Y(n_1664)
);

OAI221xp5_ASAP7_75t_SL g1665 ( 
.A1(n_1614),
.A2(n_1557),
.B1(n_1568),
.B2(n_1577),
.C(n_1576),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_L g1666 ( 
.A(n_1604),
.B(n_1543),
.C(n_1565),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1626),
.B(n_1529),
.Y(n_1667)
);

OAI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1612),
.A2(n_1508),
.B1(n_1501),
.B2(n_1587),
.C(n_1527),
.Y(n_1668)
);

OAI211xp5_ASAP7_75t_L g1669 ( 
.A1(n_1613),
.A2(n_1542),
.B(n_1535),
.C(n_1555),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1626),
.B(n_1542),
.Y(n_1670)
);

OAI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1600),
.A2(n_1508),
.B1(n_1587),
.B2(n_1527),
.C(n_1486),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1613),
.A2(n_1527),
.B1(n_1542),
.B2(n_1508),
.Y(n_1672)
);

OAI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1593),
.A2(n_1378),
.B1(n_1472),
.B2(n_1465),
.C(n_1408),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1591),
.A2(n_1567),
.B1(n_1572),
.B2(n_1561),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1591),
.B(n_1578),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1595),
.B(n_1560),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1610),
.B(n_1617),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_L g1678 ( 
.A(n_1604),
.B(n_1566),
.C(n_1565),
.Y(n_1678)
);

OAI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1588),
.A2(n_1472),
.B1(n_1408),
.B2(n_1378),
.C(n_1465),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1618),
.B(n_1619),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1597),
.A2(n_1586),
.B1(n_1561),
.B2(n_1513),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1597),
.A2(n_1586),
.B1(n_1533),
.B2(n_1575),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1617),
.B(n_1507),
.Y(n_1683)
);

OAI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1588),
.A2(n_1376),
.B1(n_1392),
.B2(n_1483),
.C(n_1562),
.Y(n_1684)
);

OAI21xp33_ASAP7_75t_SL g1685 ( 
.A1(n_1637),
.A2(n_1581),
.B(n_1553),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1622),
.B(n_1507),
.Y(n_1686)
);

NAND3xp33_ASAP7_75t_L g1687 ( 
.A(n_1625),
.B(n_1643),
.C(n_1639),
.Y(n_1687)
);

NAND2x1p5_ASAP7_75t_L g1688 ( 
.A(n_1620),
.B(n_1580),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1628),
.B(n_1632),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_SL g1690 ( 
.A1(n_1620),
.A2(n_1533),
.B1(n_1581),
.B2(n_1549),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1622),
.B(n_1511),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1627),
.B(n_1511),
.Y(n_1692)
);

NAND3xp33_ASAP7_75t_L g1693 ( 
.A(n_1625),
.B(n_1569),
.C(n_1563),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1692),
.B(n_1652),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1662),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1649),
.B(n_1616),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1645),
.A2(n_1615),
.B1(n_1599),
.B2(n_1640),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1662),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1650),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1646),
.B(n_1616),
.Y(n_1700)
);

NOR2x1p5_ASAP7_75t_L g1701 ( 
.A(n_1656),
.B(n_1623),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1692),
.B(n_1596),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1650),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1689),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1648),
.B(n_1627),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1689),
.Y(n_1706)
);

NOR2xp67_ASAP7_75t_L g1707 ( 
.A(n_1685),
.B(n_1644),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1688),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1685),
.Y(n_1709)
);

BUFx2_ASAP7_75t_L g1710 ( 
.A(n_1688),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1652),
.B(n_1680),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1678),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1658),
.B(n_1589),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1658),
.B(n_1592),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1670),
.Y(n_1715)
);

NOR2x1_ASAP7_75t_SL g1716 ( 
.A(n_1678),
.B(n_1624),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1658),
.B(n_1592),
.Y(n_1717)
);

NOR2x1p5_ASAP7_75t_L g1718 ( 
.A(n_1656),
.B(n_1623),
.Y(n_1718)
);

AND2x2_ASAP7_75t_SL g1719 ( 
.A(n_1681),
.B(n_1615),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1687),
.B(n_1609),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1663),
.Y(n_1721)
);

NAND2x1p5_ASAP7_75t_L g1722 ( 
.A(n_1651),
.B(n_1637),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_1677),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1677),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1663),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1676),
.Y(n_1726)
);

NOR2x1_ASAP7_75t_L g1727 ( 
.A(n_1666),
.B(n_1598),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1687),
.B(n_1609),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1693),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1653),
.B(n_1609),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1653),
.B(n_1631),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1693),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1712),
.Y(n_1733)
);

AOI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1697),
.A2(n_1647),
.B1(n_1657),
.B2(n_1719),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1709),
.B(n_1654),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1703),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1705),
.B(n_1667),
.Y(n_1737)
);

OAI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1727),
.A2(n_1672),
.B(n_1659),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1729),
.B(n_1654),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1705),
.B(n_1688),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1695),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1695),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1698),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1698),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1699),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1699),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1729),
.B(n_1655),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1709),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1699),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1722),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1708),
.B(n_1710),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1700),
.B(n_1690),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1704),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1703),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1703),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1704),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1706),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1696),
.B(n_1683),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1706),
.Y(n_1759)
);

INVxp67_ASAP7_75t_SL g1760 ( 
.A(n_1727),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1732),
.B(n_1686),
.Y(n_1761)
);

NOR2xp67_ASAP7_75t_L g1762 ( 
.A(n_1712),
.B(n_1669),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1715),
.B(n_1672),
.Y(n_1763)
);

OAI21xp33_ASAP7_75t_L g1764 ( 
.A1(n_1732),
.A2(n_1665),
.B(n_1657),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1723),
.B(n_1691),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1728),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1728),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1720),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1720),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1703),
.Y(n_1770)
);

INVx3_ASAP7_75t_SL g1771 ( 
.A(n_1719),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1730),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1730),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1723),
.B(n_1691),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1702),
.Y(n_1775)
);

OAI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1738),
.A2(n_1719),
.B(n_1722),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1741),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1741),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1742),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1764),
.B(n_1747),
.Y(n_1780)
);

AOI211xp5_ASAP7_75t_SL g1781 ( 
.A1(n_1762),
.A2(n_1660),
.B(n_1668),
.C(n_1671),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1751),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1764),
.B(n_1726),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1742),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1747),
.B(n_1711),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1743),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1736),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1771),
.B(n_1710),
.Y(n_1788)
);

OAI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1738),
.A2(n_1722),
.B(n_1674),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1771),
.B(n_1713),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1743),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1771),
.B(n_1713),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1744),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1744),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1736),
.Y(n_1795)
);

OAI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1734),
.A2(n_1762),
.B1(n_1701),
.B2(n_1718),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1753),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1739),
.B(n_1711),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1739),
.B(n_1694),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1752),
.B(n_1726),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1735),
.B(n_1714),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1735),
.B(n_1714),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1761),
.B(n_1721),
.Y(n_1803)
);

NOR2x1_ASAP7_75t_L g1804 ( 
.A(n_1748),
.B(n_1701),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1736),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1753),
.Y(n_1806)
);

INVx2_ASAP7_75t_SL g1807 ( 
.A(n_1751),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1735),
.B(n_1748),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1761),
.B(n_1721),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1768),
.B(n_1694),
.Y(n_1810)
);

AND2x2_ASAP7_75t_SL g1811 ( 
.A(n_1733),
.B(n_1682),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1756),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1766),
.B(n_1725),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1756),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1768),
.B(n_1731),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1757),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1757),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1769),
.B(n_1731),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1769),
.B(n_1725),
.Y(n_1819)
);

OAI21xp33_ASAP7_75t_L g1820 ( 
.A1(n_1734),
.A2(n_1674),
.B(n_1675),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1759),
.Y(n_1821)
);

INVx1_ASAP7_75t_SL g1822 ( 
.A(n_1808),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1783),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1777),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1778),
.Y(n_1825)
);

CKINVDCx16_ASAP7_75t_R g1826 ( 
.A(n_1796),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1779),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1784),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1808),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1786),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1780),
.B(n_1752),
.Y(n_1831)
);

INVx3_ASAP7_75t_L g1832 ( 
.A(n_1782),
.Y(n_1832)
);

NAND3xp33_ASAP7_75t_SL g1833 ( 
.A(n_1789),
.B(n_1733),
.C(n_1750),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1800),
.B(n_1766),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1791),
.Y(n_1835)
);

AND4x1_ASAP7_75t_L g1836 ( 
.A(n_1781),
.B(n_1804),
.C(n_1776),
.D(n_1820),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1793),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1785),
.B(n_1815),
.Y(n_1838)
);

OA21x2_ASAP7_75t_L g1839 ( 
.A1(n_1787),
.A2(n_1760),
.B(n_1755),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1794),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1797),
.Y(n_1841)
);

OR2x6_ASAP7_75t_L g1842 ( 
.A(n_1790),
.B(n_1718),
.Y(n_1842)
);

INVx3_ASAP7_75t_L g1843 ( 
.A(n_1782),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1790),
.B(n_1760),
.Y(n_1844)
);

INVx1_ASAP7_75t_SL g1845 ( 
.A(n_1811),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1792),
.B(n_1751),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1792),
.B(n_1801),
.Y(n_1847)
);

CKINVDCx16_ASAP7_75t_R g1848 ( 
.A(n_1788),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_SL g1849 ( 
.A(n_1811),
.B(n_1750),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1815),
.B(n_1767),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1801),
.B(n_1751),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1800),
.B(n_1767),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1806),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1812),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1814),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1816),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1817),
.Y(n_1857)
);

BUFx2_ASAP7_75t_L g1858 ( 
.A(n_1782),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1821),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1802),
.B(n_1740),
.Y(n_1860)
);

INVxp67_ASAP7_75t_L g1861 ( 
.A(n_1845),
.Y(n_1861)
);

AOI222xp33_ASAP7_75t_L g1862 ( 
.A1(n_1823),
.A2(n_1788),
.B1(n_1512),
.B2(n_1716),
.C1(n_1809),
.C2(n_1803),
.Y(n_1862)
);

A2O1A1Ixp33_ASAP7_75t_L g1863 ( 
.A1(n_1849),
.A2(n_1802),
.B(n_1707),
.C(n_1763),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1830),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1830),
.Y(n_1865)
);

AOI22x1_ASAP7_75t_L g1866 ( 
.A1(n_1826),
.A2(n_1807),
.B1(n_1390),
.B2(n_1818),
.Y(n_1866)
);

AO32x1_ASAP7_75t_L g1867 ( 
.A1(n_1829),
.A2(n_1807),
.A3(n_1805),
.B1(n_1795),
.B2(n_1787),
.Y(n_1867)
);

AOI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1848),
.A2(n_1763),
.B1(n_1813),
.B2(n_1708),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1849),
.A2(n_1716),
.B(n_1664),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1822),
.B(n_1759),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1835),
.Y(n_1871)
);

OAI21xp33_ASAP7_75t_SL g1872 ( 
.A1(n_1847),
.A2(n_1798),
.B(n_1799),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1833),
.A2(n_1763),
.B1(n_1708),
.B2(n_1717),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1835),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1847),
.B(n_1740),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1836),
.B(n_1485),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1837),
.Y(n_1877)
);

OA21x2_ASAP7_75t_L g1878 ( 
.A1(n_1858),
.A2(n_1805),
.B(n_1795),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1846),
.B(n_1737),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1846),
.B(n_1737),
.Y(n_1880)
);

INVx2_ASAP7_75t_SL g1881 ( 
.A(n_1858),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1831),
.A2(n_1798),
.B1(n_1724),
.B2(n_1684),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1837),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1829),
.B(n_1818),
.Y(n_1884)
);

AND2x2_ASAP7_75t_SL g1885 ( 
.A(n_1844),
.B(n_1834),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1844),
.B(n_1775),
.Y(n_1886)
);

NOR3xp33_ASAP7_75t_SL g1887 ( 
.A(n_1852),
.B(n_1673),
.C(n_1679),
.Y(n_1887)
);

AOI211xp5_ASAP7_75t_L g1888 ( 
.A1(n_1844),
.A2(n_1707),
.B(n_1375),
.C(n_1810),
.Y(n_1888)
);

BUFx2_ASAP7_75t_L g1889 ( 
.A(n_1832),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1889),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1861),
.B(n_1860),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1881),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1884),
.B(n_1838),
.Y(n_1893)
);

CKINVDCx16_ASAP7_75t_R g1894 ( 
.A(n_1876),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1885),
.B(n_1860),
.Y(n_1895)
);

NOR2x1_ASAP7_75t_L g1896 ( 
.A(n_1864),
.B(n_1832),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1865),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1878),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1879),
.B(n_1851),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1887),
.B(n_1851),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1880),
.B(n_1824),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1871),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1875),
.B(n_1832),
.Y(n_1903)
);

INVxp33_ASAP7_75t_L g1904 ( 
.A(n_1866),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1878),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1874),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1872),
.B(n_1825),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1869),
.B(n_1838),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1877),
.B(n_1827),
.Y(n_1909)
);

INVx3_ASAP7_75t_L g1910 ( 
.A(n_1883),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1863),
.B(n_1843),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1868),
.B(n_1843),
.Y(n_1912)
);

NAND3xp33_ASAP7_75t_L g1913 ( 
.A(n_1890),
.B(n_1862),
.C(n_1888),
.Y(n_1913)
);

AOI321xp33_ASAP7_75t_L g1914 ( 
.A1(n_1908),
.A2(n_1873),
.A3(n_1888),
.B1(n_1882),
.B2(n_1886),
.C(n_1862),
.Y(n_1914)
);

NAND3xp33_ASAP7_75t_SL g1915 ( 
.A(n_1904),
.B(n_1882),
.C(n_1870),
.Y(n_1915)
);

NOR2xp33_ASAP7_75t_L g1916 ( 
.A(n_1894),
.B(n_1900),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1892),
.B(n_1828),
.Y(n_1917)
);

AOI221xp5_ASAP7_75t_SL g1918 ( 
.A1(n_1907),
.A2(n_1870),
.B1(n_1854),
.B2(n_1853),
.C(n_1859),
.Y(n_1918)
);

OAI21xp5_ASAP7_75t_SL g1919 ( 
.A1(n_1895),
.A2(n_1841),
.B(n_1840),
.Y(n_1919)
);

O2A1O1Ixp33_ASAP7_75t_L g1920 ( 
.A1(n_1898),
.A2(n_1857),
.B(n_1856),
.C(n_1855),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1910),
.Y(n_1921)
);

OAI211xp5_ASAP7_75t_L g1922 ( 
.A1(n_1896),
.A2(n_1843),
.B(n_1839),
.C(n_1867),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1892),
.B(n_1850),
.Y(n_1923)
);

NOR2xp33_ASAP7_75t_L g1924 ( 
.A(n_1894),
.B(n_1842),
.Y(n_1924)
);

OAI221xp5_ASAP7_75t_L g1925 ( 
.A1(n_1891),
.A2(n_1842),
.B1(n_1850),
.B2(n_1810),
.C(n_1799),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1893),
.B(n_1842),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1916),
.B(n_1899),
.Y(n_1927)
);

NAND5xp2_ASAP7_75t_L g1928 ( 
.A(n_1914),
.B(n_1911),
.C(n_1912),
.D(n_1899),
.E(n_1901),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1921),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1924),
.B(n_1893),
.Y(n_1930)
);

NOR3xp33_ASAP7_75t_SL g1931 ( 
.A(n_1915),
.B(n_1909),
.C(n_1902),
.Y(n_1931)
);

INVxp33_ASAP7_75t_L g1932 ( 
.A(n_1926),
.Y(n_1932)
);

AOI211xp5_ASAP7_75t_L g1933 ( 
.A1(n_1913),
.A2(n_1911),
.B(n_1912),
.C(n_1905),
.Y(n_1933)
);

NAND3xp33_ASAP7_75t_SL g1934 ( 
.A(n_1922),
.B(n_1905),
.C(n_1903),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1923),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1917),
.Y(n_1936)
);

NAND3xp33_ASAP7_75t_L g1937 ( 
.A(n_1920),
.B(n_1896),
.C(n_1897),
.Y(n_1937)
);

NOR3xp33_ASAP7_75t_L g1938 ( 
.A(n_1925),
.B(n_1910),
.C(n_1902),
.Y(n_1938)
);

NAND4xp25_ASAP7_75t_SL g1939 ( 
.A(n_1933),
.B(n_1918),
.C(n_1903),
.D(n_1906),
.Y(n_1939)
);

NAND3xp33_ASAP7_75t_SL g1940 ( 
.A(n_1931),
.B(n_1919),
.C(n_1906),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1929),
.Y(n_1941)
);

AOI211xp5_ASAP7_75t_L g1942 ( 
.A1(n_1934),
.A2(n_1897),
.B(n_1910),
.C(n_1867),
.Y(n_1942)
);

NOR4xp25_ASAP7_75t_L g1943 ( 
.A(n_1937),
.B(n_1867),
.C(n_1819),
.D(n_1839),
.Y(n_1943)
);

NAND5xp2_ASAP7_75t_L g1944 ( 
.A(n_1930),
.B(n_1717),
.C(n_1630),
.D(n_1629),
.E(n_1642),
.Y(n_1944)
);

AOI32xp33_ASAP7_75t_L g1945 ( 
.A1(n_1938),
.A2(n_1708),
.A3(n_1774),
.B1(n_1765),
.B2(n_1724),
.Y(n_1945)
);

AOI211xp5_ASAP7_75t_L g1946 ( 
.A1(n_1928),
.A2(n_1819),
.B(n_1842),
.C(n_1773),
.Y(n_1946)
);

OAI211xp5_ASAP7_75t_L g1947 ( 
.A1(n_1927),
.A2(n_1839),
.B(n_1773),
.C(n_1772),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1941),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1943),
.B(n_1932),
.Y(n_1949)
);

AOI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1940),
.A2(n_1935),
.B1(n_1936),
.B2(n_1407),
.Y(n_1950)
);

NOR3xp33_ASAP7_75t_L g1951 ( 
.A(n_1939),
.B(n_1584),
.C(n_1661),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1946),
.B(n_1775),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1942),
.B(n_1758),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1947),
.Y(n_1954)
);

NOR2x1_ASAP7_75t_L g1955 ( 
.A(n_1949),
.B(n_1948),
.Y(n_1955)
);

NAND3xp33_ASAP7_75t_L g1956 ( 
.A(n_1954),
.B(n_1945),
.C(n_1944),
.Y(n_1956)
);

AOI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1953),
.A2(n_1723),
.B1(n_1772),
.B2(n_1765),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1952),
.Y(n_1958)
);

NAND4xp25_ASAP7_75t_L g1959 ( 
.A(n_1950),
.B(n_1584),
.C(n_1638),
.D(n_1635),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1951),
.B(n_1772),
.Y(n_1960)
);

OAI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1955),
.A2(n_1746),
.B(n_1745),
.Y(n_1961)
);

NOR2xp67_ASAP7_75t_L g1962 ( 
.A(n_1956),
.B(n_1754),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1958),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1957),
.B(n_1758),
.Y(n_1964)
);

AOI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1962),
.A2(n_1960),
.B1(n_1959),
.B2(n_1483),
.Y(n_1965)
);

CKINVDCx16_ASAP7_75t_R g1966 ( 
.A(n_1965),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1966),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1966),
.A2(n_1963),
.B1(n_1964),
.B2(n_1961),
.Y(n_1968)
);

OAI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1967),
.A2(n_1770),
.B1(n_1755),
.B2(n_1754),
.Y(n_1969)
);

HB1xp67_ASAP7_75t_L g1970 ( 
.A(n_1968),
.Y(n_1970)
);

NOR2xp67_ASAP7_75t_L g1971 ( 
.A(n_1970),
.B(n_1584),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1969),
.A2(n_1746),
.B(n_1745),
.Y(n_1972)
);

OAI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1971),
.A2(n_1483),
.B1(n_1770),
.B2(n_1755),
.Y(n_1973)
);

AOI22xp5_ASAP7_75t_SL g1974 ( 
.A1(n_1973),
.A2(n_1972),
.B1(n_1582),
.B2(n_1499),
.Y(n_1974)
);

OAI221xp5_ASAP7_75t_R g1975 ( 
.A1(n_1974),
.A2(n_1770),
.B1(n_1754),
.B2(n_1749),
.C(n_1571),
.Y(n_1975)
);

AOI211xp5_ASAP7_75t_L g1976 ( 
.A1(n_1975),
.A2(n_1582),
.B(n_1549),
.C(n_1499),
.Y(n_1976)
);


endmodule