module real_jpeg_4578_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_1),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_1),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_1),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_2),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_2),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_2),
.A2(n_84),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_2),
.A2(n_84),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_2),
.A2(n_84),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_3),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_3),
.A2(n_48),
.B1(n_115),
.B2(n_119),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_3),
.A2(n_48),
.B1(n_194),
.B2(n_197),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_3),
.B(n_68),
.Y(n_284)
);

O2A1O1Ixp33_ASAP7_75t_L g339 ( 
.A1(n_3),
.A2(n_340),
.B(n_342),
.C(n_348),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_3),
.B(n_98),
.C(n_188),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_3),
.B(n_21),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_3),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_3),
.B(n_102),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_4),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_5),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_5),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_5),
.A2(n_240),
.B1(n_260),
.B2(n_263),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_5),
.A2(n_240),
.B1(n_355),
.B2(n_356),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_5),
.A2(n_240),
.B1(n_376),
.B2(n_378),
.Y(n_375)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_7),
.Y(n_190)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_7),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_7),
.Y(n_393)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_8),
.Y(n_271)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_10),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_11),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_11),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_11),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_12),
.A2(n_75),
.B1(n_77),
.B2(n_80),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_12),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_12),
.A2(n_39),
.B1(n_80),
.B2(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_12),
.A2(n_80),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_12),
.A2(n_80),
.B1(n_188),
.B2(n_276),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_13),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_13),
.Y(n_104)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_13),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_438),
.B(n_440),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_156),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_154),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_134),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_18),
.B(n_134),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_89),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_53),
.B1(n_54),
.B2(n_88),
.Y(n_19)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_20),
.A2(n_88),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_34),
.B(n_45),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_21),
.B(n_125),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_21),
.A2(n_123),
.B(n_149),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_21),
.B(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_22),
.B(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_25),
.Y(n_344)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_27),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_27),
.Y(n_179)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_27),
.Y(n_347)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_28),
.Y(n_176)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g358 ( 
.A(n_30),
.Y(n_358)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_34),
.A2(n_149),
.B(n_152),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_34),
.B(n_45),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_34),
.B(n_259),
.Y(n_282)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_35),
.B(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_38),
.Y(n_341)
);

AO22x1_ASAP7_75t_SL g68 ( 
.A1(n_39),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_68)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_41),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_44),
.Y(n_151)
);

NAND2xp33_ASAP7_75t_SL g273 ( 
.A(n_44),
.B(n_69),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g122 ( 
.A(n_45),
.Y(n_122)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_46),
.Y(n_263)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_47),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_48),
.A2(n_76),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_48),
.B(n_145),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g342 ( 
.A1(n_48),
.A2(n_343),
.B(n_345),
.Y(n_342)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_74),
.B(n_81),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_55),
.A2(n_132),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_56),
.B(n_82),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_56),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_56),
.B(n_238),
.Y(n_237)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_68),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_63),
.B2(n_66),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_68),
.B(n_143),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_68),
.B(n_238),
.Y(n_254)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_74),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI32xp33_ASAP7_75t_L g267 ( 
.A1(n_79),
.A2(n_268),
.A3(n_269),
.B1(n_272),
.B2(n_273),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_81),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_81),
.B(n_237),
.Y(n_301)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_88),
.B(n_310),
.C(n_312),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_120),
.C(n_130),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_90),
.A2(n_120),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_90),
.A2(n_140),
.B1(n_148),
.B2(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_90),
.A2(n_140),
.B1(n_256),
.B2(n_264),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_90),
.B(n_253),
.C(n_256),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_112),
.B(n_113),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_91),
.A2(n_202),
.B(n_208),
.Y(n_201)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_92),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_92),
.B(n_114),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_92),
.B(n_354),
.Y(n_353)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_102),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_96),
.Y(n_355)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_100),
.Y(n_204)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_102),
.B(n_174),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_102),
.B(n_354),
.Y(n_370)
);

AO22x1_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_105),
.B1(n_108),
.B2(n_110),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_105),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_106),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_107),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_109),
.Y(n_379)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_112),
.B(n_113),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_112),
.A2(n_173),
.B(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_SL g207 ( 
.A(n_119),
.Y(n_207)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_121),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_123),
.Y(n_257)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_129),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_131),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_133),
.B(n_254),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_141),
.C(n_147),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_135),
.A2(n_136),
.B1(n_141),
.B2(n_164),
.Y(n_244)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_141),
.C(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_142),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_143),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g272 ( 
.A(n_144),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_145),
.Y(n_241)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_147),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_153),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_153),
.B(n_282),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_246),
.B(n_434),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_242),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_212),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_160),
.B(n_212),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_181),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_168),
.B2(n_169),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_163),
.B(n_168),
.C(n_181),
.Y(n_245)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_169),
.A2(n_170),
.B(n_180),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_180),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_171),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_173),
.B(n_370),
.Y(n_414)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_209),
.B(n_210),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_182),
.A2(n_183),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_201),
.Y(n_183)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_184),
.A2(n_209),
.B1(n_210),
.B2(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_184),
.A2(n_201),
.B1(n_209),
.B2(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_184),
.B(n_339),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_184),
.A2(n_209),
.B1(n_339),
.B2(n_417),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_191),
.B(n_193),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_185),
.B(n_193),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_185),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_185),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_189),
.Y(n_192)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_197),
.Y(n_276)
);

INVx4_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_201),
.Y(n_322)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g296 ( 
.A(n_208),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_208),
.B(n_353),
.Y(n_381)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.C(n_219),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_213),
.A2(n_217),
.B1(n_218),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_213),
.Y(n_326)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_219),
.B(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_233),
.C(n_235),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_220),
.A2(n_221),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_232),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_222),
.B(n_232),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_223),
.B(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_225),
.B(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_226),
.A2(n_275),
.B(n_277),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_227),
.B(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx8_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g399 ( 
.A(n_231),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_233),
.B(n_235),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_234),
.B(n_258),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_242),
.A2(n_436),
.B(n_437),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_243),
.B(n_245),
.Y(n_437)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_426),
.Y(n_247)
);

NAND3xp33_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_315),
.C(n_329),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_304),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_290),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_251),
.B(n_290),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_265),
.C(n_280),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_252),
.B(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_265),
.A2(n_266),
.B1(n_280),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_274),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_267),
.B(n_274),
.Y(n_299)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_287),
.B(n_295),
.Y(n_294)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_279),
.Y(n_401)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_280),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.C(n_285),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_281),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_285),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_286),
.B(n_391),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_287),
.B(n_374),
.Y(n_404)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_298),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_293),
.C(n_298),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_296),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_297),
.B(n_370),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_301),
.C(n_302),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_304),
.A2(n_429),
.B(n_430),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_314),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_305),
.B(n_314),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_308),
.C(n_309),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_312),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_327),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_316),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_324),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_317),
.B(n_328),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_317),
.B(n_328),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_317),
.B(n_324),
.Y(n_433)
);

FAx1_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_321),
.CI(n_323),
.CON(n_317),
.SN(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_327),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_359),
.B(n_425),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_334),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_331),
.B(n_334),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_338),
.C(n_350),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_335),
.B(n_421),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_338),
.A2(n_350),
.B1(n_351),
.B2(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_338),
.Y(n_422)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_339),
.Y(n_417)
);

INVx8_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx6_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_347),
.Y(n_367)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx6_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_419),
.B(n_424),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_361),
.A2(n_409),
.B(n_418),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_385),
.B(n_408),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_371),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_363),
.B(n_371),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_369),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_364),
.A2(n_365),
.B1(n_369),
.B2(n_388),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_368),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_369),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_380),
.Y(n_371)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_372),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_392),
.Y(n_391)
);

INVx6_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx6_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_383),
.B2(n_384),
.Y(n_380)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_381),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_382),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_382),
.B(n_383),
.C(n_411),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_386),
.A2(n_394),
.B(n_407),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_389),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_387),
.B(n_389),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_403),
.B(n_406),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_402),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_400),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_398),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_404),
.B(n_405),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_412),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_410),
.B(n_412),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_416),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_415),
.C(n_416),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_420),
.B(n_423),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_420),
.B(n_423),
.Y(n_424)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g426 ( 
.A1(n_427),
.A2(n_428),
.B(n_431),
.C(n_432),
.D(n_433),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_438),
.B(n_441),
.Y(n_440)
);

INVx6_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);


endmodule