module fake_jpeg_28724_n_476 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_476);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_476;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_10),
.B(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g56 ( 
.A1(n_31),
.A2(n_16),
.B(n_1),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_56),
.B(n_37),
.C(n_28),
.Y(n_113)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_19),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_58),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_31),
.B(n_16),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_22),
.B(n_16),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_94),
.Y(n_114)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_85),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_22),
.B(n_0),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_91),
.Y(n_117)
);

BUFx4f_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_93),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_47),
.Y(n_123)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_97),
.Y(n_146)
);

BUFx4f_ASAP7_75t_SL g97 ( 
.A(n_18),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_58),
.A2(n_21),
.B1(n_23),
.B2(n_18),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_100),
.A2(n_121),
.B1(n_122),
.B2(n_57),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_113),
.B(n_123),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_86),
.A2(n_21),
.B1(n_23),
.B2(n_18),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_68),
.A2(n_21),
.B1(n_23),
.B2(n_45),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_41),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_140),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_91),
.B(n_0),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_130),
.B(n_150),
.C(n_47),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_63),
.A2(n_26),
.B(n_46),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_136),
.A2(n_39),
.B(n_30),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_35),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_49),
.A2(n_95),
.B1(n_94),
.B2(n_88),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_54),
.B1(n_84),
.B2(n_80),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_52),
.B(n_35),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_149),
.B(n_117),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_60),
.B(n_48),
.C(n_29),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_83),
.A2(n_37),
.B1(n_28),
.B2(n_41),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_145),
.A2(n_29),
.B1(n_33),
.B2(n_30),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_153),
.B(n_188),
.Y(n_250)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_155),
.A2(n_105),
.B1(n_101),
.B2(n_106),
.Y(n_225)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_157),
.B(n_166),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_114),
.A2(n_66),
.B1(n_78),
.B2(n_82),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_158),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_206)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_160),
.A2(n_162),
.B1(n_178),
.B2(n_107),
.Y(n_213)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_59),
.B1(n_70),
.B2(n_65),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_0),
.B(n_2),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_163),
.Y(n_246)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

INVx3_ASAP7_75t_SL g222 ( 
.A(n_164),
.Y(n_222)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_167),
.Y(n_245)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_104),
.A2(n_33),
.B1(n_48),
.B2(n_46),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_170),
.A2(n_190),
.B1(n_133),
.B2(n_119),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_116),
.B(n_39),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_171),
.B(n_186),
.Y(n_226)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_172),
.Y(n_217)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_174),
.Y(n_229)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_175),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_135),
.B(n_23),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_103),
.C(n_124),
.Y(n_212)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_109),
.A2(n_55),
.B1(n_53),
.B2(n_64),
.Y(n_178)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_122),
.A2(n_61),
.B1(n_43),
.B2(n_44),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_108),
.Y(n_182)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_182),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_121),
.A2(n_100),
.B1(n_148),
.B2(n_120),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_120),
.A2(n_47),
.B1(n_45),
.B2(n_44),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_128),
.B(n_47),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_185),
.B(n_196),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_98),
.B(n_23),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_104),
.A2(n_93),
.B1(n_77),
.B2(n_63),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_137),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_195),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_139),
.A2(n_45),
.B1(n_44),
.B2(n_77),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_192),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_241)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_45),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

INVx11_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_115),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_198),
.B(n_200),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_152),
.A2(n_44),
.B1(n_93),
.B2(n_4),
.Y(n_199)
);

OA22x2_ASAP7_75t_L g221 ( 
.A1(n_199),
.A2(n_103),
.B1(n_105),
.B2(n_125),
.Y(n_221)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_132),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_201),
.B(n_204),
.Y(n_224)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_106),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_139),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_203),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_112),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_205),
.B(n_7),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_148),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_208),
.B(n_220),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_211),
.Y(n_257)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_212),
.B(n_9),
.C(n_10),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_213),
.A2(n_231),
.B1(n_232),
.B2(n_168),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_107),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_221),
.Y(n_274)
);

AO22x2_ASAP7_75t_L g223 ( 
.A1(n_174),
.A2(n_133),
.B1(n_124),
.B2(n_119),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_223),
.B(n_15),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_225),
.A2(n_199),
.B1(n_178),
.B2(n_160),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_101),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_161),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_179),
.A2(n_194),
.B1(n_153),
.B2(n_158),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_179),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_163),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_234),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_241),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_243),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_L g247 ( 
.A(n_176),
.B(n_8),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_251),
.A2(n_258),
.B1(n_260),
.B2(n_262),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_249),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_272),
.Y(n_303)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_253),
.Y(n_295)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_254),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_246),
.A2(n_188),
.B1(n_202),
.B2(n_204),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_256),
.B(n_263),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_206),
.A2(n_162),
.B1(n_172),
.B2(n_169),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_221),
.A2(n_197),
.B1(n_167),
.B2(n_156),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_259),
.A2(n_245),
.B1(n_237),
.B2(n_239),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_229),
.A2(n_223),
.B1(n_221),
.B2(n_225),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_261),
.A2(n_241),
.B1(n_227),
.B2(n_238),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_223),
.A2(n_221),
.B1(n_206),
.B2(n_213),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_175),
.B(n_173),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_270),
.Y(n_299)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_207),
.Y(n_265)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_177),
.B1(n_189),
.B2(n_154),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_266),
.A2(n_222),
.B1(n_248),
.B2(n_217),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_250),
.A2(n_164),
.B(n_159),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g325 ( 
.A(n_267),
.B(n_271),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_268),
.B(n_281),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_269),
.A2(n_273),
.B1(n_278),
.B2(n_251),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_208),
.B(n_11),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_207),
.Y(n_271)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_271),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_236),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_240),
.Y(n_275)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_275),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_220),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_230),
.B(n_212),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_282),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_219),
.B(n_215),
.C(n_226),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_235),
.C(n_245),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_234),
.A2(n_13),
.B(n_14),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_223),
.B(n_13),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_210),
.Y(n_283)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_283),
.Y(n_293)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_244),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_288),
.Y(n_294)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_285),
.B(n_287),
.Y(n_316)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_210),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_224),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_214),
.B(n_13),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_242),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_214),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_290),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_291),
.A2(n_298),
.B1(n_300),
.B2(n_304),
.Y(n_334)
);

AO22x1_ASAP7_75t_SL g292 ( 
.A1(n_262),
.A2(n_237),
.B1(n_216),
.B2(n_217),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_292),
.B(n_313),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_235),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_297),
.B(n_302),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_274),
.A2(n_232),
.B1(n_218),
.B2(n_209),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_228),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_268),
.C(n_266),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_280),
.B(n_228),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_274),
.A2(n_218),
.B1(n_209),
.B2(n_222),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_307),
.B(n_320),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_308),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_310),
.A2(n_315),
.B1(n_306),
.B2(n_305),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_311),
.A2(n_309),
.B(n_269),
.Y(n_332)
);

OAI32xp33_ASAP7_75t_L g312 ( 
.A1(n_282),
.A2(n_216),
.A3(n_239),
.B1(n_242),
.B2(n_255),
.Y(n_312)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_312),
.Y(n_330)
);

OA21x2_ASAP7_75t_L g314 ( 
.A1(n_260),
.A2(n_273),
.B(n_259),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_324),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_258),
.A2(n_257),
.B1(n_261),
.B2(n_276),
.Y(n_315)
);

OAI32xp33_ASAP7_75t_L g318 ( 
.A1(n_255),
.A2(n_264),
.A3(n_270),
.B1(n_278),
.B2(n_286),
.Y(n_318)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_256),
.B(n_268),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_267),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_281),
.Y(n_343)
);

OA21x2_ASAP7_75t_L g324 ( 
.A1(n_253),
.A2(n_254),
.B(n_263),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_325),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_327),
.B(n_340),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_301),
.B(n_252),
.C(n_265),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_331),
.B(n_335),
.C(n_351),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_332),
.A2(n_347),
.B(n_352),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_289),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_303),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_336),
.B(n_346),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_309),
.A2(n_306),
.B1(n_314),
.B2(n_292),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_337),
.A2(n_338),
.B1(n_348),
.B2(n_349),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_309),
.A2(n_286),
.B1(n_277),
.B2(n_290),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_295),
.Y(n_341)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_341),
.Y(n_359)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_295),
.Y(n_342)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_343),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_345),
.A2(n_294),
.B1(n_330),
.B2(n_339),
.Y(n_366)
);

AOI322xp5_ASAP7_75t_L g346 ( 
.A1(n_305),
.A2(n_275),
.A3(n_283),
.B1(n_285),
.B2(n_287),
.C1(n_318),
.C2(n_314),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_315),
.A2(n_326),
.B1(n_298),
.B2(n_292),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_310),
.A2(n_312),
.B1(n_325),
.B2(n_319),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_325),
.A2(n_319),
.B1(n_324),
.B2(n_326),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_296),
.Y(n_350)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_350),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_307),
.B(n_299),
.C(n_313),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_324),
.A2(n_303),
.B(n_316),
.Y(n_352)
);

NOR2x1_ASAP7_75t_L g353 ( 
.A(n_296),
.B(n_299),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_357),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_293),
.Y(n_355)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_355),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_317),
.A2(n_321),
.B1(n_322),
.B2(n_293),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_356),
.A2(n_334),
.B1(n_347),
.B2(n_333),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_321),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_322),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_361),
.B(n_365),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_336),
.B(n_353),
.Y(n_364)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_364),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_366),
.A2(n_371),
.B1(n_360),
.B2(n_358),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_370),
.A2(n_354),
.B1(n_383),
.B2(n_369),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_330),
.A2(n_339),
.B1(n_334),
.B2(n_332),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_335),
.B(n_351),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_372),
.B(n_377),
.C(n_329),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_327),
.B(n_331),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_379),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_328),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_375),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_344),
.A2(n_352),
.B(n_349),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_376),
.A2(n_368),
.B(n_370),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_337),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_333),
.Y(n_378)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_378),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_338),
.B(n_344),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_341),
.Y(n_380)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_380),
.Y(n_403)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_342),
.Y(n_382)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_382),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_356),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_383),
.B(n_329),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_350),
.Y(n_384)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_384),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_385),
.B(n_392),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_388),
.B(n_393),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_372),
.B(n_354),
.C(n_365),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_390),
.B(n_400),
.C(n_397),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_391),
.A2(n_406),
.B1(n_401),
.B2(n_405),
.Y(n_424)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_364),
.Y(n_392)
);

XNOR2x1_ASAP7_75t_L g393 ( 
.A(n_361),
.B(n_377),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_378),
.Y(n_394)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_394),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_358),
.A2(n_376),
.B(n_369),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_398),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_381),
.B(n_374),
.C(n_379),
.Y(n_400)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_402),
.Y(n_416)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_359),
.Y(n_404)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_404),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_363),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_387),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_366),
.A2(n_362),
.B1(n_375),
.B2(n_367),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_386),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_408),
.B(n_418),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_395),
.Y(n_409)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_409),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_396),
.A2(n_373),
.B1(n_381),
.B2(n_391),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_412),
.A2(n_424),
.B1(n_389),
.B2(n_404),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_389),
.C(n_403),
.Y(n_426)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_414),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_399),
.C(n_390),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_417),
.C(n_419),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_399),
.B(n_388),
.C(n_393),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_402),
.B(n_395),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_406),
.C(n_385),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_387),
.Y(n_421)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_421),
.Y(n_435)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_394),
.Y(n_423)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_423),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_420),
.B(n_417),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_425),
.B(n_428),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_426),
.B(n_430),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_416),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_429),
.Y(n_439)
);

NAND3xp33_ASAP7_75t_L g430 ( 
.A(n_416),
.B(n_410),
.C(n_408),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_407),
.Y(n_431)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_431),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_419),
.B(n_420),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_432),
.B(n_437),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_413),
.Y(n_437)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_430),
.Y(n_442)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_442),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_429),
.A2(n_407),
.B(n_423),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_447),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_431),
.A2(n_424),
.B1(n_422),
.B2(n_414),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_446),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_SL g445 ( 
.A1(n_436),
.A2(n_422),
.B1(n_421),
.B2(n_415),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_445),
.A2(n_433),
.B(n_427),
.Y(n_452)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_435),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_438),
.B(n_437),
.C(n_432),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_434),
.B(n_438),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_449),
.B(n_447),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_448),
.B(n_425),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_440),
.Y(n_465)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_452),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_441),
.B(n_442),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_453),
.B(n_456),
.Y(n_461)
);

NOR2x1_ASAP7_75t_L g455 ( 
.A(n_448),
.B(n_444),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_455),
.B(n_457),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_450),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_459),
.B(n_446),
.Y(n_460)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_460),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_461),
.B(n_464),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_457),
.B(n_450),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_465),
.B(n_440),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_468),
.B(n_454),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_462),
.A2(n_453),
.B(n_458),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_469),
.A2(n_460),
.B(n_459),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_470),
.B(n_471),
.Y(n_472)
);

BUFx24_ASAP7_75t_SL g473 ( 
.A(n_472),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_473),
.A2(n_467),
.B(n_463),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_474),
.B(n_466),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_475),
.B(n_443),
.Y(n_476)
);


endmodule