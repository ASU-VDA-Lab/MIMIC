module fake_netlist_1_6216_n_1075 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_280, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1075);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1075;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_667;
wire n_496;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_617;
wire n_384;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_303;
wire n_1042;
wire n_1060;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_529;
wire n_312;
wire n_1025;
wire n_1011;
wire n_880;
wire n_630;
wire n_511;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_769;
wire n_844;
wire n_1018;
wire n_738;
wire n_979;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_1046;
wire n_478;
wire n_482;
wire n_415;
wire n_703;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_805;
wire n_729;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_704;
wire n_611;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_601;
wire n_439;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_666;
wire n_423;
wire n_342;
wire n_621;
wire n_799;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_716;
wire n_653;
wire n_899;
wire n_806;
wire n_881;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_955;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_924;
wire n_912;
wire n_947;
wire n_1043;
wire n_582;
wire n_378;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_695;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_992;
INVx1_ASAP7_75t_L g286 ( .A(n_40), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_181), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_234), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_184), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_273), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_106), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_99), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_204), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_38), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_167), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_199), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_178), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_227), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_70), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_16), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_89), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_166), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_76), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_205), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_280), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_255), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_86), .Y(n_307) );
BUFx3_ASAP7_75t_L g308 ( .A(n_190), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_100), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_179), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_146), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_143), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_120), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_27), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_141), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_209), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_176), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_104), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_43), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_256), .Y(n_320) );
CKINVDCx16_ASAP7_75t_R g321 ( .A(n_22), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_66), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_79), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_182), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_172), .Y(n_325) );
CKINVDCx16_ASAP7_75t_R g326 ( .A(n_249), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_284), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_165), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_75), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_57), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_259), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_107), .Y(n_332) );
CKINVDCx16_ASAP7_75t_R g333 ( .A(n_191), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_245), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_260), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_112), .Y(n_336) );
INVx4_ASAP7_75t_R g337 ( .A(n_105), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_116), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_23), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_238), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_196), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_19), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_7), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_220), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_177), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_136), .Y(n_346) );
NOR2xp67_ASAP7_75t_L g347 ( .A(n_189), .B(n_31), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_266), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_281), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_85), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_168), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_212), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_244), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_221), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_110), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_274), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_80), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_92), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_84), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_119), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_67), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_45), .Y(n_362) );
CKINVDCx16_ASAP7_75t_R g363 ( .A(n_113), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_55), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_3), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_66), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_65), .B(n_197), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_77), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_12), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_17), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_203), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_153), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_250), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_265), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_26), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_257), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_228), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_258), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_170), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_242), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_0), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_42), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_222), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_269), .Y(n_384) );
INVxp67_ASAP7_75t_SL g385 ( .A(n_279), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_20), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_124), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_28), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_282), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_152), .Y(n_390) );
INVx1_ASAP7_75t_SL g391 ( .A(n_38), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_186), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_271), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_267), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_98), .Y(n_395) );
CKINVDCx16_ASAP7_75t_R g396 ( .A(n_171), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_37), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_31), .Y(n_398) );
INVxp67_ASAP7_75t_SL g399 ( .A(n_4), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_87), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_188), .Y(n_401) );
INVxp67_ASAP7_75t_L g402 ( .A(n_59), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_233), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_29), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_79), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_51), .Y(n_406) );
CKINVDCx16_ASAP7_75t_R g407 ( .A(n_111), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_4), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_68), .Y(n_409) );
BUFx2_ASAP7_75t_L g410 ( .A(n_251), .Y(n_410) );
CKINVDCx14_ASAP7_75t_R g411 ( .A(n_8), .Y(n_411) );
CKINVDCx16_ASAP7_75t_R g412 ( .A(n_246), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_217), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_210), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_164), .Y(n_415) );
NOR2xp67_ASAP7_75t_L g416 ( .A(n_23), .B(n_175), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_58), .Y(n_417) );
BUFx3_ASAP7_75t_L g418 ( .A(n_232), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_237), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_50), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_17), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_37), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_47), .Y(n_423) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_169), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_103), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_93), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_192), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_121), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_215), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_145), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_56), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_53), .Y(n_432) );
INVxp67_ASAP7_75t_SL g433 ( .A(n_229), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_11), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_150), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_138), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_133), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_127), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_226), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_35), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_69), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_154), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_62), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_326), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_411), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_303), .Y(n_446) );
INVx3_ASAP7_75t_L g447 ( .A(n_290), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_333), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_411), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_303), .Y(n_450) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_328), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_329), .Y(n_452) );
INVx4_ASAP7_75t_L g453 ( .A(n_401), .Y(n_453) );
NOR2xp33_ASAP7_75t_R g454 ( .A(n_363), .B(n_95), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_410), .B(n_0), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_328), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_321), .B(n_1), .Y(n_457) );
OA21x2_ASAP7_75t_L g458 ( .A1(n_290), .A2(n_1), .B(n_2), .Y(n_458) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_328), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_320), .B(n_2), .Y(n_460) );
NOR2xp33_ASAP7_75t_R g461 ( .A(n_396), .B(n_96), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_323), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_328), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_323), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_358), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_338), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_358), .Y(n_467) );
INVx3_ASAP7_75t_L g468 ( .A(n_292), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_394), .B(n_3), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_292), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_388), .Y(n_471) );
BUFx2_ASAP7_75t_L g472 ( .A(n_407), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_338), .Y(n_473) );
OAI22xp5_ASAP7_75t_SL g474 ( .A1(n_314), .A2(n_7), .B1(n_5), .B2(n_6), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_388), .B(n_5), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_408), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_408), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_432), .B(n_6), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_338), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_412), .Y(n_480) );
INVx4_ASAP7_75t_L g481 ( .A(n_308), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_419), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_419), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_453), .B(n_445), .Y(n_484) );
BUFx3_ASAP7_75t_L g485 ( .A(n_475), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_453), .B(n_437), .Y(n_486) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_451), .Y(n_487) );
BUFx3_ASAP7_75t_L g488 ( .A(n_475), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_453), .B(n_432), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_458), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_466), .Y(n_491) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_451), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_458), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_458), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_472), .Y(n_495) );
BUFx10_ASAP7_75t_L g496 ( .A(n_445), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_449), .B(n_441), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_466), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_453), .B(n_441), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_458), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_451), .Y(n_501) );
AND2x2_ASAP7_75t_SL g502 ( .A(n_458), .B(n_367), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_449), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_472), .A2(n_295), .B1(n_324), .B2(n_288), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_466), .Y(n_505) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_472), .A2(n_330), .B1(n_343), .B2(n_329), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_453), .B(n_291), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_458), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_447), .Y(n_509) );
AND2x6_ASAP7_75t_L g510 ( .A(n_475), .B(n_308), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_447), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_447), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_452), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_455), .B(n_330), .Y(n_514) );
INVxp33_ASAP7_75t_L g515 ( .A(n_452), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_451), .Y(n_516) );
AND2x6_ASAP7_75t_L g517 ( .A(n_475), .B(n_353), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_455), .B(n_343), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_447), .Y(n_519) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_451), .Y(n_520) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_451), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_482), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_457), .B(n_361), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_451), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_444), .B(n_293), .Y(n_525) );
INVx4_ASAP7_75t_SL g526 ( .A(n_475), .Y(n_526) );
INVx6_ASAP7_75t_L g527 ( .A(n_481), .Y(n_527) );
BUFx10_ASAP7_75t_L g528 ( .A(n_448), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_447), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_468), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_480), .B(n_297), .Y(n_531) );
AND2x4_ASAP7_75t_L g532 ( .A(n_497), .B(n_455), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_489), .B(n_469), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_495), .B(n_457), .Y(n_534) );
NOR2xp33_ASAP7_75t_SL g535 ( .A(n_502), .B(n_288), .Y(n_535) );
AND2x6_ASAP7_75t_L g536 ( .A(n_485), .B(n_478), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_489), .B(n_478), .Y(n_537) );
AO22x1_ASAP7_75t_L g538 ( .A1(n_504), .A2(n_457), .B1(n_370), .B2(n_375), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_526), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_515), .B(n_460), .Y(n_540) );
NOR2xp33_ASAP7_75t_R g541 ( .A(n_528), .B(n_295), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_514), .B(n_460), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_503), .Y(n_543) );
NOR2xp67_ASAP7_75t_L g544 ( .A(n_513), .B(n_468), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_526), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_489), .B(n_478), .Y(n_546) );
INVx5_ASAP7_75t_L g547 ( .A(n_510), .Y(n_547) );
INVx5_ASAP7_75t_L g548 ( .A(n_510), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_484), .B(n_478), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_489), .B(n_481), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_510), .A2(n_481), .B1(n_470), .B2(n_468), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_486), .B(n_287), .Y(n_552) );
INVx4_ASAP7_75t_L g553 ( .A(n_510), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_499), .B(n_510), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_509), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_509), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_499), .B(n_481), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_511), .Y(n_558) );
INVx5_ASAP7_75t_L g559 ( .A(n_510), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_511), .Y(n_560) );
NOR2x1p5_ASAP7_75t_L g561 ( .A(n_523), .B(n_361), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_510), .A2(n_481), .B1(n_470), .B2(n_468), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_512), .Y(n_563) );
AND2x4_ASAP7_75t_L g564 ( .A(n_499), .B(n_446), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_518), .A2(n_474), .B1(n_375), .B2(n_404), .Y(n_565) );
INVx3_ASAP7_75t_L g566 ( .A(n_488), .Y(n_566) );
OAI22xp5_ASAP7_75t_SL g567 ( .A1(n_523), .A2(n_474), .B1(n_314), .B2(n_397), .Y(n_567) );
AND2x4_ASAP7_75t_L g568 ( .A(n_499), .B(n_446), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_517), .A2(n_470), .B1(n_468), .B2(n_286), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_519), .Y(n_570) );
INVxp67_ASAP7_75t_L g571 ( .A(n_496), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_488), .Y(n_572) );
OR2x6_ASAP7_75t_L g573 ( .A(n_528), .B(n_402), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_525), .B(n_454), .Y(n_574) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_502), .Y(n_575) );
BUFx3_ASAP7_75t_L g576 ( .A(n_528), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_531), .B(n_461), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_506), .B(n_461), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_517), .B(n_507), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_517), .B(n_470), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_517), .B(n_470), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_517), .B(n_502), .Y(n_582) );
INVx3_ASAP7_75t_L g583 ( .A(n_517), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_528), .Y(n_584) );
BUFx8_ASAP7_75t_L g585 ( .A(n_517), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_490), .B(n_287), .Y(n_586) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_490), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_493), .B(n_289), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_494), .B(n_289), .Y(n_589) );
INVx2_ASAP7_75t_SL g590 ( .A(n_494), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_529), .B(n_370), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_529), .Y(n_592) );
INVxp67_ASAP7_75t_L g593 ( .A(n_530), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_500), .B(n_450), .Y(n_594) );
INVxp67_ASAP7_75t_L g595 ( .A(n_530), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_508), .A2(n_406), .B1(n_421), .B2(n_404), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_508), .A2(n_421), .B1(n_423), .B2(n_406), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_527), .B(n_296), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_527), .A2(n_443), .B1(n_423), .B2(n_342), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_527), .A2(n_397), .B1(n_322), .B2(n_294), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_491), .A2(n_299), .B1(n_307), .B2(n_301), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_491), .B(n_296), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_498), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_498), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_505), .B(n_304), .Y(n_605) );
AND2x6_ASAP7_75t_SL g606 ( .A(n_522), .B(n_319), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_501), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_541), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_566), .Y(n_609) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_587), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_543), .B(n_339), .Y(n_611) );
AO22x1_ASAP7_75t_L g612 ( .A1(n_585), .A2(n_316), .B1(n_318), .B2(n_304), .Y(n_612) );
INVx4_ASAP7_75t_L g613 ( .A(n_573), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_564), .Y(n_614) );
INVx5_ASAP7_75t_L g615 ( .A(n_573), .Y(n_615) );
O2A1O1Ixp33_ASAP7_75t_L g616 ( .A1(n_533), .A2(n_399), .B(n_350), .C(n_359), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_533), .B(n_532), .Y(n_617) );
INVxp33_ASAP7_75t_L g618 ( .A(n_534), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_590), .A2(n_524), .B(n_516), .Y(n_619) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_587), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g621 ( .A1(n_537), .A2(n_362), .B(n_364), .C(n_357), .Y(n_621) );
O2A1O1Ixp33_ASAP7_75t_L g622 ( .A1(n_537), .A2(n_546), .B(n_578), .C(n_600), .Y(n_622) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_587), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_535), .A2(n_424), .B1(n_433), .B2(n_385), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_566), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_532), .B(n_300), .Y(n_626) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_553), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_564), .Y(n_628) );
AND2x4_ASAP7_75t_L g629 ( .A(n_576), .B(n_365), .Y(n_629) );
INVx1_ASAP7_75t_SL g630 ( .A(n_554), .Y(n_630) );
BUFx3_ASAP7_75t_L g631 ( .A(n_584), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_591), .B(n_327), .Y(n_632) );
INVx5_ASAP7_75t_L g633 ( .A(n_536), .Y(n_633) );
BUFx12f_ASAP7_75t_L g634 ( .A(n_606), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_575), .A2(n_349), .B1(n_356), .B2(n_332), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_546), .A2(n_368), .B(n_369), .C(n_366), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_600), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_540), .B(n_391), .Y(n_638) );
OR2x6_ASAP7_75t_L g639 ( .A(n_538), .B(n_381), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_568), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_594), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_586), .A2(n_589), .B(n_588), .Y(n_642) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_547), .Y(n_643) );
INVx5_ASAP7_75t_L g644 ( .A(n_536), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_571), .B(n_371), .Y(n_645) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_544), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_550), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_586), .A2(n_524), .B(n_516), .Y(n_648) );
INVx4_ASAP7_75t_L g649 ( .A(n_547), .Y(n_649) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_567), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_542), .B(n_382), .Y(n_651) );
INVxp67_ASAP7_75t_L g652 ( .A(n_561), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g653 ( .A1(n_549), .A2(n_386), .B(n_400), .C(n_398), .Y(n_653) );
BUFx2_ASAP7_75t_L g654 ( .A(n_585), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_596), .B(n_373), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_550), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_597), .B(n_373), .Y(n_657) );
BUFx8_ASAP7_75t_L g658 ( .A(n_536), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_580), .Y(n_659) );
AOI222xp33_ASAP7_75t_L g660 ( .A1(n_535), .A2(n_465), .B1(n_462), .B2(n_467), .C1(n_464), .C2(n_450), .Y(n_660) );
A2O1A1Ixp33_ASAP7_75t_L g661 ( .A1(n_589), .A2(n_405), .B(n_417), .C(n_409), .Y(n_661) );
INVx1_ASAP7_75t_SL g662 ( .A(n_580), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_557), .Y(n_663) );
AO22x1_ASAP7_75t_L g664 ( .A1(n_536), .A2(n_374), .B1(n_413), .B2(n_376), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_582), .A2(n_524), .B(n_302), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_555), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_579), .A2(n_422), .B1(n_426), .B2(n_420), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_556), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_574), .B(n_431), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_582), .A2(n_305), .B(n_298), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_558), .Y(n_671) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_581), .Y(n_672) );
BUFx12f_ASAP7_75t_L g673 ( .A(n_547), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_595), .A2(n_309), .B(n_306), .Y(n_674) );
AOI222xp33_ASAP7_75t_L g675 ( .A1(n_601), .A2(n_465), .B1(n_477), .B2(n_471), .C1(n_462), .C2(n_464), .Y(n_675) );
BUFx2_ASAP7_75t_L g676 ( .A(n_579), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g677 ( .A1(n_581), .A2(n_440), .B(n_434), .C(n_467), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_565), .A2(n_311), .B1(n_312), .B2(n_310), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_560), .Y(n_679) );
AND2x4_ASAP7_75t_L g680 ( .A(n_548), .B(n_471), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_599), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_572), .Y(n_682) );
AO22x1_ASAP7_75t_L g683 ( .A1(n_548), .A2(n_374), .B1(n_413), .B2(n_376), .Y(n_683) );
INVxp67_ASAP7_75t_L g684 ( .A(n_602), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_569), .A2(n_315), .B1(n_317), .B2(n_313), .Y(n_685) );
BUFx6f_ASAP7_75t_L g686 ( .A(n_548), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_563), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g688 ( .A1(n_552), .A2(n_415), .B1(n_427), .B2(n_414), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_577), .B(n_415), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g690 ( .A1(n_570), .A2(n_416), .B(n_347), .C(n_476), .Y(n_690) );
CKINVDCx5p33_ASAP7_75t_R g691 ( .A(n_605), .Y(n_691) );
O2A1O1Ixp33_ASAP7_75t_L g692 ( .A1(n_605), .A2(n_477), .B(n_331), .C(n_335), .Y(n_692) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_559), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_593), .B(n_551), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_592), .Y(n_695) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_559), .Y(n_696) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_559), .Y(n_697) );
A2O1A1Ixp33_ASAP7_75t_L g698 ( .A1(n_562), .A2(n_334), .B(n_341), .C(n_336), .Y(n_698) );
INVxp67_ASAP7_75t_SL g699 ( .A(n_583), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_598), .B(n_427), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_539), .A2(n_345), .B1(n_346), .B2(n_344), .Y(n_701) );
BUFx2_ASAP7_75t_SL g702 ( .A(n_545), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_603), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_604), .A2(n_351), .B1(n_352), .B2(n_348), .Y(n_704) );
BUFx6f_ASAP7_75t_L g705 ( .A(n_607), .Y(n_705) );
OR2x6_ASAP7_75t_L g706 ( .A(n_573), .B(n_354), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_566), .Y(n_707) );
O2A1O1Ixp33_ASAP7_75t_L g708 ( .A1(n_533), .A2(n_372), .B(n_377), .C(n_360), .Y(n_708) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_587), .Y(n_709) );
NAND2xp33_ASAP7_75t_L g710 ( .A(n_587), .B(n_419), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_535), .A2(n_379), .B1(n_387), .B2(n_378), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_575), .A2(n_390), .B1(n_392), .B2(n_389), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_543), .B(n_393), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_566), .Y(n_714) );
BUFx12f_ASAP7_75t_L g715 ( .A(n_573), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_534), .B(n_8), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_617), .B(n_428), .Y(n_717) );
INVxp67_ASAP7_75t_SL g718 ( .A(n_610), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_637), .A2(n_380), .B1(n_418), .B2(n_353), .Y(n_719) );
OAI21x1_ASAP7_75t_L g720 ( .A1(n_648), .A2(n_340), .B(n_325), .Y(n_720) );
CKINVDCx11_ASAP7_75t_R g721 ( .A(n_715), .Y(n_721) );
CKINVDCx16_ASAP7_75t_R g722 ( .A(n_706), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_618), .B(n_9), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g724 ( .A1(n_642), .A2(n_430), .B(n_429), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_660), .A2(n_436), .B1(n_438), .B2(n_435), .Y(n_725) );
AOI21x1_ASAP7_75t_L g726 ( .A1(n_670), .A2(n_383), .B(n_355), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_716), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g728 ( .A(n_610), .B(n_439), .Y(n_728) );
NAND2x1p5_ASAP7_75t_L g729 ( .A(n_633), .B(n_380), .Y(n_729) );
OAI21x1_ASAP7_75t_L g730 ( .A1(n_619), .A2(n_384), .B(n_383), .Y(n_730) );
AO21x2_ASAP7_75t_L g731 ( .A1(n_690), .A2(n_395), .B(n_384), .Y(n_731) );
AO21x2_ASAP7_75t_L g732 ( .A1(n_711), .A2(n_425), .B(n_403), .Y(n_732) );
NAND2xp33_ASAP7_75t_L g733 ( .A(n_610), .B(n_419), .Y(n_733) );
OA21x2_ASAP7_75t_L g734 ( .A1(n_665), .A2(n_442), .B(n_456), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_626), .B(n_9), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_706), .B(n_10), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_674), .A2(n_463), .B(n_456), .Y(n_737) );
AND2x4_ASAP7_75t_L g738 ( .A(n_615), .B(n_10), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_647), .B(n_11), .Y(n_739) );
OA21x2_ASAP7_75t_L g740 ( .A1(n_661), .A2(n_463), .B(n_456), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_666), .Y(n_741) );
INVx3_ASAP7_75t_L g742 ( .A(n_673), .Y(n_742) );
O2A1O1Ixp33_ASAP7_75t_L g743 ( .A1(n_653), .A2(n_482), .B(n_463), .C(n_473), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_691), .B(n_13), .Y(n_744) );
INVx3_ASAP7_75t_SL g745 ( .A(n_706), .Y(n_745) );
INVx8_ASAP7_75t_L g746 ( .A(n_633), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_668), .Y(n_747) );
NOR2xp67_ASAP7_75t_SL g748 ( .A(n_613), .B(n_337), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_671), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_624), .A2(n_483), .B1(n_479), .B2(n_482), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_681), .A2(n_483), .B1(n_479), .B2(n_459), .Y(n_751) );
AOI21x1_ASAP7_75t_L g752 ( .A1(n_679), .A2(n_459), .B(n_451), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_641), .A2(n_459), .B1(n_492), .B2(n_487), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_695), .Y(n_754) );
OAI21xp5_ASAP7_75t_L g755 ( .A1(n_622), .A2(n_459), .B(n_13), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_656), .B(n_14), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_704), .A2(n_459), .B1(n_492), .B2(n_487), .Y(n_757) );
AND2x4_ASAP7_75t_L g758 ( .A(n_613), .B(n_14), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_687), .Y(n_759) );
BUFx3_ASAP7_75t_L g760 ( .A(n_631), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_704), .A2(n_459), .B1(n_492), .B2(n_487), .Y(n_761) );
NAND2x1p5_ASAP7_75t_L g762 ( .A(n_633), .B(n_15), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_703), .Y(n_763) );
OA21x2_ASAP7_75t_L g764 ( .A1(n_698), .A2(n_521), .B(n_520), .Y(n_764) );
INVx3_ASAP7_75t_L g765 ( .A(n_644), .Y(n_765) );
NAND4xp25_ASAP7_75t_L g766 ( .A(n_678), .B(n_18), .C(n_15), .D(n_16), .Y(n_766) );
NAND2xp5_ASAP7_75t_SL g767 ( .A(n_620), .B(n_492), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_614), .Y(n_768) );
AO21x1_ASAP7_75t_L g769 ( .A1(n_692), .A2(n_101), .B(n_97), .Y(n_769) );
AND2x6_ASAP7_75t_L g770 ( .A(n_627), .B(n_520), .Y(n_770) );
AND2x4_ASAP7_75t_L g771 ( .A(n_644), .B(n_20), .Y(n_771) );
OAI21x1_ASAP7_75t_L g772 ( .A1(n_682), .A2(n_521), .B(n_108), .Y(n_772) );
NAND3xp33_ASAP7_75t_L g773 ( .A(n_688), .B(n_521), .C(n_21), .Y(n_773) );
BUFx2_ASAP7_75t_SL g774 ( .A(n_644), .Y(n_774) );
OA21x2_ASAP7_75t_L g775 ( .A1(n_694), .A2(n_109), .B(n_102), .Y(n_775) );
BUFx3_ASAP7_75t_L g776 ( .A(n_658), .Y(n_776) );
OAI21x1_ASAP7_75t_L g777 ( .A1(n_609), .A2(n_115), .B(n_114), .Y(n_777) );
AO31x2_ASAP7_75t_L g778 ( .A1(n_669), .A2(n_24), .A3(n_21), .B(n_22), .Y(n_778) );
OAI21xp5_ASAP7_75t_L g779 ( .A1(n_684), .A2(n_24), .B(n_25), .Y(n_779) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_663), .A2(n_27), .B1(n_25), .B2(n_26), .Y(n_780) );
INVx4_ASAP7_75t_L g781 ( .A(n_639), .Y(n_781) );
OAI21x1_ASAP7_75t_L g782 ( .A1(n_625), .A2(n_118), .B(n_117), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_611), .A2(n_28), .B1(n_29), .B2(n_30), .Y(n_783) );
OAI22xp33_ASAP7_75t_L g784 ( .A1(n_639), .A2(n_32), .B1(n_33), .B2(n_34), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_628), .Y(n_785) );
AND2x4_ASAP7_75t_L g786 ( .A(n_654), .B(n_34), .Y(n_786) );
OAI21x1_ASAP7_75t_L g787 ( .A1(n_707), .A2(n_123), .B(n_122), .Y(n_787) );
INVx3_ASAP7_75t_L g788 ( .A(n_627), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_705), .Y(n_789) );
AO21x2_ASAP7_75t_L g790 ( .A1(n_708), .A2(n_126), .B(n_125), .Y(n_790) );
OAI21x1_ASAP7_75t_L g791 ( .A1(n_714), .A2(n_129), .B(n_128), .Y(n_791) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_634), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_640), .Y(n_793) );
OAI21x1_ASAP7_75t_L g794 ( .A1(n_677), .A2(n_131), .B(n_130), .Y(n_794) );
OAI22xp33_ASAP7_75t_L g795 ( .A1(n_678), .A2(n_36), .B1(n_39), .B2(n_40), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_630), .B(n_39), .Y(n_796) );
OAI21x1_ASAP7_75t_L g797 ( .A1(n_701), .A2(n_636), .B(n_621), .Y(n_797) );
OA21x2_ASAP7_75t_L g798 ( .A1(n_712), .A2(n_134), .B(n_132), .Y(n_798) );
CKINVDCx6p67_ASAP7_75t_R g799 ( .A(n_629), .Y(n_799) );
AO221x2_ASAP7_75t_L g800 ( .A1(n_664), .A2(n_41), .B1(n_42), .B2(n_43), .C(n_44), .Y(n_800) );
OAI21x1_ASAP7_75t_L g801 ( .A1(n_693), .A2(n_700), .B(n_699), .Y(n_801) );
NAND2xp33_ASAP7_75t_L g802 ( .A(n_620), .B(n_135), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_651), .A2(n_46), .B1(n_47), .B2(n_48), .Y(n_803) );
OAI21x1_ASAP7_75t_L g804 ( .A1(n_616), .A2(n_139), .B(n_137), .Y(n_804) );
AND2x2_ASAP7_75t_SL g805 ( .A(n_620), .B(n_46), .Y(n_805) );
NOR2xp33_ASAP7_75t_R g806 ( .A(n_608), .B(n_48), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_675), .Y(n_807) );
A2O1A1Ixp33_ASAP7_75t_L g808 ( .A1(n_713), .A2(n_49), .B(n_50), .C(n_51), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_646), .Y(n_809) );
OAI21x1_ASAP7_75t_L g810 ( .A1(n_667), .A2(n_142), .B(n_140), .Y(n_810) );
NAND2x1_ASAP7_75t_L g811 ( .A(n_649), .B(n_144), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_659), .B(n_49), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_662), .B(n_52), .Y(n_813) );
OAI21x1_ASAP7_75t_L g814 ( .A1(n_685), .A2(n_148), .B(n_147), .Y(n_814) );
INVxp67_ASAP7_75t_L g815 ( .A(n_672), .Y(n_815) );
AND2x4_ASAP7_75t_L g816 ( .A(n_676), .B(n_52), .Y(n_816) );
INVx4_ASAP7_75t_L g817 ( .A(n_623), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_632), .Y(n_818) );
OAI21x1_ASAP7_75t_L g819 ( .A1(n_645), .A2(n_151), .B(n_149), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_652), .B(n_54), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_635), .A2(n_54), .B1(n_55), .B2(n_56), .Y(n_821) );
AOI21xp5_ASAP7_75t_L g822 ( .A1(n_710), .A2(n_156), .B(n_155), .Y(n_822) );
OAI21x1_ASAP7_75t_SL g823 ( .A1(n_649), .A2(n_57), .B(n_58), .Y(n_823) );
OAI21xp5_ASAP7_75t_L g824 ( .A1(n_655), .A2(n_59), .B(n_60), .Y(n_824) );
OAI21x1_ASAP7_75t_L g825 ( .A1(n_623), .A2(n_158), .B(n_157), .Y(n_825) );
BUFx6f_ASAP7_75t_L g826 ( .A(n_623), .Y(n_826) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_650), .Y(n_827) );
AOI21xp5_ASAP7_75t_L g828 ( .A1(n_709), .A2(n_160), .B(n_159), .Y(n_828) );
OAI21xp5_ASAP7_75t_L g829 ( .A1(n_657), .A2(n_60), .B(n_61), .Y(n_829) );
OAI21x1_ASAP7_75t_L g830 ( .A1(n_709), .A2(n_162), .B(n_161), .Y(n_830) );
OAI21x1_ASAP7_75t_L g831 ( .A1(n_689), .A2(n_187), .B(n_283), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_680), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_680), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_683), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_702), .Y(n_835) );
AND2x2_ASAP7_75t_L g836 ( .A(n_612), .B(n_63), .Y(n_836) );
AOI222xp33_ASAP7_75t_L g837 ( .A1(n_807), .A2(n_697), .B1(n_696), .B2(n_686), .C1(n_643), .C2(n_68), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_722), .A2(n_697), .B1(n_696), .B2(n_686), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_805), .A2(n_697), .B1(n_696), .B2(n_686), .Y(n_839) );
BUFx12f_ASAP7_75t_L g840 ( .A(n_721), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_759), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_741), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_747), .Y(n_843) );
INVx2_ASAP7_75t_L g844 ( .A(n_763), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_749), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_754), .Y(n_846) );
AOI21xp5_ASAP7_75t_L g847 ( .A1(n_724), .A2(n_185), .B(n_278), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_745), .B(n_64), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_768), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_744), .A2(n_816), .B1(n_818), .B2(n_766), .Y(n_850) );
AOI21xp5_ASAP7_75t_L g851 ( .A1(n_724), .A2(n_183), .B(n_277), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_780), .Y(n_852) );
INVx4_ASAP7_75t_L g853 ( .A(n_746), .Y(n_853) );
OA21x2_ASAP7_75t_L g854 ( .A1(n_720), .A2(n_193), .B(n_276), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_725), .A2(n_71), .B1(n_72), .B2(n_73), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_744), .A2(n_72), .B1(n_73), .B2(n_74), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_780), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_816), .A2(n_74), .B1(n_75), .B2(n_76), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_725), .A2(n_77), .B1(n_78), .B2(n_80), .Y(n_859) );
AOI22xp33_ASAP7_75t_SL g860 ( .A1(n_781), .A2(n_78), .B1(n_81), .B2(n_82), .Y(n_860) );
AND2x4_ASAP7_75t_SL g861 ( .A(n_799), .B(n_81), .Y(n_861) );
OAI21xp5_ASAP7_75t_L g862 ( .A1(n_739), .A2(n_82), .B(n_83), .Y(n_862) );
AND2x4_ASAP7_75t_L g863 ( .A(n_776), .B(n_83), .Y(n_863) );
AOI221xp5_ASAP7_75t_L g864 ( .A1(n_727), .A2(n_87), .B1(n_88), .B2(n_89), .C(n_90), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_800), .A2(n_88), .B1(n_90), .B2(n_91), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_815), .B(n_91), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_800), .A2(n_93), .B1(n_94), .B2(n_163), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_739), .Y(n_868) );
OA21x2_ASAP7_75t_L g869 ( .A1(n_730), .A2(n_173), .B(n_174), .Y(n_869) );
BUFx6f_ASAP7_75t_L g870 ( .A(n_826), .Y(n_870) );
AND2x4_ASAP7_75t_L g871 ( .A(n_776), .B(n_180), .Y(n_871) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_762), .A2(n_194), .B1(n_195), .B2(n_198), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_762), .A2(n_200), .B1(n_201), .B2(n_202), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_756), .A2(n_206), .B1(n_207), .B2(n_208), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_785), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_800), .A2(n_211), .B1(n_213), .B2(n_214), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_735), .A2(n_216), .B1(n_218), .B2(n_219), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_717), .B(n_223), .Y(n_878) );
BUFx5_ASAP7_75t_L g879 ( .A(n_770), .Y(n_879) );
AOI221xp5_ASAP7_75t_L g880 ( .A1(n_795), .A2(n_224), .B1(n_225), .B2(n_230), .C(n_231), .Y(n_880) );
AOI221xp5_ASAP7_75t_L g881 ( .A1(n_820), .A2(n_235), .B1(n_236), .B2(n_239), .C(n_240), .Y(n_881) );
AND2x4_ASAP7_75t_L g882 ( .A(n_815), .B(n_241), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_723), .A2(n_243), .B1(n_247), .B2(n_248), .Y(n_883) );
A2O1A1Ixp33_ASAP7_75t_L g884 ( .A1(n_779), .A2(n_252), .B(n_253), .C(n_254), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_793), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_786), .A2(n_261), .B1(n_262), .B2(n_263), .Y(n_886) );
AOI211xp5_ASAP7_75t_SL g887 ( .A1(n_784), .A2(n_264), .B(n_268), .C(n_270), .Y(n_887) );
OA21x2_ASAP7_75t_L g888 ( .A1(n_772), .A2(n_272), .B(n_275), .Y(n_888) );
INVx6_ASAP7_75t_L g889 ( .A(n_760), .Y(n_889) );
OAI211xp5_ASAP7_75t_L g890 ( .A1(n_806), .A2(n_285), .B(n_783), .C(n_803), .Y(n_890) );
AOI21xp5_ASAP7_75t_L g891 ( .A1(n_767), .A2(n_734), .B(n_801), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_834), .A2(n_736), .B1(n_836), .B2(n_738), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_758), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_758), .Y(n_894) );
AOI21xp5_ASAP7_75t_L g895 ( .A1(n_734), .A2(n_718), .B(n_728), .Y(n_895) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_771), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_812), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_835), .B(n_809), .Y(n_898) );
AND2x4_ASAP7_75t_L g899 ( .A(n_832), .B(n_833), .Y(n_899) );
XOR2xp5_ASAP7_75t_L g900 ( .A(n_792), .B(n_827), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_813), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_813), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_750), .A2(n_731), .B1(n_797), .B2(n_773), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_731), .A2(n_829), .B1(n_824), .B2(n_732), .Y(n_904) );
BUFx12f_ASAP7_75t_L g905 ( .A(n_721), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_796), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_719), .A2(n_742), .B1(n_748), .B2(n_740), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_808), .B(n_778), .Y(n_908) );
AO21x2_ASAP7_75t_L g909 ( .A1(n_769), .A2(n_726), .B(n_790), .Y(n_909) );
INVx3_ASAP7_75t_L g910 ( .A(n_746), .Y(n_910) );
OAI22xp33_ASAP7_75t_L g911 ( .A1(n_821), .A2(n_746), .B1(n_729), .B2(n_765), .Y(n_911) );
AOI22xp33_ASAP7_75t_SL g912 ( .A1(n_823), .A2(n_774), .B1(n_761), .B2(n_757), .Y(n_912) );
OAI22xp33_ASAP7_75t_L g913 ( .A1(n_765), .A2(n_798), .B1(n_728), .B2(n_811), .Y(n_913) );
AND2x2_ASAP7_75t_L g914 ( .A(n_778), .B(n_788), .Y(n_914) );
OAI221xp5_ASAP7_75t_L g915 ( .A1(n_743), .A2(n_751), .B1(n_737), .B2(n_798), .C(n_802), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_778), .B(n_789), .Y(n_916) );
OAI221xp5_ASAP7_75t_L g917 ( .A1(n_737), .A2(n_802), .B1(n_753), .B2(n_828), .C(n_764), .Y(n_917) );
INVx2_ASAP7_75t_SL g918 ( .A(n_817), .Y(n_918) );
OA21x2_ASAP7_75t_L g919 ( .A1(n_777), .A2(n_791), .B(n_787), .Y(n_919) );
AOI21xp5_ASAP7_75t_L g920 ( .A1(n_775), .A2(n_733), .B(n_753), .Y(n_920) );
A2O1A1Ixp33_ASAP7_75t_L g921 ( .A1(n_804), .A2(n_814), .B(n_794), .C(n_810), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_819), .Y(n_922) );
AO21x2_ASAP7_75t_L g923 ( .A1(n_752), .A2(n_782), .B(n_831), .Y(n_923) );
INVx4_ASAP7_75t_L g924 ( .A(n_770), .Y(n_924) );
INVx4_ASAP7_75t_SL g925 ( .A(n_770), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_770), .B(n_826), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_825), .Y(n_927) );
INVx4_ASAP7_75t_SL g928 ( .A(n_830), .Y(n_928) );
OAI21xp5_ASAP7_75t_L g929 ( .A1(n_822), .A2(n_755), .B(n_642), .Y(n_929) );
INVx2_ASAP7_75t_L g930 ( .A(n_759), .Y(n_930) );
INVx2_ASAP7_75t_L g931 ( .A(n_759), .Y(n_931) );
AOI221xp5_ASAP7_75t_L g932 ( .A1(n_818), .A2(n_651), .B1(n_618), .B2(n_638), .C(n_600), .Y(n_932) );
OR2x2_ASAP7_75t_L g933 ( .A(n_852), .B(n_857), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_841), .B(n_844), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_932), .B(n_850), .Y(n_935) );
INVx4_ASAP7_75t_L g936 ( .A(n_925), .Y(n_936) );
BUFx2_ASAP7_75t_L g937 ( .A(n_879), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_930), .B(n_931), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_908), .B(n_868), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_842), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_843), .Y(n_941) );
INVx2_ASAP7_75t_L g942 ( .A(n_927), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_845), .B(n_846), .Y(n_943) );
AND2x2_ASAP7_75t_L g944 ( .A(n_897), .B(n_901), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_902), .B(n_849), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_875), .B(n_885), .Y(n_946) );
NOR2xp33_ASAP7_75t_L g947 ( .A(n_893), .B(n_894), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_906), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_862), .B(n_837), .Y(n_949) );
OR2x2_ASAP7_75t_L g950 ( .A(n_892), .B(n_896), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_914), .Y(n_951) );
BUFx2_ASAP7_75t_L g952 ( .A(n_879), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_916), .Y(n_953) );
HB1xp67_ASAP7_75t_L g954 ( .A(n_882), .Y(n_954) );
INVx3_ASAP7_75t_L g955 ( .A(n_924), .Y(n_955) );
NAND2xp5_ASAP7_75t_SL g956 ( .A(n_839), .B(n_871), .Y(n_956) );
INVx2_ASAP7_75t_L g957 ( .A(n_922), .Y(n_957) );
OAI221xp5_ASAP7_75t_L g958 ( .A1(n_865), .A2(n_867), .B1(n_890), .B2(n_858), .C(n_912), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_870), .Y(n_959) );
INVx2_ASAP7_75t_L g960 ( .A(n_870), .Y(n_960) );
OR2x2_ASAP7_75t_L g961 ( .A(n_839), .B(n_898), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_899), .B(n_855), .Y(n_962) );
BUFx2_ASAP7_75t_SL g963 ( .A(n_853), .Y(n_963) );
AOI222xp33_ASAP7_75t_L g964 ( .A1(n_855), .A2(n_859), .B1(n_861), .B2(n_840), .C1(n_905), .C2(n_863), .Y(n_964) );
INVx2_ASAP7_75t_L g965 ( .A(n_923), .Y(n_965) );
AND2x4_ASAP7_75t_L g966 ( .A(n_925), .B(n_926), .Y(n_966) );
INVx2_ASAP7_75t_L g967 ( .A(n_923), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_887), .B(n_918), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_887), .B(n_904), .Y(n_969) );
INVxp67_ASAP7_75t_L g970 ( .A(n_848), .Y(n_970) );
INVx2_ASAP7_75t_L g971 ( .A(n_919), .Y(n_971) );
AOI21xp33_ASAP7_75t_SL g972 ( .A1(n_872), .A2(n_873), .B(n_911), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_854), .Y(n_973) );
AND2x4_ASAP7_75t_L g974 ( .A(n_925), .B(n_928), .Y(n_974) );
BUFx2_ASAP7_75t_L g975 ( .A(n_879), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_854), .Y(n_976) );
INVx2_ASAP7_75t_L g977 ( .A(n_909), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_866), .B(n_910), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_856), .B(n_864), .Y(n_979) );
OR2x2_ASAP7_75t_L g980 ( .A(n_838), .B(n_907), .Y(n_980) );
AO21x2_ASAP7_75t_L g981 ( .A1(n_929), .A2(n_891), .B(n_920), .Y(n_981) );
INVx2_ASAP7_75t_L g982 ( .A(n_888), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_876), .B(n_860), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_895), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_889), .B(n_903), .Y(n_985) );
AND2x4_ASAP7_75t_L g986 ( .A(n_928), .B(n_929), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_878), .B(n_880), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_869), .Y(n_988) );
INVx2_ASAP7_75t_L g989 ( .A(n_928), .Y(n_989) );
INVx2_ASAP7_75t_L g990 ( .A(n_917), .Y(n_990) );
AND2x4_ASAP7_75t_L g991 ( .A(n_921), .B(n_884), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_874), .B(n_886), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_939), .B(n_874), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_943), .Y(n_994) );
INVx1_ASAP7_75t_SL g995 ( .A(n_963), .Y(n_995) );
AOI221xp5_ASAP7_75t_L g996 ( .A1(n_935), .A2(n_881), .B1(n_915), .B2(n_913), .C(n_900), .Y(n_996) );
AO21x2_ASAP7_75t_L g997 ( .A1(n_973), .A2(n_847), .B(n_851), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_939), .B(n_877), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_933), .Y(n_999) );
OR2x2_ASAP7_75t_L g1000 ( .A(n_953), .B(n_883), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_953), .B(n_951), .Y(n_1001) );
BUFx2_ASAP7_75t_L g1002 ( .A(n_937), .Y(n_1002) );
AND2x4_ASAP7_75t_L g1003 ( .A(n_974), .B(n_966), .Y(n_1003) );
INVx4_ASAP7_75t_L g1004 ( .A(n_936), .Y(n_1004) );
INVxp67_ASAP7_75t_L g1005 ( .A(n_963), .Y(n_1005) );
HB1xp67_ASAP7_75t_L g1006 ( .A(n_946), .Y(n_1006) );
NAND3xp33_ASAP7_75t_L g1007 ( .A(n_964), .B(n_972), .C(n_985), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_942), .Y(n_1008) );
AOI33xp33_ASAP7_75t_L g1009 ( .A1(n_944), .A2(n_940), .A3(n_941), .B1(n_949), .B2(n_948), .B3(n_945), .Y(n_1009) );
OAI221xp5_ASAP7_75t_L g1010 ( .A1(n_970), .A2(n_958), .B1(n_978), .B2(n_979), .C(n_954), .Y(n_1010) );
BUFx2_ASAP7_75t_L g1011 ( .A(n_937), .Y(n_1011) );
OR2x6_ASAP7_75t_L g1012 ( .A(n_956), .B(n_974), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_957), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_934), .B(n_938), .Y(n_1014) );
NAND3xp33_ASAP7_75t_L g1015 ( .A(n_947), .B(n_983), .C(n_968), .Y(n_1015) );
HB1xp67_ASAP7_75t_L g1016 ( .A(n_961), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_990), .B(n_969), .Y(n_1017) );
OR2x2_ASAP7_75t_L g1018 ( .A(n_950), .B(n_962), .Y(n_1018) );
AND2x4_ASAP7_75t_L g1019 ( .A(n_974), .B(n_966), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_992), .B(n_980), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_990), .B(n_986), .Y(n_1021) );
AND2x4_ASAP7_75t_L g1022 ( .A(n_1003), .B(n_986), .Y(n_1022) );
INVx1_ASAP7_75t_SL g1023 ( .A(n_995), .Y(n_1023) );
AND2x4_ASAP7_75t_L g1024 ( .A(n_1003), .B(n_986), .Y(n_1024) );
NAND4xp25_ASAP7_75t_L g1025 ( .A(n_1007), .B(n_986), .C(n_987), .D(n_991), .Y(n_1025) );
AND2x4_ASAP7_75t_L g1026 ( .A(n_1003), .B(n_989), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_994), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_1006), .B(n_960), .Y(n_1028) );
O2A1O1Ixp33_ASAP7_75t_L g1029 ( .A1(n_1010), .A2(n_965), .B(n_967), .C(n_984), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_1021), .B(n_967), .Y(n_1030) );
OR2x2_ASAP7_75t_L g1031 ( .A(n_1018), .B(n_967), .Y(n_1031) );
AND2x4_ASAP7_75t_L g1032 ( .A(n_1019), .B(n_989), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_1001), .B(n_965), .Y(n_1033) );
INVx3_ASAP7_75t_L g1034 ( .A(n_1004), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_1001), .B(n_965), .Y(n_1035) );
AOI31xp33_ASAP7_75t_L g1036 ( .A1(n_1005), .A2(n_989), .A3(n_991), .B(n_936), .Y(n_1036) );
OR2x2_ASAP7_75t_L g1037 ( .A(n_1016), .B(n_981), .Y(n_1037) );
NAND2x1p5_ASAP7_75t_L g1038 ( .A(n_1004), .B(n_936), .Y(n_1038) );
AND2x4_ASAP7_75t_L g1039 ( .A(n_1019), .B(n_952), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_1017), .B(n_981), .Y(n_1040) );
NAND2xp33_ASAP7_75t_L g1041 ( .A(n_1038), .B(n_1015), .Y(n_1041) );
NAND2x1_ASAP7_75t_SL g1042 ( .A(n_1034), .B(n_1004), .Y(n_1042) );
AND2x4_ASAP7_75t_L g1043 ( .A(n_1022), .B(n_1012), .Y(n_1043) );
NOR3xp33_ASAP7_75t_L g1044 ( .A(n_1025), .B(n_996), .C(n_1020), .Y(n_1044) );
NOR2x1_ASAP7_75t_L g1045 ( .A(n_1034), .B(n_955), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_1027), .B(n_1009), .Y(n_1046) );
NOR3xp33_ASAP7_75t_L g1047 ( .A(n_1029), .B(n_999), .C(n_1000), .Y(n_1047) );
NOR3xp33_ASAP7_75t_L g1048 ( .A(n_1023), .B(n_1000), .C(n_1014), .Y(n_1048) );
O2A1O1Ixp33_ASAP7_75t_L g1049 ( .A1(n_1044), .A2(n_1036), .B(n_1037), .C(n_1028), .Y(n_1049) );
AOI32xp33_ASAP7_75t_L g1050 ( .A1(n_1041), .A2(n_993), .A3(n_1024), .B1(n_1022), .B2(n_1039), .Y(n_1050) );
NAND2xp5_ASAP7_75t_SL g1051 ( .A(n_1047), .B(n_1039), .Y(n_1051) );
OAI21xp33_ASAP7_75t_SL g1052 ( .A1(n_1042), .A2(n_1012), .B(n_1035), .Y(n_1052) );
NAND2x1p5_ASAP7_75t_L g1053 ( .A(n_1045), .B(n_1002), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_1048), .A2(n_1040), .B1(n_998), .B2(n_1012), .Y(n_1054) );
OAI21xp5_ASAP7_75t_L g1055 ( .A1(n_1041), .A2(n_1011), .B(n_1002), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_1048), .B(n_1033), .Y(n_1056) );
NOR2xp33_ASAP7_75t_L g1057 ( .A(n_1046), .B(n_1031), .Y(n_1057) );
NOR2x1_ASAP7_75t_L g1058 ( .A(n_1051), .B(n_1043), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_1057), .B(n_1056), .Y(n_1059) );
INVx2_ASAP7_75t_L g1060 ( .A(n_1053), .Y(n_1060) );
INVx2_ASAP7_75t_L g1061 ( .A(n_1053), .Y(n_1061) );
NAND2xp5_ASAP7_75t_SL g1062 ( .A(n_1052), .B(n_1050), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_1054), .A2(n_1032), .B1(n_1026), .B2(n_1030), .Y(n_1063) );
AOI21xp5_ASAP7_75t_L g1064 ( .A1(n_1062), .A2(n_1049), .B(n_1055), .Y(n_1064) );
AOI321xp33_ASAP7_75t_L g1065 ( .A1(n_1064), .A2(n_1058), .A3(n_1063), .B1(n_1059), .B2(n_1060), .C(n_1061), .Y(n_1065) );
OR3x1_ASAP7_75t_L g1066 ( .A(n_1065), .B(n_1013), .C(n_1008), .Y(n_1066) );
HB1xp67_ASAP7_75t_L g1067 ( .A(n_1066), .Y(n_1067) );
BUFx2_ASAP7_75t_L g1068 ( .A(n_1067), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1067), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1068), .Y(n_1070) );
OAI22xp5_ASAP7_75t_SL g1071 ( .A1(n_1069), .A2(n_975), .B1(n_976), .B2(n_973), .Y(n_1071) );
OAI22xp5_ASAP7_75t_SL g1072 ( .A1(n_1070), .A2(n_982), .B1(n_959), .B2(n_988), .Y(n_1072) );
NOR3xp33_ASAP7_75t_L g1073 ( .A(n_1072), .B(n_1071), .C(n_977), .Y(n_1073) );
INVxp67_ASAP7_75t_L g1074 ( .A(n_1073), .Y(n_1074) );
AOI21xp5_ASAP7_75t_L g1075 ( .A1(n_1074), .A2(n_997), .B(n_971), .Y(n_1075) );
endmodule