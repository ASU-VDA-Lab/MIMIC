module fake_aes_9123_n_15 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_15);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_9;
wire n_14;
wire n_7;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
NAND2xp5_ASAP7_75t_L g8 ( .A(n_2), .B(n_4), .Y(n_8) );
NAND2xp5_ASAP7_75t_SL g9 ( .A(n_1), .B(n_0), .Y(n_9) );
AOI22xp33_ASAP7_75t_L g10 ( .A1(n_7), .A2(n_3), .B1(n_5), .B2(n_9), .Y(n_10) );
INVx2_ASAP7_75t_SL g11 ( .A(n_8), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
XOR2xp5_ASAP7_75t_L g15 ( .A(n_14), .B(n_10), .Y(n_15) );
endmodule