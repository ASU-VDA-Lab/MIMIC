module fake_jpeg_9349_n_173 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_32),
.Y(n_46)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_36),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_0),
.Y(n_35)
);

OR2x2_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_37),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_23),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_27),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_32),
.A2(n_21),
.B1(n_16),
.B2(n_26),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_41),
.B1(n_29),
.B2(n_31),
.Y(n_68)
);

HAxp5_ASAP7_75t_SL g40 ( 
.A(n_38),
.B(n_26),
.CON(n_40),
.SN(n_40)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_33),
.B1(n_31),
.B2(n_19),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_21),
.B1(n_14),
.B2(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_51),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_21),
.B1(n_14),
.B2(n_16),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_50),
.B1(n_22),
.B2(n_30),
.Y(n_56)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_16),
.B1(n_22),
.B2(n_23),
.Y(n_50)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_53),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_58),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_57),
.B1(n_54),
.B2(n_47),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_33),
.B1(n_30),
.B2(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_35),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_37),
.B(n_30),
.C(n_28),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_19),
.B(n_15),
.C(n_25),
.Y(n_87)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_60),
.B(n_61),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_34),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_71),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_54),
.B1(n_47),
.B2(n_19),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_37),
.B(n_33),
.C(n_29),
.Y(n_69)
);

OAI32xp33_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_48),
.A3(n_34),
.B1(n_31),
.B2(n_52),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_37),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_SL g73 ( 
.A(n_72),
.B(n_45),
.C(n_53),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_82),
.B(n_78),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_39),
.B1(n_53),
.B2(n_48),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_72),
.B1(n_67),
.B2(n_61),
.Y(n_95)
);

XNOR2x2_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_69),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_78),
.B1(n_82),
.B2(n_62),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_54),
.B1(n_47),
.B2(n_18),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_65),
.B1(n_25),
.B2(n_15),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_13),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_80),
.B(n_87),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_18),
.B1(n_19),
.B2(n_25),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_88),
.Y(n_96)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_66),
.B(n_2),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_3),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_15),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_64),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_102),
.B1(n_109),
.B2(n_74),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_98),
.B(n_99),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_60),
.B(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_62),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_107),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_89),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_85),
.B(n_92),
.Y(n_122)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_105),
.B(n_108),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_15),
.Y(n_106)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_81),
.B(n_2),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_77),
.Y(n_110)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

XNOR2x1_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_87),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_103),
.B(n_96),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_84),
.C(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_124),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_84),
.C(n_81),
.Y(n_114)
);

AO21x1_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_122),
.B(n_97),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_115),
.B(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_93),
.A3(n_107),
.B1(n_102),
.B2(n_90),
.C1(n_80),
.C2(n_108),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_95),
.C(n_98),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_137),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_124),
.B(n_117),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_129),
.B(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_130),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_85),
.B1(n_65),
.B2(n_76),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_113),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_93),
.B1(n_97),
.B2(n_116),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_132),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_112),
.C(n_4),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_134),
.B(n_118),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_138),
.B(n_140),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_135),
.B(n_123),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_131),
.B(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_143),
.A2(n_126),
.B(n_136),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_128),
.B(n_127),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_125),
.B(n_4),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_34),
.C(n_15),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_34),
.C(n_4),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_148),
.A2(n_149),
.B(n_152),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_34),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_151),
.C(n_5),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_3),
.B(n_5),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_147),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_154),
.B(n_145),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_159),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_5),
.Y(n_159)
);

NAND4xp25_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_143),
.C(n_6),
.D(n_8),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_160),
.A2(n_156),
.B(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_6),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_165),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_161),
.A2(n_8),
.B(n_9),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_167),
.A2(n_10),
.B(n_11),
.Y(n_171)
);

BUFx4f_ASAP7_75t_SL g168 ( 
.A(n_164),
.Y(n_168)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_168),
.A2(n_163),
.B(n_10),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_171),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_169),
.Y(n_173)
);


endmodule