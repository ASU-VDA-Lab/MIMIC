module fake_jpeg_26354_n_155 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_155);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_18),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_66),
.Y(n_71)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_82),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_55),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_70),
.A2(n_41),
.B1(n_62),
.B2(n_49),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_75),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_41),
.B1(n_58),
.B2(n_52),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_45),
.B1(n_4),
.B2(n_5),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_59),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_59),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_45),
.B(n_48),
.C(n_51),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_43),
.B1(n_46),
.B2(n_54),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_60),
.B1(n_57),
.B2(n_53),
.Y(n_92)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_95),
.B1(n_6),
.B2(n_7),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_1),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_3),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_98),
.Y(n_108)
);

CKINVDCx11_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_99),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_109),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_112),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_86),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_13),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_108),
.B(n_94),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_83),
.B(n_95),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_115),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_7),
.B(n_8),
.C(n_10),
.Y(n_115)
);

CKINVDCx6p67_ASAP7_75t_R g116 ( 
.A(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_102),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_117),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_87),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_14),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_113),
.A2(n_106),
.B(n_107),
.Y(n_120)
);

AO21x1_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_122),
.B(n_132),
.Y(n_136)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_130),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_113),
.B(n_12),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_111),
.B(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_124),
.B(n_125),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_114),
.A2(n_109),
.B1(n_93),
.B2(n_85),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_16),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_20),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_21),
.C(n_22),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_133),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_SL g143 ( 
.A(n_135),
.B(n_128),
.C(n_133),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_142),
.C(n_131),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_129),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_144),
.C(n_145),
.Y(n_146)
);

XNOR2x1_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_126),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_140),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_136),
.Y(n_148)
);

NAND2xp33_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_141),
.B1(n_137),
.B2(n_134),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_24),
.C(n_28),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_38),
.B(n_30),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_29),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_31),
.Y(n_155)
);


endmodule