module fake_ibex_45_n_665 (n_85, n_84, n_64, n_3, n_73, n_65, n_55, n_63, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_70, n_7, n_20, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_13, n_61, n_14, n_0, n_12, n_42, n_77, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_83, n_32, n_53, n_50, n_11, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_54, n_19, n_665);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_55;
input n_63;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_70;
input n_7;
input n_20;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_13;
input n_61;
input n_14;
input n_0;
input n_12;
input n_42;
input n_77;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_83;
input n_32;
input n_53;
input n_50;
input n_11;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_54;
input n_19;

output n_665;

wire n_151;
wire n_599;
wire n_507;
wire n_540;
wire n_395;
wire n_171;
wire n_103;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_130;
wire n_177;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_124;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_108;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_452;
wire n_86;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_638;
wire n_398;
wire n_125;
wire n_304;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_94;
wire n_134;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_412;
wire n_88;
wire n_357;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_90;
wire n_449;
wire n_547;
wire n_176;
wire n_216;
wire n_652;
wire n_421;
wire n_475;
wire n_166;
wire n_163;
wire n_645;
wire n_500;
wire n_542;
wire n_114;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_556;
wire n_189;
wire n_498;
wire n_317;
wire n_280;
wire n_340;
wire n_375;
wire n_105;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_89;
wire n_144;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_113;
wire n_561;
wire n_117;
wire n_417;
wire n_471;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_91;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_228;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_426;
wire n_323;
wire n_469;
wire n_598;
wire n_143;
wire n_106;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_110;
wire n_306;
wire n_400;
wire n_550;
wire n_169;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_109;
wire n_127;
wire n_121;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_120;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_122;
wire n_523;
wire n_116;
wire n_614;
wire n_370;
wire n_431;
wire n_574;
wire n_289;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_136;
wire n_261;
wire n_521;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_654;
wire n_656;
wire n_437;
wire n_602;
wire n_355;
wire n_474;
wire n_594;
wire n_636;
wire n_407;
wire n_102;
wire n_490;
wire n_568;
wire n_448;
wire n_646;
wire n_595;
wire n_99;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_126;
wire n_623;
wire n_585;
wire n_530;
wire n_356;
wire n_104;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_141;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_331;
wire n_576;
wire n_230;
wire n_96;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_618;
wire n_514;
wire n_139;
wire n_488;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_129;
wire n_98;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_347;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_299;
wire n_87;
wire n_262;
wire n_433;
wire n_439;
wire n_643;
wire n_137;
wire n_338;
wire n_173;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_401;
wire n_554;
wire n_553;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_605;
wire n_539;
wire n_100;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_546;
wire n_199;
wire n_592;
wire n_495;
wire n_410;
wire n_308;
wire n_463;
wire n_624;
wire n_411;
wire n_135;
wire n_520;
wire n_658;
wire n_512;
wire n_615;
wire n_283;
wire n_366;
wire n_397;
wire n_111;
wire n_627;
wire n_322;
wire n_227;
wire n_499;
wire n_115;
wire n_248;
wire n_92;
wire n_451;
wire n_101;
wire n_190;
wire n_138;
wire n_650;
wire n_409;
wire n_582;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_332;
wire n_517;
wire n_211;
wire n_218;
wire n_314;
wire n_563;
wire n_132;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_633;
wire n_532;
wire n_95;
wire n_405;
wire n_415;
wire n_597;
wire n_320;
wire n_288;
wire n_247;
wire n_285;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_385;
wire n_233;
wire n_342;
wire n_414;
wire n_430;
wire n_118;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_639;
wire n_303;
wire n_362;
wire n_93;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_501;
wire n_266;
wire n_294;
wire n_112;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_119;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_97;
wire n_197;
wire n_528;
wire n_181;
wire n_131;
wire n_123;
wire n_631;
wire n_260;
wire n_620;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_107;
wire n_149;
wire n_489;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_159;
wire n_231;
wire n_202;
wire n_298;
wire n_587;
wire n_160;
wire n_657;
wire n_184;
wire n_492;
wire n_649;
wire n_232;
wire n_380;
wire n_281;
wire n_559;
wire n_425;

INVxp67_ASAP7_75t_SL g86 ( 
.A(n_15),
.Y(n_86)
);

INVxp67_ASAP7_75t_SL g87 ( 
.A(n_4),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_0),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_8),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_9),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVxp67_ASAP7_75t_SL g98 ( 
.A(n_16),
.Y(n_98)
);

INVxp33_ASAP7_75t_SL g99 ( 
.A(n_12),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_27),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_45),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_3),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_30),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVxp67_ASAP7_75t_SL g112 ( 
.A(n_47),
.Y(n_112)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_34),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_5),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_0),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g117 ( 
.A(n_23),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_21),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_25),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_36),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_50),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_17),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_2),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_24),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

INVxp67_ASAP7_75t_SL g131 ( 
.A(n_65),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_20),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_26),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_48),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_6),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_57),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_28),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_16),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_51),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_38),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_3),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_42),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_78),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_7),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g150 ( 
.A(n_52),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_5),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_18),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_4),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_12),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_44),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_82),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_31),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_2),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_1),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_159),
.Y(n_162)
);

AND2x4_ASAP7_75t_L g163 ( 
.A(n_102),
.B(n_1),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_88),
.B(n_7),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_114),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_103),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_88),
.B(n_8),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_122),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_96),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_94),
.B(n_39),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_117),
.B(n_9),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_90),
.B(n_10),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_110),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_95),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_89),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_110),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_129),
.B(n_10),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_92),
.B(n_11),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_95),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_97),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_11),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_124),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_97),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_104),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_124),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_143),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_13),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_152),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_105),
.B(n_13),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_120),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_133),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_99),
.A2(n_154),
.B1(n_153),
.B2(n_87),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_133),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_138),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_138),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_145),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_140),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_100),
.B(n_14),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_86),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_93),
.B(n_14),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_106),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_107),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_108),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_145),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_109),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_156),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_111),
.B(n_15),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_118),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_98),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_119),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_121),
.B(n_17),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_127),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_130),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_132),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_156),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_163),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_165),
.Y(n_239)
);

AO22x2_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_158),
.B1(n_135),
.B2(n_137),
.Y(n_240)
);

OAI221xp5_ASAP7_75t_L g241 ( 
.A1(n_175),
.A2(n_134),
.B1(n_150),
.B2(n_113),
.C(n_131),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_147),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_163),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_163),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_142),
.Y(n_246)
);

AND2x4_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_141),
.Y(n_247)
);

AND2x6_ASAP7_75t_L g248 ( 
.A(n_177),
.B(n_157),
.Y(n_248)
);

AND2x6_ASAP7_75t_L g249 ( 
.A(n_177),
.B(n_112),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_205),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_123),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_197),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_168),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_123),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_165),
.B(n_100),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_169),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_182),
.A2(n_99),
.B1(n_101),
.B2(n_18),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_178),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_213),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_167),
.B(n_19),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_174),
.Y(n_265)
);

AND2x4_ASAP7_75t_L g266 ( 
.A(n_182),
.B(n_19),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_168),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_196),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_199),
.B(n_33),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_196),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_181),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_169),
.Y(n_272)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_206),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_200),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_167),
.B(n_37),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_178),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_200),
.Y(n_277)
);

NAND2x1p5_ASAP7_75t_L g278 ( 
.A(n_219),
.B(n_43),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_193),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_171),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_215),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_171),
.Y(n_282)
);

AND2x4_ASAP7_75t_L g283 ( 
.A(n_199),
.B(n_46),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_201),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_208),
.B(n_49),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_183),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_172),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_172),
.B(n_54),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_208),
.B(n_55),
.Y(n_289)
);

AND2x4_ASAP7_75t_L g290 ( 
.A(n_193),
.B(n_58),
.Y(n_290)
);

OA22x2_ASAP7_75t_L g291 ( 
.A1(n_234),
.A2(n_236),
.B1(n_218),
.B2(n_222),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_201),
.Y(n_292)
);

AND2x6_ASAP7_75t_L g293 ( 
.A(n_219),
.B(n_61),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_178),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_234),
.B(n_68),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_173),
.B(n_85),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_183),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_203),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_176),
.A2(n_72),
.B1(n_76),
.B2(n_185),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_186),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_186),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_236),
.B(n_211),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_160),
.Y(n_303)
);

AO21x2_ASAP7_75t_L g304 ( 
.A1(n_221),
.A2(n_233),
.B(n_229),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_174),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_187),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_206),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_187),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_184),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_206),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_188),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_173),
.B(n_190),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_206),
.B(n_217),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_230),
.B(n_235),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_224),
.B(n_232),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_228),
.A2(n_198),
.B1(n_226),
.B2(n_216),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_176),
.A2(n_191),
.B1(n_192),
.B2(n_166),
.Y(n_317)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_206),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_225),
.B(n_227),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_162),
.B(n_202),
.Y(n_320)
);

NAND2x1p5_ASAP7_75t_L g321 ( 
.A(n_207),
.B(n_230),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_235),
.B(n_161),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_178),
.Y(n_323)
);

AO22x2_ASAP7_75t_L g324 ( 
.A1(n_170),
.A2(n_204),
.B1(n_164),
.B2(n_202),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_178),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_180),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_179),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_194),
.B(n_180),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_189),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_189),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_198),
.B(n_237),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_279),
.B(n_209),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_209),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_239),
.B(n_214),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_214),
.B1(n_216),
.B2(n_226),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_239),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_317),
.A2(n_237),
.B1(n_249),
.B2(n_303),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_266),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_304),
.B(n_257),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_R g341 ( 
.A(n_262),
.B(n_281),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_283),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_278),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_283),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_250),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_322),
.Y(n_346)
);

NOR3xp33_ASAP7_75t_SL g347 ( 
.A(n_299),
.B(n_331),
.C(n_241),
.Y(n_347)
);

BUFx2_ASAP7_75t_SL g348 ( 
.A(n_293),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_272),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_326),
.Y(n_350)
);

NOR2xp67_ASAP7_75t_L g351 ( 
.A(n_299),
.B(n_241),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_314),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_259),
.A2(n_254),
.B1(n_252),
.B2(n_279),
.Y(n_353)
);

OR2x2_ASAP7_75t_SL g354 ( 
.A(n_331),
.B(n_271),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_322),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_312),
.Y(n_356)
);

BUFx4_ASAP7_75t_SL g357 ( 
.A(n_298),
.Y(n_357)
);

AND2x4_ASAP7_75t_L g358 ( 
.A(n_246),
.B(n_247),
.Y(n_358)
);

INVx5_ASAP7_75t_L g359 ( 
.A(n_293),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_304),
.B(n_257),
.Y(n_360)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_293),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_244),
.A2(n_245),
.B(n_302),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_R g363 ( 
.A(n_258),
.B(n_287),
.Y(n_363)
);

AO22x1_ASAP7_75t_L g364 ( 
.A1(n_293),
.A2(n_249),
.B1(n_248),
.B2(n_320),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_253),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_246),
.B(n_247),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_302),
.B(n_256),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_291),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_263),
.B(n_290),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_328),
.B(n_265),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_243),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_249),
.A2(n_291),
.B1(n_293),
.B2(n_248),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_253),
.B(n_256),
.Y(n_373)
);

OR2x6_ASAP7_75t_L g374 ( 
.A(n_316),
.B(n_329),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_305),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_290),
.B(n_315),
.Y(n_376)
);

BUFx12f_ASAP7_75t_L g377 ( 
.A(n_248),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_248),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_R g379 ( 
.A(n_330),
.B(n_238),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_251),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_314),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_278),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_248),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_238),
.B(n_311),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_300),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_288),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_309),
.B(n_315),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_249),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_321),
.B(n_275),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_328),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_301),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_321),
.Y(n_392)
);

AO22x1_ASAP7_75t_L g393 ( 
.A1(n_249),
.A2(n_296),
.B1(n_319),
.B2(n_242),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_261),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_306),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_308),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_319),
.B(n_240),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_260),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_318),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_264),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_268),
.B(n_284),
.Y(n_401)
);

INVx5_ASAP7_75t_L g402 ( 
.A(n_307),
.Y(n_402)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_307),
.Y(n_403)
);

NAND3xp33_ASAP7_75t_SL g404 ( 
.A(n_259),
.B(n_295),
.C(n_285),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_R g405 ( 
.A(n_242),
.B(n_274),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_255),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_318),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_270),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_295),
.B(n_292),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_269),
.B(n_289),
.Y(n_410)
);

NOR3xp33_ASAP7_75t_SL g411 ( 
.A(n_269),
.B(n_289),
.C(n_285),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_267),
.B(n_286),
.Y(n_412)
);

A2O1A1Ixp33_ASAP7_75t_L g413 ( 
.A1(n_340),
.A2(n_360),
.B(n_362),
.C(n_373),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_358),
.B(n_324),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_343),
.B(n_280),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_382),
.B(n_297),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_385),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_358),
.B(n_282),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_361),
.Y(n_419)
);

INVx5_ASAP7_75t_L g420 ( 
.A(n_361),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_346),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_351),
.A2(n_324),
.B1(n_240),
.B2(n_277),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_355),
.A2(n_324),
.B1(n_240),
.B2(n_313),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_363),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_349),
.B(n_313),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_350),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_387),
.Y(n_427)
);

AND2x2_ASAP7_75t_SL g428 ( 
.A(n_372),
.B(n_310),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_376),
.B(n_273),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_366),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_412),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_390),
.A2(n_273),
.B1(n_323),
.B2(n_325),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_367),
.B(n_273),
.Y(n_433)
);

NAND2xp33_ASAP7_75t_L g434 ( 
.A(n_342),
.B(n_261),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_368),
.A2(n_273),
.B1(n_261),
.B2(n_276),
.Y(n_435)
);

INVx3_ASAP7_75t_SL g436 ( 
.A(n_375),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_369),
.B(n_276),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_340),
.A2(n_360),
.B(n_373),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_369),
.B(n_276),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_412),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_367),
.A2(n_294),
.B(n_410),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_376),
.B(n_294),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_348),
.B(n_294),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_387),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_406),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g446 ( 
.A(n_332),
.B(n_294),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_341),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_352),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_364),
.B(n_377),
.Y(n_449)
);

AND2x2_ASAP7_75t_SL g450 ( 
.A(n_335),
.B(n_388),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_336),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_338),
.B(n_339),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_342),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_342),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_356),
.B(n_370),
.Y(n_455)
);

AOI222xp33_ASAP7_75t_L g456 ( 
.A1(n_353),
.A2(n_397),
.B1(n_334),
.B2(n_333),
.C1(n_365),
.C2(n_352),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_334),
.B(n_365),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_338),
.B(n_339),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_359),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_357),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_354),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_357),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_392),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_344),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_381),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_386),
.B(n_347),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_379),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_388),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_344),
.A2(n_347),
.B1(n_353),
.B2(n_337),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_405),
.Y(n_470)
);

CKINVDCx8_ASAP7_75t_R g471 ( 
.A(n_374),
.Y(n_471)
);

O2A1O1Ixp33_ASAP7_75t_L g472 ( 
.A1(n_404),
.A2(n_362),
.B(n_401),
.C(n_408),
.Y(n_472)
);

NOR3xp33_ASAP7_75t_L g473 ( 
.A(n_393),
.B(n_404),
.C(n_389),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_374),
.B(n_381),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_401),
.A2(n_409),
.B1(n_359),
.B2(n_400),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_406),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_399),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_391),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_359),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_374),
.B(n_383),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_384),
.A2(n_345),
.B(n_396),
.Y(n_481)
);

CKINVDCx8_ASAP7_75t_R g482 ( 
.A(n_378),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_395),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_398),
.B(n_371),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_380),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_427),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_444),
.Y(n_487)
);

AOI221xp5_ASAP7_75t_L g488 ( 
.A1(n_455),
.A2(n_411),
.B1(n_407),
.B2(n_403),
.C(n_402),
.Y(n_488)
);

AO21x2_ASAP7_75t_L g489 ( 
.A1(n_473),
.A2(n_411),
.B(n_394),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_421),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_457),
.B(n_402),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_438),
.B(n_402),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_419),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_451),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_426),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_478),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_468),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_433),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_433),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_483),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_484),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_485),
.Y(n_502)
);

AND2x2_ASAP7_75t_SL g503 ( 
.A(n_422),
.B(n_403),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_456),
.B(n_413),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_424),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_472),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_470),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_466),
.A2(n_414),
.B1(n_460),
.B2(n_461),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_479),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_472),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_420),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_420),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_442),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_468),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_446),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_479),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_456),
.A2(n_450),
.B1(n_430),
.B2(n_469),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_480),
.B(n_474),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_442),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_436),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_419),
.Y(n_521)
);

NAND3xp33_ASAP7_75t_SL g522 ( 
.A(n_422),
.B(n_471),
.C(n_462),
.Y(n_522)
);

OA21x2_ASAP7_75t_L g523 ( 
.A1(n_441),
.A2(n_473),
.B(n_475),
.Y(n_523)
);

OR2x6_ASAP7_75t_L g524 ( 
.A(n_449),
.B(n_480),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_423),
.B(n_440),
.Y(n_525)
);

AO21x2_ASAP7_75t_L g526 ( 
.A1(n_423),
.A2(n_481),
.B(n_429),
.Y(n_526)
);

NAND2x1p5_ASAP7_75t_L g527 ( 
.A(n_420),
.B(n_419),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_449),
.A2(n_440),
.B1(n_431),
.B2(n_417),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_436),
.A2(n_447),
.B1(n_467),
.B2(n_452),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_452),
.A2(n_458),
.B1(n_418),
.B2(n_416),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_418),
.B(n_415),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_458),
.A2(n_448),
.B1(n_465),
.B2(n_425),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_448),
.A2(n_465),
.B1(n_416),
.B2(n_415),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_453),
.Y(n_534)
);

AO21x2_ASAP7_75t_L g535 ( 
.A1(n_481),
.A2(n_432),
.B(n_434),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_477),
.A2(n_428),
.B1(n_449),
.B2(n_437),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_420),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_477),
.A2(n_437),
.B1(n_439),
.B2(n_463),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_453),
.A2(n_454),
.B1(n_464),
.B2(n_482),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_439),
.B(n_476),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_453),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_454),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_459),
.B(n_445),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_464),
.A2(n_459),
.B1(n_479),
.B2(n_435),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_435),
.A2(n_444),
.B1(n_427),
.B2(n_438),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_443),
.Y(n_547)
);

AND2x4_ASAP7_75t_SL g548 ( 
.A(n_443),
.B(n_427),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_522),
.A2(n_517),
.B1(n_504),
.B2(n_487),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_486),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_486),
.B(n_487),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_512),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_R g553 ( 
.A(n_547),
.B(n_504),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_498),
.A2(n_499),
.B1(n_503),
.B2(n_501),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_501),
.B(n_490),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_490),
.B(n_494),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_503),
.A2(n_499),
.B1(n_498),
.B2(n_524),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_524),
.A2(n_508),
.B1(n_514),
.B2(n_497),
.Y(n_558)
);

OAI221xp5_ASAP7_75t_L g559 ( 
.A1(n_532),
.A2(n_507),
.B1(n_530),
.B2(n_529),
.C(n_533),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_546),
.A2(n_514),
.B1(n_497),
.B2(n_525),
.Y(n_560)
);

OAI221xp5_ASAP7_75t_L g561 ( 
.A1(n_536),
.A2(n_520),
.B1(n_495),
.B2(n_538),
.C(n_502),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_512),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_502),
.Y(n_563)
);

OAI211xp5_ASAP7_75t_L g564 ( 
.A1(n_488),
.A2(n_515),
.B(n_505),
.C(n_540),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_524),
.A2(n_518),
.B1(n_531),
.B2(n_528),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_524),
.A2(n_518),
.B1(n_531),
.B2(n_519),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_534),
.Y(n_567)
);

AOI222xp33_ASAP7_75t_L g568 ( 
.A1(n_494),
.A2(n_518),
.B1(n_519),
.B2(n_513),
.C1(n_506),
.C2(n_510),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_496),
.A2(n_500),
.B1(n_513),
.B2(n_491),
.Y(n_569)
);

BUFx4f_ASAP7_75t_SL g570 ( 
.A(n_512),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_496),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_548),
.A2(n_547),
.B1(n_492),
.B2(n_511),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_492),
.Y(n_573)
);

AOI221xp5_ASAP7_75t_L g574 ( 
.A1(n_526),
.A2(n_539),
.B1(n_543),
.B2(n_489),
.C(n_545),
.Y(n_574)
);

AOI221xp5_ASAP7_75t_L g575 ( 
.A1(n_526),
.A2(n_543),
.B1(n_489),
.B2(n_511),
.C(n_537),
.Y(n_575)
);

OAI221xp5_ASAP7_75t_L g576 ( 
.A1(n_523),
.A2(n_537),
.B1(n_527),
.B2(n_521),
.C(n_493),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_527),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_489),
.A2(n_543),
.B1(n_526),
.B2(n_537),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_523),
.A2(n_535),
.B1(n_493),
.B2(n_521),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_523),
.A2(n_535),
.B1(n_493),
.B2(n_521),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_534),
.Y(n_581)
);

AOI31xp33_ASAP7_75t_L g582 ( 
.A1(n_527),
.A2(n_541),
.A3(n_516),
.B(n_509),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_542),
.A2(n_522),
.B1(n_455),
.B2(n_466),
.Y(n_583)
);

AOI222xp33_ASAP7_75t_L g584 ( 
.A1(n_548),
.A2(n_351),
.B1(n_455),
.B2(n_353),
.C1(n_316),
.C2(n_466),
.Y(n_584)
);

OAI31xp33_ASAP7_75t_L g585 ( 
.A1(n_564),
.A2(n_542),
.A3(n_544),
.B(n_554),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_573),
.B(n_542),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_573),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_571),
.B(n_544),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_559),
.B(n_561),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_571),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_584),
.A2(n_549),
.B1(n_568),
.B2(n_560),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_550),
.Y(n_592)
);

BUFx2_ASAP7_75t_SL g593 ( 
.A(n_562),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_551),
.B(n_550),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_557),
.A2(n_583),
.B1(n_551),
.B2(n_558),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_563),
.B(n_556),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_578),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_555),
.B(n_569),
.Y(n_598)
);

AOI33xp33_ASAP7_75t_L g599 ( 
.A1(n_566),
.A2(n_565),
.A3(n_580),
.B1(n_579),
.B2(n_575),
.B3(n_574),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_576),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_562),
.B(n_552),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_562),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_572),
.B(n_581),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_552),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_581),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_L g606 ( 
.A1(n_582),
.A2(n_577),
.B(n_553),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_594),
.B(n_567),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_592),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_592),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_594),
.B(n_567),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_602),
.Y(n_611)
);

AOI221xp5_ASAP7_75t_L g612 ( 
.A1(n_591),
.A2(n_553),
.B1(n_567),
.B2(n_570),
.C(n_589),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_591),
.A2(n_567),
.B1(n_589),
.B2(n_595),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_590),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_594),
.B(n_567),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_595),
.A2(n_606),
.B1(n_598),
.B2(n_593),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_606),
.A2(n_598),
.B1(n_593),
.B2(n_600),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_592),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_607),
.B(n_596),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_607),
.B(n_596),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_611),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_610),
.B(n_596),
.Y(n_622)
);

NOR4xp25_ASAP7_75t_SL g623 ( 
.A(n_612),
.B(n_605),
.C(n_602),
.D(n_585),
.Y(n_623)
);

INVxp67_ASAP7_75t_SL g624 ( 
.A(n_614),
.Y(n_624)
);

NAND4xp25_ASAP7_75t_L g625 ( 
.A(n_616),
.B(n_599),
.C(n_585),
.D(n_600),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_614),
.A2(n_601),
.B(n_602),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_619),
.B(n_618),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_624),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_620),
.Y(n_629)
);

OAI211xp5_ASAP7_75t_L g630 ( 
.A1(n_625),
.A2(n_612),
.B(n_613),
.C(n_617),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_622),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_626),
.B(n_621),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_623),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_623),
.A2(n_611),
.B1(n_602),
.B2(n_604),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_627),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_628),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_629),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_631),
.B(n_615),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_628),
.B(n_615),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_632),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_638),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_635),
.B(n_632),
.Y(n_642)
);

AOI221xp5_ASAP7_75t_L g643 ( 
.A1(n_640),
.A2(n_630),
.B1(n_633),
.B2(n_634),
.C(n_600),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_R g644 ( 
.A(n_637),
.B(n_611),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_636),
.B(n_618),
.Y(n_645)
);

AOI322xp5_ASAP7_75t_L g646 ( 
.A1(n_640),
.A2(n_610),
.A3(n_600),
.B1(n_597),
.B2(n_601),
.C1(n_609),
.C2(n_608),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_645),
.Y(n_647)
);

INVxp33_ASAP7_75t_L g648 ( 
.A(n_644),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_641),
.Y(n_649)
);

AOI311xp33_ASAP7_75t_L g650 ( 
.A1(n_643),
.A2(n_609),
.A3(n_608),
.B(n_605),
.C(n_603),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_642),
.A2(n_639),
.B1(n_636),
.B2(n_601),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_649),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_647),
.Y(n_653)
);

NOR3xp33_ASAP7_75t_L g654 ( 
.A(n_651),
.B(n_650),
.C(n_648),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_653),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_652),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_656),
.B(n_648),
.Y(n_657)
);

OAI222xp33_ASAP7_75t_L g658 ( 
.A1(n_655),
.A2(n_654),
.B1(n_639),
.B2(n_646),
.C1(n_601),
.C2(n_603),
.Y(n_658)
);

NOR3xp33_ASAP7_75t_L g659 ( 
.A(n_655),
.B(n_599),
.C(n_601),
.Y(n_659)
);

AND2x4_ASAP7_75t_SL g660 ( 
.A(n_657),
.B(n_588),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_659),
.Y(n_661)
);

OAI222xp33_ASAP7_75t_L g662 ( 
.A1(n_661),
.A2(n_658),
.B1(n_586),
.B2(n_604),
.C1(n_597),
.C2(n_587),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_660),
.Y(n_663)
);

AOI222xp33_ASAP7_75t_L g664 ( 
.A1(n_663),
.A2(n_604),
.B1(n_588),
.B2(n_597),
.C1(n_590),
.C2(n_587),
.Y(n_664)
);

AOI221xp5_ASAP7_75t_L g665 ( 
.A1(n_664),
.A2(n_663),
.B1(n_662),
.B2(n_604),
.C(n_588),
.Y(n_665)
);


endmodule