module real_jpeg_7550_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_1),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_2),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_2),
.A2(n_44),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_2),
.A2(n_44),
.B1(n_72),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_2),
.A2(n_44),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_2),
.B(n_127),
.C(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_2),
.B(n_242),
.Y(n_241)
);

O2A1O1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_2),
.A2(n_249),
.B(n_251),
.C(n_252),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_2),
.B(n_262),
.C(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_2),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_2),
.B(n_136),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_2),
.B(n_23),
.Y(n_288)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_4),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_4),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_4),
.Y(n_275)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_5),
.Y(n_231)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_7),
.A2(n_79),
.B1(n_83),
.B2(n_86),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_7),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_7),
.A2(n_86),
.B1(n_104),
.B2(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_7),
.A2(n_86),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_8),
.Y(n_227)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_9),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_10),
.A2(n_71),
.B1(n_74),
.B2(n_76),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_10),
.A2(n_76),
.B1(n_112),
.B2(n_116),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_10),
.A2(n_76),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_11),
.Y(n_338)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_333),
.B(n_336),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_168),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_167),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_18),
.B(n_128),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_122),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_22),
.B2(n_121),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_46),
.B1(n_47),
.B2(n_121),
.Y(n_21)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_22),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_22),
.A2(n_121),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_22),
.A2(n_143),
.B(n_166),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_L g176 ( 
.A(n_22),
.B(n_137),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_22),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_22),
.B(n_204),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_22),
.A2(n_121),
.B1(n_145),
.B2(n_166),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_22),
.A2(n_121),
.B1(n_245),
.B2(n_255),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_22),
.B(n_186),
.Y(n_318)
);

OA21x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_33),
.B(n_42),
.Y(n_22)
);

NOR2x1_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_34),
.Y(n_33)
);

AO22x1_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_29),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_29),
.Y(n_126)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_34)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_44),
.A2(n_101),
.B(n_104),
.Y(n_251)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_77),
.B1(n_119),
.B2(n_120),
.Y(n_47)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_48),
.B(n_121),
.C(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_48),
.A2(n_119),
.B1(n_123),
.B2(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_59),
.B(n_70),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_49),
.A2(n_59),
.B1(n_161),
.B2(n_165),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_49),
.B(n_59),
.Y(n_187)
);

NAND2x1_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_59),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_58),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_53),
.Y(n_263)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_56),
.Y(n_164)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_65),
.B2(n_69),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_60),
.B(n_272),
.Y(n_271)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_62),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_62),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_68),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g264 ( 
.A(n_73),
.Y(n_264)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_87),
.B1(n_100),
.B2(n_111),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_78),
.A2(n_87),
.B1(n_100),
.B2(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AO21x2_ASAP7_75t_SL g137 ( 
.A1(n_88),
.A2(n_100),
.B(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_100),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_89)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_90),
.Y(n_250)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_100),
.Y(n_242)
);

OA22x2_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_103),
.B1(n_105),
.B2(n_108),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_118),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_121),
.A2(n_137),
.B(n_206),
.C(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_128),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_128),
.B(n_331),
.Y(n_332)
);

FAx1_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_138),
.CI(n_142),
.CON(n_128),
.SN(n_128)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_129),
.A2(n_204),
.B(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_137),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_130),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_130)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_137),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_137),
.A2(n_186),
.B1(n_204),
.B2(n_221),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_137),
.A2(n_204),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_143),
.A2(n_144),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_160),
.Y(n_144)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_160),
.B1(n_166),
.B2(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_154),
.Y(n_145)
);

INVxp33_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_147),
.B(n_196),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_154),
.B1(n_179),
.B2(n_182),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_179),
.B1(n_195),
.B2(n_201),
.Y(n_194)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_152),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AND2x4_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_187),
.Y(n_186)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_330),
.B(n_332),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI211xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_235),
.B(n_324),
.C(n_329),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_217),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g324 ( 
.A1(n_173),
.A2(n_217),
.B(n_325),
.C(n_328),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_207),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_174),
.B(n_207),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_190),
.C(n_192),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_175),
.B(n_190),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_188),
.B2(n_189),
.Y(n_175)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_176),
.B(n_193),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_176),
.A2(n_188),
.B1(n_224),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_177),
.A2(n_203),
.B(n_205),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_186),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_178),
.A2(n_186),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_186),
.B(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_186),
.A2(n_221),
.B1(n_241),
.B2(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_186),
.A2(n_221),
.B1(n_259),
.B2(n_260),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_186),
.A2(n_221),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

O2A1O1Ixp33_ASAP7_75t_L g292 ( 
.A1(n_186),
.A2(n_204),
.B(n_247),
.C(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_186),
.B(n_204),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_186),
.A2(n_194),
.B1(n_221),
.B2(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_203),
.B(n_205),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_194),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_204),
.B(n_232),
.C(n_287),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AND3x1_ASAP7_75t_L g317 ( 
.A(n_206),
.B(n_294),
.C(n_318),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_216),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_211),
.B(n_213),
.C(n_216),
.Y(n_331)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_233),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_218),
.B(n_233),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.C(n_223),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_219),
.B(n_220),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_241),
.C(n_243),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_221),
.B(n_284),
.C(n_291),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_223),
.B(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_224),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_232),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_225),
.A2(n_226),
.B1(n_232),
.B2(n_243),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_232),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_232),
.A2(n_243),
.B1(n_248),
.B2(n_254),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_232),
.B(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_232),
.A2(n_243),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_232),
.B(n_248),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_306),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_296),
.B(n_305),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_282),
.B(n_295),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_256),
.B(n_281),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_240),
.B(n_244),
.Y(n_281)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_243),
.B(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_243),
.B(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_255),
.Y(n_244)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_268),
.B(n_280),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_265),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_265),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_278),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_276),
.Y(n_269)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_292),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_292),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_289),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_298),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_302),
.C(n_303),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NOR2x1_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_319),
.Y(n_306)
);

NOR2x1_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_309),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_316),
.B2(n_317),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_316),
.C(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_319),
.A2(n_326),
.B(n_327),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_322),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx12f_ASAP7_75t_L g337 ( 
.A(n_334),
.Y(n_337)
);

INVx13_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);


endmodule