module real_jpeg_14652_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_286, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_286;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_249;
wire n_78;
wire n_83;
wire n_176;
wire n_215;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_271;
wire n_47;
wire n_131;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_205;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_244;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_181;
wire n_85;
wire n_102;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_3),
.A2(n_15),
.B(n_282),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_3),
.B(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_6),
.A2(n_23),
.B1(n_26),
.B2(n_36),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_6),
.A2(n_8),
.B(n_32),
.C(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_6),
.A2(n_36),
.B1(n_56),
.B2(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_6),
.B(n_37),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_6),
.B(n_54),
.C(n_57),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_6),
.B(n_44),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_6),
.B(n_29),
.C(n_33),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

AO22x1_ASAP7_75t_L g44 ( 
.A1(n_8),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g283 ( 
.A(n_9),
.Y(n_283)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_11),
.A2(n_23),
.B1(n_26),
.B2(n_48),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_11),
.A2(n_48),
.B1(n_56),
.B2(n_57),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_12),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_12),
.A2(n_25),
.B1(n_45),
.B2(n_46),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_12),
.A2(n_25),
.B1(n_56),
.B2(n_57),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_13),
.A2(n_23),
.B1(n_26),
.B2(n_40),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_13),
.A2(n_40),
.B1(n_56),
.B2(n_57),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_13),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_74),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_72),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_69),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_18),
.B(n_69),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_62),
.C(n_66),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_19),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_38),
.C(n_49),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_20),
.A2(n_108),
.B1(n_118),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_20),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_20),
.B(n_118),
.C(n_181),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_20),
.A2(n_84),
.B1(n_85),
.B2(n_183),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_20),
.A2(n_183),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B1(n_35),
.B2(n_37),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g171 ( 
.A1(n_22),
.A2(n_31),
.B(n_68),
.Y(n_171)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_26),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_27),
.B(n_35),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_27),
.B(n_37),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_31),
.A2(n_67),
.B(n_68),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_31),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_42),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g239 ( 
.A(n_35),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_SL g97 ( 
.A1(n_36),
.A2(n_42),
.B(n_45),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_36),
.B(n_104),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_36),
.B(n_60),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_38),
.A2(n_49),
.B1(n_257),
.B2(n_271),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_38),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_44),
.B2(n_47),
.Y(n_38)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_39),
.Y(n_259)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_41),
.B(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_46),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_49),
.A2(n_257),
.B1(n_258),
.B2(n_260),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_49),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_49),
.B(n_171),
.C(n_258),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_60),
.B(n_61),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_50),
.A2(n_60),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_93),
.Y(n_92)
);

AO22x1_ASAP7_75t_SL g123 ( 
.A1(n_51),
.A2(n_55),
.B1(n_91),
.B2(n_93),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_51),
.A2(n_55),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

AO22x1_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_56),
.B(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OA21x2_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_90),
.B(n_92),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_60),
.A2(n_92),
.B(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_61),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_62),
.B(n_66),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_64),
.A2(n_65),
.B1(n_86),
.B2(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_64),
.A2(n_65),
.B(n_109),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_65),
.A2(n_87),
.B(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_277),
.B(n_281),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_249),
.B(n_274),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_227),
.B(n_248),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_210),
.B(n_226),
.Y(n_78)
);

OAI321xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_178),
.A3(n_205),
.B1(n_208),
.B2(n_209),
.C(n_286),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_160),
.B(n_177),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_126),
.B(n_159),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_105),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_83),
.B(n_105),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.C(n_94),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_84),
.A2(n_85),
.B1(n_89),
.B2(n_143),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_84),
.A2(n_85),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_85),
.B(n_170),
.C(n_175),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_85),
.B(n_183),
.C(n_215),
.Y(n_247)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_89),
.B(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_89),
.A2(n_130),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_89),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_89),
.A2(n_143),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_94),
.A2(n_95),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_98),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_100),
.B(n_203),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_103),
.A2(n_104),
.B1(n_186),
.B2(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_104),
.A2(n_116),
.B(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_120),
.B2(n_121),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_106),
.B(n_123),
.C(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_110),
.B1(n_118),
.B2(n_119),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_108),
.B(n_111),
.C(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_113),
.B(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_114),
.B(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_118),
.A2(n_243),
.B(n_246),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_118),
.B(n_243),
.Y(n_246)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_122),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_123),
.A2(n_125),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_135),
.C(n_137),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_123),
.A2(n_125),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_123),
.B(n_202),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_153),
.B(n_158),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_139),
.B(n_152),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_132),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_130),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_132)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_134),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_137),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_137),
.B(n_149),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_166),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_144),
.B(n_151),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_185),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_148),
.B(n_150),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_154),
.B(n_155),
.Y(n_158)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_162),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_169),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_165),
.C(n_169),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_170),
.A2(n_171),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_170),
.B(n_193),
.C(n_198),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_170),
.A2(n_171),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_170),
.A2(n_171),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_171),
.B(n_268),
.C(n_272),
.Y(n_280)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_189),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_189),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.C(n_188),
.Y(n_179)
);

FAx1_ASAP7_75t_SL g207 ( 
.A(n_180),
.B(n_184),
.CI(n_188),
.CON(n_207),
.SN(n_207)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_185),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_204),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_199),
.B2(n_200),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_200),
.C(n_204),
.Y(n_225)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_206),
.B(n_207),
.Y(n_208)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_207),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_225),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_225),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_214),
.C(n_219),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_219),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_224),
.Y(n_219)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_220),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_222),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_220),
.A2(n_224),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_224),
.A2(n_233),
.B(n_238),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_229),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_247),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_241),
.B2(n_242),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_241),
.C(n_247),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_246),
.A2(n_253),
.B1(n_254),
.B2(n_261),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_246),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_264),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_263),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_263),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_262),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_261),
.C(n_262),
.Y(n_273)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_258),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_273),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_273),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_272),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_280),
.Y(n_281)
);


endmodule