module fake_jpeg_22924_n_303 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_265;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_41),
.Y(n_49)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_20),
.B1(n_33),
.B2(n_19),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_55),
.B(n_62),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_24),
.B1(n_33),
.B2(n_31),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_53),
.A2(n_54),
.B1(n_62),
.B2(n_26),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_18),
.B1(n_21),
.B2(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_28),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_59),
.Y(n_88)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_24),
.B1(n_27),
.B2(n_30),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_44),
.B1(n_28),
.B2(n_36),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_69),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_19),
.B1(n_30),
.B2(n_22),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_65),
.A2(n_67),
.B1(n_70),
.B2(n_73),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_36),
.B1(n_31),
.B2(n_25),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_68),
.A2(n_74),
.B1(n_42),
.B2(n_37),
.Y(n_122)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_17),
.B1(n_23),
.B2(n_29),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_77),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_17),
.B1(n_35),
.B2(n_32),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_31),
.B1(n_35),
.B2(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_83),
.B1(n_98),
.B2(n_25),
.Y(n_103)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_80),
.Y(n_116)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_35),
.B(n_32),
.C(n_26),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_81),
.B(n_94),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_84),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_54),
.A2(n_35),
.B1(n_32),
.B2(n_26),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_53),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_86),
.B(n_87),
.Y(n_113)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_89),
.B(n_95),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_46),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_0),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_96),
.B(n_99),
.Y(n_114)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_62),
.A2(n_26),
.B1(n_25),
.B2(n_31),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_55),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_9),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_0),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_8),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_103),
.A2(n_105),
.B1(n_92),
.B2(n_91),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_25),
.B1(n_42),
.B2(n_37),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_78),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_100),
.A2(n_42),
.B1(n_37),
.B2(n_3),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_130),
.B1(n_72),
.B2(n_94),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_87),
.C(n_68),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_123),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_99),
.B(n_63),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_121),
.A2(n_126),
.B(n_128),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_122),
.A2(n_81),
.B1(n_97),
.B2(n_64),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_8),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_88),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_1),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_1),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_2),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_88),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_79),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_132),
.B(n_136),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_134),
.A2(n_140),
.B1(n_148),
.B2(n_156),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_153),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_72),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_144),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_138),
.B(n_149),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_89),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_141),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_77),
.B1(n_69),
.B2(n_93),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_96),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_146),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_90),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_112),
.B(n_110),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_95),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_75),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_150),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_75),
.B1(n_91),
.B2(n_80),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_75),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_131),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_151),
.Y(n_169)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_117),
.B(n_2),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_155),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_112),
.B(n_3),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_157),
.B(n_160),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_85),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_143),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_111),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_108),
.Y(n_172)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_133),
.B(n_123),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_143),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_111),
.B(n_128),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_162),
.A2(n_118),
.B(n_102),
.Y(n_209)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_167),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_122),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_176),
.C(n_126),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_166),
.Y(n_213)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_187),
.B(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_173),
.B(n_175),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_110),
.C(n_119),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_178),
.B(n_182),
.Y(n_206)
);

INVx3_ASAP7_75t_SL g181 ( 
.A(n_153),
.Y(n_181)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_119),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_127),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_185),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_152),
.A2(n_128),
.B(n_130),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_188),
.A2(n_126),
.B(n_127),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_156),
.A2(n_130),
.B1(n_126),
.B2(n_120),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_189),
.A2(n_145),
.B1(n_135),
.B2(n_106),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_128),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_191),
.B(n_198),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_184),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_194),
.B(n_163),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_197),
.B1(n_170),
.B2(n_167),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_160),
.B1(n_149),
.B2(n_146),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_209),
.B1(n_211),
.B2(n_169),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_SL g197 ( 
.A1(n_190),
.A2(n_144),
.B(n_134),
.C(n_154),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_137),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_155),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_207),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_142),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_208),
.C(n_216),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_138),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_204),
.B(n_171),
.Y(n_221)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_129),
.B(n_125),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_164),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_118),
.C(n_102),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_212),
.C(n_179),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_175),
.A2(n_85),
.B(n_66),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_104),
.C(n_66),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_174),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_218),
.A2(n_209),
.B(n_213),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_219),
.A2(n_226),
.B1(n_228),
.B2(n_207),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_222),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_221),
.B(n_224),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_189),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_223),
.A2(n_162),
.B(n_202),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_169),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_178),
.B1(n_171),
.B2(n_186),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_186),
.B1(n_162),
.B2(n_179),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_180),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_232),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g230 ( 
.A(n_192),
.B(n_183),
.CI(n_162),
.CON(n_230),
.SN(n_230)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_233),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_204),
.B(n_180),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_211),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_235),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_208),
.C(n_210),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_246),
.C(n_231),
.Y(n_259)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_216),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_244),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_198),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_245),
.A2(n_227),
.B1(n_228),
.B2(n_226),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_201),
.C(n_202),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_247),
.A2(n_249),
.B1(n_251),
.B2(n_219),
.Y(n_255)
);

NOR3xp33_ASAP7_75t_SL g248 ( 
.A(n_220),
.B(n_164),
.C(n_197),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_11),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_197),
.B(n_215),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_200),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_254),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_SL g251 ( 
.A(n_218),
.B(n_197),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_206),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_259),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_256),
.A2(n_263),
.B1(n_12),
.B2(n_16),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_242),
.A2(n_230),
.B1(n_218),
.B2(n_222),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_258),
.A2(n_252),
.B1(n_254),
.B2(n_244),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_230),
.C(n_214),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_262),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_214),
.C(n_183),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_181),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_264),
.B(n_266),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_243),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

OAI221xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_11),
.B1(n_16),
.B2(n_15),
.C(n_14),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_181),
.C(n_104),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_268),
.A2(n_240),
.B(n_250),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_275),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_SL g273 ( 
.A1(n_261),
.A2(n_242),
.B(n_248),
.C(n_237),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_273),
.A2(n_265),
.B1(n_260),
.B2(n_12),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_8),
.C(n_15),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_277),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_9),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_278),
.B(n_11),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_262),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_279),
.B(n_283),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_271),
.A2(n_259),
.B(n_265),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_273),
.B(n_104),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_3),
.Y(n_283)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_284),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_260),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_285),
.B(n_278),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_12),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_280),
.C(n_279),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_293),
.C(n_13),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_294),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_292),
.B(n_283),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_273),
.B(n_7),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_298),
.C(n_291),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_7),
.Y(n_297)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_297),
.Y(n_301)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_299),
.A2(n_300),
.B(n_4),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_296),
.A2(n_288),
.B(n_5),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_301),
.Y(n_303)
);


endmodule