module fake_jpeg_14404_n_489 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_489);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_489;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_SL g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_95),
.Y(n_101)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_55),
.Y(n_152)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_61),
.B(n_63),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_21),
.B(n_17),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_72),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_71),
.A2(n_33),
.B1(n_36),
.B2(n_26),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_32),
.B(n_16),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_73),
.Y(n_151)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

CKINVDCx9p33_ASAP7_75t_R g123 ( 
.A(n_75),
.Y(n_123)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

BUFx4f_ASAP7_75t_SL g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_24),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_78),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_84),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_22),
.B(n_16),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_91),
.Y(n_119)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_33),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_39),
.B1(n_44),
.B2(n_46),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_100),
.A2(n_23),
.B1(n_20),
.B2(n_95),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_44),
.C(n_48),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_108),
.A2(n_112),
.B(n_4),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_48),
.C(n_38),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_57),
.A2(n_25),
.B1(n_19),
.B2(n_30),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_114),
.A2(n_141),
.B(n_11),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_122),
.B(n_130),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_148),
.B1(n_149),
.B2(n_96),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_78),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_133),
.B(n_142),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_53),
.A2(n_30),
.B1(n_37),
.B2(n_36),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_75),
.Y(n_142)
);

AO22x1_ASAP7_75t_SL g143 ( 
.A1(n_71),
.A2(n_30),
.B1(n_35),
.B2(n_49),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_94),
.A2(n_46),
.B1(n_37),
.B2(n_20),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_52),
.A2(n_30),
.B1(n_35),
.B2(n_49),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_87),
.B1(n_55),
.B2(n_65),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_154),
.A2(n_167),
.B1(n_168),
.B2(n_172),
.Y(n_215)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_158),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_159),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_160),
.Y(n_228)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_161),
.Y(n_225)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_101),
.A2(n_51),
.B(n_77),
.C(n_90),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_SL g245 ( 
.A1(n_163),
.A2(n_173),
.B(n_165),
.C(n_188),
.Y(n_245)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_165),
.B(n_189),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_23),
.B1(n_70),
.B2(n_98),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_166),
.A2(n_174),
.B1(n_175),
.B2(n_186),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_80),
.B1(n_79),
.B2(n_69),
.Y(n_168)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_169),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_126),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_170),
.B(n_171),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_126),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_120),
.A2(n_82),
.B1(n_67),
.B2(n_62),
.Y(n_172)
);

AOI32xp33_ASAP7_75t_L g173 ( 
.A1(n_117),
.A2(n_91),
.A3(n_14),
.B1(n_13),
.B2(n_85),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_143),
.A2(n_49),
.B1(n_35),
.B2(n_3),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_116),
.A2(n_49),
.B1(n_35),
.B2(n_3),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_108),
.B(n_0),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_195),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_109),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_177),
.B(n_185),
.Y(n_238)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_179),
.Y(n_249)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_182),
.A2(n_188),
.B1(n_196),
.B2(n_177),
.Y(n_248)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_115),
.Y(n_183)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_184),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_109),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_L g187 ( 
.A1(n_113),
.A2(n_14),
.B(n_8),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_192),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_141),
.A2(n_14),
.B1(n_8),
.B2(n_10),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_119),
.B(n_7),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_139),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_194),
.A2(n_140),
.B1(n_146),
.B2(n_173),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_112),
.B(n_153),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_L g196 ( 
.A1(n_114),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_197),
.A2(n_198),
.B1(n_102),
.B2(n_147),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_102),
.A2(n_11),
.B1(n_12),
.B2(n_106),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_144),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_206),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_150),
.B(n_11),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_202),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_120),
.A2(n_121),
.B1(n_127),
.B2(n_135),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_201),
.A2(n_208),
.B1(n_159),
.B2(n_170),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_121),
.B(n_127),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_128),
.Y(n_203)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_203),
.Y(n_251)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_104),
.Y(n_204)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_106),
.B(n_103),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_132),
.C(n_124),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_115),
.B(n_140),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_144),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_146),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_135),
.A2(n_152),
.B1(n_111),
.B2(n_103),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_167),
.A2(n_152),
.B1(n_111),
.B2(n_138),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_209),
.A2(n_222),
.B1(n_233),
.B2(n_244),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_107),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_241),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_220),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_195),
.A2(n_197),
.B1(n_194),
.B2(n_176),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_232),
.B(n_245),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_202),
.A2(n_138),
.B1(n_145),
.B2(n_107),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_236),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_182),
.A2(n_147),
.B1(n_145),
.B2(n_140),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_239),
.A2(n_169),
.B(n_184),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_185),
.B(n_200),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_189),
.B(n_146),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_256),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_163),
.A2(n_160),
.B1(n_206),
.B2(n_156),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_246),
.B(n_254),
.Y(n_286)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_248),
.B(n_250),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_205),
.B(n_191),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_181),
.B(n_180),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_252),
.B(n_253),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_203),
.B(n_207),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_171),
.A2(n_205),
.B1(n_199),
.B2(n_157),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_254),
.A2(n_239),
.B1(n_218),
.B2(n_226),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_179),
.B(n_190),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_258),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_217),
.B(n_155),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_259),
.B(n_264),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_158),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_260),
.B(n_265),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_241),
.A2(n_160),
.B1(n_164),
.B2(n_204),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_261),
.A2(n_283),
.B1(n_293),
.B2(n_227),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_217),
.B(n_193),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_216),
.B(n_183),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_266),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_229),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_267),
.B(n_274),
.Y(n_324)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_227),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_269),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_212),
.B(n_161),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_270),
.B(n_271),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_222),
.B(n_162),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_272),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_209),
.A2(n_178),
.B1(n_184),
.B2(n_233),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_273),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_213),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_276),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_256),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_289),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_244),
.A2(n_238),
.B1(n_250),
.B2(n_219),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_280),
.A2(n_281),
.B(n_284),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_238),
.A2(n_221),
.B(n_245),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_214),
.Y(n_282)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_282),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_238),
.A2(n_248),
.B(n_210),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_284),
.A2(n_286),
.B(n_275),
.Y(n_321)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_214),
.Y(n_285)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_285),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_245),
.B(n_232),
.C(n_218),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_223),
.C(n_225),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_230),
.B(n_226),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_240),
.B(n_255),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_291),
.B(n_249),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_231),
.B(n_237),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_298),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_215),
.A2(n_235),
.B1(n_240),
.B2(n_242),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_230),
.Y(n_294)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_242),
.B(n_255),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_295),
.B(n_299),
.Y(n_337)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_211),
.Y(n_296)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_211),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_224),
.B(n_249),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_224),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_228),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_303),
.B(n_315),
.Y(n_358)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_308),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_278),
.B(n_228),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_309),
.B(n_312),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_310),
.A2(n_335),
.B1(n_287),
.B2(n_262),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_237),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_277),
.B(n_223),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_320),
.C(n_323),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_299),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_318),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_259),
.B(n_225),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_285),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_257),
.B(n_288),
.C(n_290),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_321),
.A2(n_330),
.B(n_280),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_257),
.B(n_290),
.C(n_281),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_295),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_326),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_327),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_270),
.B(n_263),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_329),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_286),
.A2(n_258),
.B(n_275),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_297),
.Y(n_331)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_331),
.Y(n_342)
);

INVx13_ASAP7_75t_L g334 ( 
.A(n_294),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_334),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_262),
.A2(n_297),
.B1(n_271),
.B2(n_283),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_264),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_336),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_279),
.B(n_263),
.Y(n_339)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_339),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_343),
.B(n_350),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_321),
.A2(n_286),
.B(n_290),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_344),
.A2(n_349),
.B(n_313),
.Y(n_374)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_328),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_348),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_335),
.A2(n_287),
.B1(n_297),
.B2(n_293),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_320),
.B(n_261),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_351),
.B(n_353),
.C(n_359),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_317),
.B(n_282),
.C(n_268),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_356),
.B(n_337),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_330),
.A2(n_276),
.B(n_272),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_357),
.A2(n_305),
.B(n_315),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_323),
.B(n_331),
.C(n_327),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_336),
.A2(n_266),
.B1(n_294),
.B2(n_300),
.Y(n_360)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_360),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_339),
.B(n_296),
.C(n_298),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_367),
.C(n_369),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_304),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_371),
.Y(n_379)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_301),
.Y(n_364)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_364),
.Y(n_382)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_301),
.Y(n_366)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_366),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_329),
.B(n_269),
.C(n_326),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_302),
.Y(n_368)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_368),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_332),
.B(n_304),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_302),
.Y(n_370)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_370),
.Y(n_390)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_306),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_310),
.A2(n_325),
.B1(n_333),
.B2(n_307),
.Y(n_372)
);

CKINVDCx14_ASAP7_75t_R g396 ( 
.A(n_372),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_374),
.A2(n_395),
.B(n_357),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_332),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_375),
.B(n_398),
.C(n_314),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_365),
.A2(n_318),
.B1(n_333),
.B2(n_337),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_377),
.A2(n_384),
.B1(n_387),
.B2(n_322),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_378),
.B(n_386),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_354),
.Y(n_380)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_380),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_361),
.B(n_324),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_381),
.B(n_397),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_345),
.A2(n_325),
.B1(n_307),
.B2(n_319),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_360),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_345),
.A2(n_324),
.B1(n_312),
.B2(n_305),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_340),
.Y(n_391)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_391),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_393),
.A2(n_308),
.B(n_316),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_358),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_394),
.B(n_399),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_355),
.A2(n_309),
.B(n_303),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_361),
.B(n_369),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_347),
.B(n_306),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_358),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_381),
.B(n_367),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_400),
.B(n_402),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_380),
.Y(n_401)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_401),
.Y(n_424)
);

AOI321xp33_ASAP7_75t_L g402 ( 
.A1(n_379),
.A2(n_342),
.A3(n_359),
.B1(n_344),
.B2(n_347),
.C(n_349),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_392),
.A2(n_355),
.B1(n_365),
.B2(n_341),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_403),
.A2(n_407),
.B1(n_384),
.B2(n_373),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_404),
.B(n_408),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_396),
.A2(n_341),
.B1(n_362),
.B2(n_371),
.Y(n_406)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_406),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_392),
.A2(n_350),
.B1(n_353),
.B2(n_342),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_375),
.B(n_356),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_394),
.A2(n_370),
.B1(n_368),
.B2(n_364),
.Y(n_409)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_409),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_366),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_411),
.B(n_414),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_377),
.B(n_348),
.Y(n_415)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_415),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_417),
.A2(n_420),
.B1(n_379),
.B2(n_395),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_373),
.A2(n_328),
.B1(n_352),
.B2(n_314),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_418),
.A2(n_385),
.B1(n_389),
.B2(n_390),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_383),
.B(n_338),
.C(n_322),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_419),
.B(n_422),
.C(n_378),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_383),
.B(n_388),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_374),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_388),
.B(n_338),
.C(n_316),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_426),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_407),
.A2(n_403),
.B1(n_386),
.B2(n_415),
.Y(n_427)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_416),
.A2(n_387),
.B1(n_399),
.B2(n_397),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_429),
.B(n_417),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_414),
.C(n_422),
.Y(n_447)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_412),
.Y(n_433)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_433),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_405),
.B(n_382),
.Y(n_434)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_434),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_382),
.Y(n_436)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_436),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_419),
.B(n_393),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_438),
.B(n_440),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_439),
.B(n_413),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_412),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_441),
.A2(n_390),
.B1(n_385),
.B2(n_389),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_443),
.B(n_452),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_445),
.B(n_430),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_450),
.Y(n_461)
);

INVxp33_ASAP7_75t_L g450 ( 
.A(n_434),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_451),
.B(n_453),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_425),
.A2(n_404),
.B1(n_402),
.B2(n_420),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_437),
.A2(n_418),
.B(n_421),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_411),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_455),
.A2(n_423),
.B(n_433),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_443),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_464),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_465),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_449),
.A2(n_431),
.B(n_432),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_459),
.A2(n_460),
.B(n_462),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_451),
.A2(n_428),
.B(n_427),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_453),
.A2(n_430),
.B(n_424),
.Y(n_463)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_463),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_447),
.B(n_435),
.C(n_428),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_435),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_442),
.A2(n_441),
.B1(n_436),
.B2(n_376),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_467),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_461),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_470),
.B(n_471),
.Y(n_477)
);

AOI322xp5_ASAP7_75t_L g471 ( 
.A1(n_462),
.A2(n_448),
.A3(n_444),
.B1(n_446),
.B2(n_454),
.C1(n_450),
.C2(n_445),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_452),
.C(n_448),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_473),
.B(n_476),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_408),
.C(n_376),
.Y(n_476)
);

OAI21x1_ASAP7_75t_L g478 ( 
.A1(n_472),
.A2(n_466),
.B(n_457),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_478),
.B(n_479),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_474),
.B(n_466),
.C(n_458),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_468),
.A2(n_458),
.B(n_376),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_480),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_477),
.A2(n_472),
.B(n_469),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_483),
.Y(n_485)
);

AOI321xp33_ASAP7_75t_L g486 ( 
.A1(n_484),
.A2(n_481),
.A3(n_475),
.B1(n_471),
.B2(n_334),
.C(n_311),
.Y(n_486)
);

O2A1O1Ixp33_ASAP7_75t_SL g487 ( 
.A1(n_486),
.A2(n_482),
.B(n_334),
.C(n_311),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_487),
.B(n_485),
.C(n_311),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_488),
.Y(n_489)
);


endmodule