module fake_jpeg_7080_n_280 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_10),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_36),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx12f_ASAP7_75t_SL g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp67_ASAP7_75t_R g53 ( 
.A(n_39),
.B(n_28),
.Y(n_53)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_36),
.Y(n_62)
);

CKINVDCx12_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_19),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_54),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_31),
.Y(n_80)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_21),
.B1(n_32),
.B2(n_18),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_26),
.B1(n_22),
.B2(n_16),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_39),
.B1(n_18),
.B2(n_32),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_62),
.A2(n_75),
.B(n_86),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_35),
.B1(n_37),
.B2(n_36),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_63),
.A2(n_65),
.B1(n_69),
.B2(n_73),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_56),
.B1(n_57),
.B2(n_47),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_32),
.B1(n_18),
.B2(n_21),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_83),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_78),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_41),
.B1(n_30),
.B2(n_17),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_41),
.B1(n_50),
.B2(n_30),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_34),
.B1(n_17),
.B2(n_35),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_76),
.B1(n_79),
.B2(n_84),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_34),
.B1(n_41),
.B2(n_19),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_37),
.C(n_35),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_82),
.C(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_31),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_34),
.B1(n_41),
.B2(n_25),
.Y(n_79)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_38),
.B(n_24),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_38),
.C(n_25),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_44),
.A2(n_34),
.B1(n_23),
.B2(n_26),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_38),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_92),
.B1(n_20),
.B2(n_27),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_22),
.B1(n_31),
.B2(n_27),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_91),
.B1(n_80),
.B2(n_63),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_53),
.A2(n_29),
.B(n_38),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_54),
.A2(n_31),
.B1(n_27),
.B2(n_20),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_105),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_107),
.B1(n_83),
.B2(n_68),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_104),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_60),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_24),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

NAND3xp33_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_62),
.C(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_110),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_24),
.C(n_0),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_119),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_24),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_111),
.Y(n_137)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_24),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_66),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_0),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_59),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_82),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_118),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_L g119 ( 
.A1(n_63),
.A2(n_15),
.B(n_2),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g120 ( 
.A1(n_63),
.A2(n_15),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_140),
.B1(n_148),
.B2(n_86),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_114),
.A2(n_64),
.B1(n_92),
.B2(n_68),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_129),
.Y(n_157)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_100),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_133),
.B(n_139),
.Y(n_152)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_135),
.Y(n_175)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_110),
.B1(n_105),
.B2(n_93),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_98),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_111),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_71),
.B1(n_75),
.B2(n_59),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_71),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_149),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_147),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_102),
.A2(n_87),
.B1(n_88),
.B2(n_86),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_81),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_119),
.B(n_106),
.C(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_150),
.B(n_153),
.Y(n_198)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_125),
.A2(n_107),
.B1(n_96),
.B2(n_103),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_164),
.B1(n_167),
.B2(n_126),
.Y(n_181)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_103),
.C(n_113),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_172),
.C(n_130),
.Y(n_189)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_165),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_141),
.A2(n_147),
.B1(n_128),
.B2(n_149),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_170),
.B(n_173),
.Y(n_183)
);

OR2x4_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_120),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_101),
.B(n_144),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_108),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_94),
.C(n_101),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_176),
.Y(n_191)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_175),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_188),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_168),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_98),
.B1(n_95),
.B2(n_136),
.Y(n_182)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_143),
.B(n_135),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_186),
.B(n_195),
.Y(n_205)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_196),
.C(n_201),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_171),
.A2(n_174),
.B1(n_157),
.B2(n_150),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_186),
.B1(n_194),
.B2(n_198),
.Y(n_214)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_194),
.Y(n_209)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_124),
.B(n_122),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_130),
.C(n_122),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_122),
.B1(n_93),
.B2(n_81),
.Y(n_197)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_200),
.Y(n_216)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_72),
.C(n_2),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_172),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_207),
.B(n_214),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_176),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_210),
.Y(n_237)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_217),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_161),
.C(n_159),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_219),
.C(n_201),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_183),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_168),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_179),
.B1(n_185),
.B2(n_151),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_184),
.C(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_179),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_197),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_R g222 ( 
.A(n_207),
.B(n_190),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_SL g238 ( 
.A(n_222),
.B(n_230),
.C(n_231),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_215),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_234),
.C(n_212),
.Y(n_242)
);

OA21x2_ASAP7_75t_L g227 ( 
.A1(n_218),
.A2(n_169),
.B(n_202),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_227),
.B(n_221),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_211),
.A2(n_199),
.B1(n_202),
.B2(n_169),
.Y(n_228)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_214),
.B(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_208),
.A2(n_160),
.B1(n_165),
.B2(n_159),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_217),
.B1(n_203),
.B2(n_5),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_219),
.B(n_160),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_72),
.C(n_4),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_216),
.C(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_246),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_244),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_237),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_204),
.C(n_206),
.Y(n_244)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_14),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g248 ( 
.A(n_225),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_248),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_14),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_235),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_243),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_250),
.B(n_251),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_247),
.B(n_229),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_238),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_255),
.B(n_256),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_244),
.B(n_236),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_226),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_261),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_226),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_231),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_253),
.C(n_227),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_239),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_264),
.A2(n_266),
.B(n_254),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_227),
.B(n_258),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_267),
.B(n_268),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_262),
.B1(n_6),
.B2(n_7),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_L g276 ( 
.A1(n_273),
.A2(n_1),
.B(n_7),
.Y(n_276)
);

O2A1O1Ixp33_ASAP7_75t_SL g275 ( 
.A1(n_272),
.A2(n_269),
.B(n_7),
.C(n_8),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_276),
.C(n_274),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_9),
.B(n_10),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_9),
.B(n_11),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_11),
.Y(n_280)
);


endmodule